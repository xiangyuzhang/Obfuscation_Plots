module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate911(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate912(.a(gate12inter0), .b(s_52), .O(gate12inter1));
  and2  gate913(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate914(.a(s_52), .O(gate12inter3));
  inv1  gate915(.a(s_53), .O(gate12inter4));
  nand2 gate916(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate917(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate918(.a(G7), .O(gate12inter7));
  inv1  gate919(.a(G8), .O(gate12inter8));
  nand2 gate920(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate921(.a(s_53), .b(gate12inter3), .O(gate12inter10));
  nor2  gate922(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate923(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate924(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1513(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1514(.a(gate22inter0), .b(s_138), .O(gate22inter1));
  and2  gate1515(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1516(.a(s_138), .O(gate22inter3));
  inv1  gate1517(.a(s_139), .O(gate22inter4));
  nand2 gate1518(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1519(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1520(.a(G27), .O(gate22inter7));
  inv1  gate1521(.a(G28), .O(gate22inter8));
  nand2 gate1522(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1523(.a(s_139), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1524(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1525(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1526(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate617(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate618(.a(gate26inter0), .b(s_10), .O(gate26inter1));
  and2  gate619(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate620(.a(s_10), .O(gate26inter3));
  inv1  gate621(.a(s_11), .O(gate26inter4));
  nand2 gate622(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate623(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate624(.a(G9), .O(gate26inter7));
  inv1  gate625(.a(G13), .O(gate26inter8));
  nand2 gate626(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate627(.a(s_11), .b(gate26inter3), .O(gate26inter10));
  nor2  gate628(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate629(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate630(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1569(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1570(.a(gate33inter0), .b(s_146), .O(gate33inter1));
  and2  gate1571(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1572(.a(s_146), .O(gate33inter3));
  inv1  gate1573(.a(s_147), .O(gate33inter4));
  nand2 gate1574(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1575(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1576(.a(G17), .O(gate33inter7));
  inv1  gate1577(.a(G21), .O(gate33inter8));
  nand2 gate1578(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1579(.a(s_147), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1580(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1581(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1582(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1219(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1220(.a(gate34inter0), .b(s_96), .O(gate34inter1));
  and2  gate1221(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1222(.a(s_96), .O(gate34inter3));
  inv1  gate1223(.a(s_97), .O(gate34inter4));
  nand2 gate1224(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1225(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1226(.a(G25), .O(gate34inter7));
  inv1  gate1227(.a(G29), .O(gate34inter8));
  nand2 gate1228(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1229(.a(s_97), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1230(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1231(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1232(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate827(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate828(.a(gate36inter0), .b(s_40), .O(gate36inter1));
  and2  gate829(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate830(.a(s_40), .O(gate36inter3));
  inv1  gate831(.a(s_41), .O(gate36inter4));
  nand2 gate832(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate833(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate834(.a(G26), .O(gate36inter7));
  inv1  gate835(.a(G30), .O(gate36inter8));
  nand2 gate836(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate837(.a(s_41), .b(gate36inter3), .O(gate36inter10));
  nor2  gate838(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate839(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate840(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1317(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1318(.a(gate38inter0), .b(s_110), .O(gate38inter1));
  and2  gate1319(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1320(.a(s_110), .O(gate38inter3));
  inv1  gate1321(.a(s_111), .O(gate38inter4));
  nand2 gate1322(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1323(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1324(.a(G27), .O(gate38inter7));
  inv1  gate1325(.a(G31), .O(gate38inter8));
  nand2 gate1326(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1327(.a(s_111), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1328(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1329(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1330(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate743(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate744(.a(gate39inter0), .b(s_28), .O(gate39inter1));
  and2  gate745(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate746(.a(s_28), .O(gate39inter3));
  inv1  gate747(.a(s_29), .O(gate39inter4));
  nand2 gate748(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate749(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate750(.a(G20), .O(gate39inter7));
  inv1  gate751(.a(G24), .O(gate39inter8));
  nand2 gate752(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate753(.a(s_29), .b(gate39inter3), .O(gate39inter10));
  nor2  gate754(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate755(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate756(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1177(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1178(.a(gate45inter0), .b(s_90), .O(gate45inter1));
  and2  gate1179(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1180(.a(s_90), .O(gate45inter3));
  inv1  gate1181(.a(s_91), .O(gate45inter4));
  nand2 gate1182(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1183(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1184(.a(G5), .O(gate45inter7));
  inv1  gate1185(.a(G272), .O(gate45inter8));
  nand2 gate1186(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1187(.a(s_91), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1188(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1189(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1190(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate575(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate576(.a(gate48inter0), .b(s_4), .O(gate48inter1));
  and2  gate577(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate578(.a(s_4), .O(gate48inter3));
  inv1  gate579(.a(s_5), .O(gate48inter4));
  nand2 gate580(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate581(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate582(.a(G8), .O(gate48inter7));
  inv1  gate583(.a(G275), .O(gate48inter8));
  nand2 gate584(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate585(.a(s_5), .b(gate48inter3), .O(gate48inter10));
  nor2  gate586(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate587(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate588(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate939(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate940(.a(gate63inter0), .b(s_56), .O(gate63inter1));
  and2  gate941(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate942(.a(s_56), .O(gate63inter3));
  inv1  gate943(.a(s_57), .O(gate63inter4));
  nand2 gate944(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate945(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate946(.a(G23), .O(gate63inter7));
  inv1  gate947(.a(G299), .O(gate63inter8));
  nand2 gate948(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate949(.a(s_57), .b(gate63inter3), .O(gate63inter10));
  nor2  gate950(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate951(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate952(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1611(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1612(.a(gate67inter0), .b(s_152), .O(gate67inter1));
  and2  gate1613(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1614(.a(s_152), .O(gate67inter3));
  inv1  gate1615(.a(s_153), .O(gate67inter4));
  nand2 gate1616(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1617(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1618(.a(G27), .O(gate67inter7));
  inv1  gate1619(.a(G305), .O(gate67inter8));
  nand2 gate1620(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1621(.a(s_153), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1622(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1623(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1624(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate841(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate842(.a(gate71inter0), .b(s_42), .O(gate71inter1));
  and2  gate843(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate844(.a(s_42), .O(gate71inter3));
  inv1  gate845(.a(s_43), .O(gate71inter4));
  nand2 gate846(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate847(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate848(.a(G31), .O(gate71inter7));
  inv1  gate849(.a(G311), .O(gate71inter8));
  nand2 gate850(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate851(.a(s_43), .b(gate71inter3), .O(gate71inter10));
  nor2  gate852(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate853(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate854(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1653(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1654(.a(gate86inter0), .b(s_158), .O(gate86inter1));
  and2  gate1655(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1656(.a(s_158), .O(gate86inter3));
  inv1  gate1657(.a(s_159), .O(gate86inter4));
  nand2 gate1658(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1659(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1660(.a(G8), .O(gate86inter7));
  inv1  gate1661(.a(G332), .O(gate86inter8));
  nand2 gate1662(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1663(.a(s_159), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1664(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1665(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1666(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1093(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1094(.a(gate88inter0), .b(s_78), .O(gate88inter1));
  and2  gate1095(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1096(.a(s_78), .O(gate88inter3));
  inv1  gate1097(.a(s_79), .O(gate88inter4));
  nand2 gate1098(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1099(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1100(.a(G16), .O(gate88inter7));
  inv1  gate1101(.a(G335), .O(gate88inter8));
  nand2 gate1102(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1103(.a(s_79), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1104(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1105(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1106(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate673(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate674(.a(gate92inter0), .b(s_18), .O(gate92inter1));
  and2  gate675(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate676(.a(s_18), .O(gate92inter3));
  inv1  gate677(.a(s_19), .O(gate92inter4));
  nand2 gate678(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate679(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate680(.a(G29), .O(gate92inter7));
  inv1  gate681(.a(G341), .O(gate92inter8));
  nand2 gate682(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate683(.a(s_19), .b(gate92inter3), .O(gate92inter10));
  nor2  gate684(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate685(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate686(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1471(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1472(.a(gate93inter0), .b(s_132), .O(gate93inter1));
  and2  gate1473(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1474(.a(s_132), .O(gate93inter3));
  inv1  gate1475(.a(s_133), .O(gate93inter4));
  nand2 gate1476(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1477(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1478(.a(G18), .O(gate93inter7));
  inv1  gate1479(.a(G344), .O(gate93inter8));
  nand2 gate1480(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1481(.a(s_133), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1482(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1483(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1484(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1247(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1248(.a(gate96inter0), .b(s_100), .O(gate96inter1));
  and2  gate1249(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1250(.a(s_100), .O(gate96inter3));
  inv1  gate1251(.a(s_101), .O(gate96inter4));
  nand2 gate1252(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1253(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1254(.a(G30), .O(gate96inter7));
  inv1  gate1255(.a(G347), .O(gate96inter8));
  nand2 gate1256(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1257(.a(s_101), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1258(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1259(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1260(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate729(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate730(.a(gate106inter0), .b(s_26), .O(gate106inter1));
  and2  gate731(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate732(.a(s_26), .O(gate106inter3));
  inv1  gate733(.a(s_27), .O(gate106inter4));
  nand2 gate734(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate735(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate736(.a(G364), .O(gate106inter7));
  inv1  gate737(.a(G365), .O(gate106inter8));
  nand2 gate738(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate739(.a(s_27), .b(gate106inter3), .O(gate106inter10));
  nor2  gate740(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate741(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate742(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate561(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate562(.a(gate108inter0), .b(s_2), .O(gate108inter1));
  and2  gate563(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate564(.a(s_2), .O(gate108inter3));
  inv1  gate565(.a(s_3), .O(gate108inter4));
  nand2 gate566(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate567(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate568(.a(G368), .O(gate108inter7));
  inv1  gate569(.a(G369), .O(gate108inter8));
  nand2 gate570(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate571(.a(s_3), .b(gate108inter3), .O(gate108inter10));
  nor2  gate572(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate573(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate574(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1429(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1430(.a(gate113inter0), .b(s_126), .O(gate113inter1));
  and2  gate1431(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1432(.a(s_126), .O(gate113inter3));
  inv1  gate1433(.a(s_127), .O(gate113inter4));
  nand2 gate1434(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1435(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1436(.a(G378), .O(gate113inter7));
  inv1  gate1437(.a(G379), .O(gate113inter8));
  nand2 gate1438(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1439(.a(s_127), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1440(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1441(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1442(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1415(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1416(.a(gate117inter0), .b(s_124), .O(gate117inter1));
  and2  gate1417(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1418(.a(s_124), .O(gate117inter3));
  inv1  gate1419(.a(s_125), .O(gate117inter4));
  nand2 gate1420(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1421(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1422(.a(G386), .O(gate117inter7));
  inv1  gate1423(.a(G387), .O(gate117inter8));
  nand2 gate1424(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1425(.a(s_125), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1426(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1427(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1428(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate701(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate702(.a(gate120inter0), .b(s_22), .O(gate120inter1));
  and2  gate703(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate704(.a(s_22), .O(gate120inter3));
  inv1  gate705(.a(s_23), .O(gate120inter4));
  nand2 gate706(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate707(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate708(.a(G392), .O(gate120inter7));
  inv1  gate709(.a(G393), .O(gate120inter8));
  nand2 gate710(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate711(.a(s_23), .b(gate120inter3), .O(gate120inter10));
  nor2  gate712(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate713(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate714(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1261(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1262(.a(gate122inter0), .b(s_102), .O(gate122inter1));
  and2  gate1263(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1264(.a(s_102), .O(gate122inter3));
  inv1  gate1265(.a(s_103), .O(gate122inter4));
  nand2 gate1266(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1267(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1268(.a(G396), .O(gate122inter7));
  inv1  gate1269(.a(G397), .O(gate122inter8));
  nand2 gate1270(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1271(.a(s_103), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1272(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1273(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1274(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1597(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1598(.a(gate125inter0), .b(s_150), .O(gate125inter1));
  and2  gate1599(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1600(.a(s_150), .O(gate125inter3));
  inv1  gate1601(.a(s_151), .O(gate125inter4));
  nand2 gate1602(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1603(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1604(.a(G402), .O(gate125inter7));
  inv1  gate1605(.a(G403), .O(gate125inter8));
  nand2 gate1606(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1607(.a(s_151), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1608(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1609(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1610(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate631(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate632(.a(gate126inter0), .b(s_12), .O(gate126inter1));
  and2  gate633(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate634(.a(s_12), .O(gate126inter3));
  inv1  gate635(.a(s_13), .O(gate126inter4));
  nand2 gate636(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate637(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate638(.a(G404), .O(gate126inter7));
  inv1  gate639(.a(G405), .O(gate126inter8));
  nand2 gate640(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate641(.a(s_13), .b(gate126inter3), .O(gate126inter10));
  nor2  gate642(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate643(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate644(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate869(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate870(.a(gate127inter0), .b(s_46), .O(gate127inter1));
  and2  gate871(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate872(.a(s_46), .O(gate127inter3));
  inv1  gate873(.a(s_47), .O(gate127inter4));
  nand2 gate874(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate875(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate876(.a(G406), .O(gate127inter7));
  inv1  gate877(.a(G407), .O(gate127inter8));
  nand2 gate878(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate879(.a(s_47), .b(gate127inter3), .O(gate127inter10));
  nor2  gate880(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate881(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate882(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate603(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate604(.a(gate129inter0), .b(s_8), .O(gate129inter1));
  and2  gate605(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate606(.a(s_8), .O(gate129inter3));
  inv1  gate607(.a(s_9), .O(gate129inter4));
  nand2 gate608(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate609(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate610(.a(G410), .O(gate129inter7));
  inv1  gate611(.a(G411), .O(gate129inter8));
  nand2 gate612(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate613(.a(s_9), .b(gate129inter3), .O(gate129inter10));
  nor2  gate614(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate615(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate616(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1275(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1276(.a(gate131inter0), .b(s_104), .O(gate131inter1));
  and2  gate1277(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1278(.a(s_104), .O(gate131inter3));
  inv1  gate1279(.a(s_105), .O(gate131inter4));
  nand2 gate1280(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1281(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1282(.a(G414), .O(gate131inter7));
  inv1  gate1283(.a(G415), .O(gate131inter8));
  nand2 gate1284(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1285(.a(s_105), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1286(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1287(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1288(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1667(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1668(.a(gate136inter0), .b(s_160), .O(gate136inter1));
  and2  gate1669(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1670(.a(s_160), .O(gate136inter3));
  inv1  gate1671(.a(s_161), .O(gate136inter4));
  nand2 gate1672(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1673(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1674(.a(G424), .O(gate136inter7));
  inv1  gate1675(.a(G425), .O(gate136inter8));
  nand2 gate1676(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1677(.a(s_161), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1678(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1679(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1680(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1457(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1458(.a(gate139inter0), .b(s_130), .O(gate139inter1));
  and2  gate1459(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1460(.a(s_130), .O(gate139inter3));
  inv1  gate1461(.a(s_131), .O(gate139inter4));
  nand2 gate1462(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1463(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1464(.a(G438), .O(gate139inter7));
  inv1  gate1465(.a(G441), .O(gate139inter8));
  nand2 gate1466(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1467(.a(s_131), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1468(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1469(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1470(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate659(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate660(.a(gate147inter0), .b(s_16), .O(gate147inter1));
  and2  gate661(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate662(.a(s_16), .O(gate147inter3));
  inv1  gate663(.a(s_17), .O(gate147inter4));
  nand2 gate664(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate665(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate666(.a(G486), .O(gate147inter7));
  inv1  gate667(.a(G489), .O(gate147inter8));
  nand2 gate668(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate669(.a(s_17), .b(gate147inter3), .O(gate147inter10));
  nor2  gate670(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate671(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate672(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1289(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1290(.a(gate151inter0), .b(s_106), .O(gate151inter1));
  and2  gate1291(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1292(.a(s_106), .O(gate151inter3));
  inv1  gate1293(.a(s_107), .O(gate151inter4));
  nand2 gate1294(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1295(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1296(.a(G510), .O(gate151inter7));
  inv1  gate1297(.a(G513), .O(gate151inter8));
  nand2 gate1298(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1299(.a(s_107), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1300(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1301(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1302(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1345(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1346(.a(gate154inter0), .b(s_114), .O(gate154inter1));
  and2  gate1347(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1348(.a(s_114), .O(gate154inter3));
  inv1  gate1349(.a(s_115), .O(gate154inter4));
  nand2 gate1350(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1351(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1352(.a(G429), .O(gate154inter7));
  inv1  gate1353(.a(G522), .O(gate154inter8));
  nand2 gate1354(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1355(.a(s_115), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1356(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1357(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1358(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1499(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1500(.a(gate155inter0), .b(s_136), .O(gate155inter1));
  and2  gate1501(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1502(.a(s_136), .O(gate155inter3));
  inv1  gate1503(.a(s_137), .O(gate155inter4));
  nand2 gate1504(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1505(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1506(.a(G432), .O(gate155inter7));
  inv1  gate1507(.a(G525), .O(gate155inter8));
  nand2 gate1508(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1509(.a(s_137), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1510(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1511(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1512(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate855(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate856(.a(gate158inter0), .b(s_44), .O(gate158inter1));
  and2  gate857(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate858(.a(s_44), .O(gate158inter3));
  inv1  gate859(.a(s_45), .O(gate158inter4));
  nand2 gate860(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate861(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate862(.a(G441), .O(gate158inter7));
  inv1  gate863(.a(G528), .O(gate158inter8));
  nand2 gate864(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate865(.a(s_45), .b(gate158inter3), .O(gate158inter10));
  nor2  gate866(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate867(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate868(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate715(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate716(.a(gate164inter0), .b(s_24), .O(gate164inter1));
  and2  gate717(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate718(.a(s_24), .O(gate164inter3));
  inv1  gate719(.a(s_25), .O(gate164inter4));
  nand2 gate720(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate721(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate722(.a(G459), .O(gate164inter7));
  inv1  gate723(.a(G537), .O(gate164inter8));
  nand2 gate724(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate725(.a(s_25), .b(gate164inter3), .O(gate164inter10));
  nor2  gate726(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate727(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate728(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate813(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate814(.a(gate166inter0), .b(s_38), .O(gate166inter1));
  and2  gate815(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate816(.a(s_38), .O(gate166inter3));
  inv1  gate817(.a(s_39), .O(gate166inter4));
  nand2 gate818(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate819(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate820(.a(G465), .O(gate166inter7));
  inv1  gate821(.a(G540), .O(gate166inter8));
  nand2 gate822(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate823(.a(s_39), .b(gate166inter3), .O(gate166inter10));
  nor2  gate824(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate825(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate826(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate757(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate758(.a(gate169inter0), .b(s_30), .O(gate169inter1));
  and2  gate759(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate760(.a(s_30), .O(gate169inter3));
  inv1  gate761(.a(s_31), .O(gate169inter4));
  nand2 gate762(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate763(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate764(.a(G474), .O(gate169inter7));
  inv1  gate765(.a(G546), .O(gate169inter8));
  nand2 gate766(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate767(.a(s_31), .b(gate169inter3), .O(gate169inter10));
  nor2  gate768(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate769(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate770(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1485(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1486(.a(gate184inter0), .b(s_134), .O(gate184inter1));
  and2  gate1487(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1488(.a(s_134), .O(gate184inter3));
  inv1  gate1489(.a(s_135), .O(gate184inter4));
  nand2 gate1490(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1491(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1492(.a(G519), .O(gate184inter7));
  inv1  gate1493(.a(G567), .O(gate184inter8));
  nand2 gate1494(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1495(.a(s_135), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1496(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1497(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1498(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate785(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate786(.a(gate189inter0), .b(s_34), .O(gate189inter1));
  and2  gate787(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate788(.a(s_34), .O(gate189inter3));
  inv1  gate789(.a(s_35), .O(gate189inter4));
  nand2 gate790(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate791(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate792(.a(G578), .O(gate189inter7));
  inv1  gate793(.a(G579), .O(gate189inter8));
  nand2 gate794(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate795(.a(s_35), .b(gate189inter3), .O(gate189inter10));
  nor2  gate796(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate797(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate798(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1191(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1192(.a(gate192inter0), .b(s_92), .O(gate192inter1));
  and2  gate1193(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1194(.a(s_92), .O(gate192inter3));
  inv1  gate1195(.a(s_93), .O(gate192inter4));
  nand2 gate1196(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1197(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1198(.a(G584), .O(gate192inter7));
  inv1  gate1199(.a(G585), .O(gate192inter8));
  nand2 gate1200(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1201(.a(s_93), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1202(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1203(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1204(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1625(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1626(.a(gate196inter0), .b(s_154), .O(gate196inter1));
  and2  gate1627(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1628(.a(s_154), .O(gate196inter3));
  inv1  gate1629(.a(s_155), .O(gate196inter4));
  nand2 gate1630(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1631(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1632(.a(G592), .O(gate196inter7));
  inv1  gate1633(.a(G593), .O(gate196inter8));
  nand2 gate1634(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1635(.a(s_155), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1636(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1637(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1638(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate771(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate772(.a(gate204inter0), .b(s_32), .O(gate204inter1));
  and2  gate773(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate774(.a(s_32), .O(gate204inter3));
  inv1  gate775(.a(s_33), .O(gate204inter4));
  nand2 gate776(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate777(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate778(.a(G607), .O(gate204inter7));
  inv1  gate779(.a(G617), .O(gate204inter8));
  nand2 gate780(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate781(.a(s_33), .b(gate204inter3), .O(gate204inter10));
  nor2  gate782(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate783(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate784(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1163(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1164(.a(gate209inter0), .b(s_88), .O(gate209inter1));
  and2  gate1165(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1166(.a(s_88), .O(gate209inter3));
  inv1  gate1167(.a(s_89), .O(gate209inter4));
  nand2 gate1168(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1169(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1170(.a(G602), .O(gate209inter7));
  inv1  gate1171(.a(G666), .O(gate209inter8));
  nand2 gate1172(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1173(.a(s_89), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1174(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1175(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1176(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1233(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1234(.a(gate210inter0), .b(s_98), .O(gate210inter1));
  and2  gate1235(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1236(.a(s_98), .O(gate210inter3));
  inv1  gate1237(.a(s_99), .O(gate210inter4));
  nand2 gate1238(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1239(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1240(.a(G607), .O(gate210inter7));
  inv1  gate1241(.a(G666), .O(gate210inter8));
  nand2 gate1242(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1243(.a(s_99), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1244(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1245(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1246(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1065(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1066(.a(gate211inter0), .b(s_74), .O(gate211inter1));
  and2  gate1067(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1068(.a(s_74), .O(gate211inter3));
  inv1  gate1069(.a(s_75), .O(gate211inter4));
  nand2 gate1070(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1071(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1072(.a(G612), .O(gate211inter7));
  inv1  gate1073(.a(G669), .O(gate211inter8));
  nand2 gate1074(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1075(.a(s_75), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1076(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1077(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1078(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1023(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1024(.a(gate212inter0), .b(s_68), .O(gate212inter1));
  and2  gate1025(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1026(.a(s_68), .O(gate212inter3));
  inv1  gate1027(.a(s_69), .O(gate212inter4));
  nand2 gate1028(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1029(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1030(.a(G617), .O(gate212inter7));
  inv1  gate1031(.a(G669), .O(gate212inter8));
  nand2 gate1032(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1033(.a(s_69), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1034(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1035(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1036(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1037(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1038(.a(gate215inter0), .b(s_70), .O(gate215inter1));
  and2  gate1039(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1040(.a(s_70), .O(gate215inter3));
  inv1  gate1041(.a(s_71), .O(gate215inter4));
  nand2 gate1042(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1043(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1044(.a(G607), .O(gate215inter7));
  inv1  gate1045(.a(G675), .O(gate215inter8));
  nand2 gate1046(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1047(.a(s_71), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1048(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1049(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1050(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1373(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1374(.a(gate227inter0), .b(s_118), .O(gate227inter1));
  and2  gate1375(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1376(.a(s_118), .O(gate227inter3));
  inv1  gate1377(.a(s_119), .O(gate227inter4));
  nand2 gate1378(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1379(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1380(.a(G694), .O(gate227inter7));
  inv1  gate1381(.a(G695), .O(gate227inter8));
  nand2 gate1382(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1383(.a(s_119), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1384(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1385(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1386(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate589(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate590(.a(gate231inter0), .b(s_6), .O(gate231inter1));
  and2  gate591(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate592(.a(s_6), .O(gate231inter3));
  inv1  gate593(.a(s_7), .O(gate231inter4));
  nand2 gate594(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate595(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate596(.a(G702), .O(gate231inter7));
  inv1  gate597(.a(G703), .O(gate231inter8));
  nand2 gate598(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate599(.a(s_7), .b(gate231inter3), .O(gate231inter10));
  nor2  gate600(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate601(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate602(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate687(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate688(.a(gate233inter0), .b(s_20), .O(gate233inter1));
  and2  gate689(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate690(.a(s_20), .O(gate233inter3));
  inv1  gate691(.a(s_21), .O(gate233inter4));
  nand2 gate692(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate693(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate694(.a(G242), .O(gate233inter7));
  inv1  gate695(.a(G718), .O(gate233inter8));
  nand2 gate696(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate697(.a(s_21), .b(gate233inter3), .O(gate233inter10));
  nor2  gate698(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate699(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate700(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate897(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate898(.a(gate248inter0), .b(s_50), .O(gate248inter1));
  and2  gate899(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate900(.a(s_50), .O(gate248inter3));
  inv1  gate901(.a(s_51), .O(gate248inter4));
  nand2 gate902(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate903(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate904(.a(G727), .O(gate248inter7));
  inv1  gate905(.a(G739), .O(gate248inter8));
  nand2 gate906(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate907(.a(s_51), .b(gate248inter3), .O(gate248inter10));
  nor2  gate908(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate909(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate910(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate547(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate548(.a(gate252inter0), .b(s_0), .O(gate252inter1));
  and2  gate549(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate550(.a(s_0), .O(gate252inter3));
  inv1  gate551(.a(s_1), .O(gate252inter4));
  nand2 gate552(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate553(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate554(.a(G709), .O(gate252inter7));
  inv1  gate555(.a(G745), .O(gate252inter8));
  nand2 gate556(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate557(.a(s_1), .b(gate252inter3), .O(gate252inter10));
  nor2  gate558(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate559(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate560(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate799(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate800(.a(gate253inter0), .b(s_36), .O(gate253inter1));
  and2  gate801(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate802(.a(s_36), .O(gate253inter3));
  inv1  gate803(.a(s_37), .O(gate253inter4));
  nand2 gate804(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate805(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate806(.a(G260), .O(gate253inter7));
  inv1  gate807(.a(G748), .O(gate253inter8));
  nand2 gate808(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate809(.a(s_37), .b(gate253inter3), .O(gate253inter10));
  nor2  gate810(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate811(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate812(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1331(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1332(.a(gate264inter0), .b(s_112), .O(gate264inter1));
  and2  gate1333(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1334(.a(s_112), .O(gate264inter3));
  inv1  gate1335(.a(s_113), .O(gate264inter4));
  nand2 gate1336(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1337(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1338(.a(G768), .O(gate264inter7));
  inv1  gate1339(.a(G769), .O(gate264inter8));
  nand2 gate1340(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1341(.a(s_113), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1342(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1343(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1344(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate925(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate926(.a(gate265inter0), .b(s_54), .O(gate265inter1));
  and2  gate927(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate928(.a(s_54), .O(gate265inter3));
  inv1  gate929(.a(s_55), .O(gate265inter4));
  nand2 gate930(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate931(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate932(.a(G642), .O(gate265inter7));
  inv1  gate933(.a(G770), .O(gate265inter8));
  nand2 gate934(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate935(.a(s_55), .b(gate265inter3), .O(gate265inter10));
  nor2  gate936(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate937(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate938(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1639(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1640(.a(gate284inter0), .b(s_156), .O(gate284inter1));
  and2  gate1641(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1642(.a(s_156), .O(gate284inter3));
  inv1  gate1643(.a(s_157), .O(gate284inter4));
  nand2 gate1644(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1645(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1646(.a(G785), .O(gate284inter7));
  inv1  gate1647(.a(G809), .O(gate284inter8));
  nand2 gate1648(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1649(.a(s_157), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1650(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1651(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1652(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate645(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate646(.a(gate290inter0), .b(s_14), .O(gate290inter1));
  and2  gate647(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate648(.a(s_14), .O(gate290inter3));
  inv1  gate649(.a(s_15), .O(gate290inter4));
  nand2 gate650(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate651(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate652(.a(G820), .O(gate290inter7));
  inv1  gate653(.a(G821), .O(gate290inter8));
  nand2 gate654(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate655(.a(s_15), .b(gate290inter3), .O(gate290inter10));
  nor2  gate656(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate657(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate658(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1583(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1584(.a(gate292inter0), .b(s_148), .O(gate292inter1));
  and2  gate1585(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1586(.a(s_148), .O(gate292inter3));
  inv1  gate1587(.a(s_149), .O(gate292inter4));
  nand2 gate1588(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1589(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1590(.a(G824), .O(gate292inter7));
  inv1  gate1591(.a(G825), .O(gate292inter8));
  nand2 gate1592(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1593(.a(s_149), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1594(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1595(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1596(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate967(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate968(.a(gate389inter0), .b(s_60), .O(gate389inter1));
  and2  gate969(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate970(.a(s_60), .O(gate389inter3));
  inv1  gate971(.a(s_61), .O(gate389inter4));
  nand2 gate972(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate973(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate974(.a(G3), .O(gate389inter7));
  inv1  gate975(.a(G1042), .O(gate389inter8));
  nand2 gate976(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate977(.a(s_61), .b(gate389inter3), .O(gate389inter10));
  nor2  gate978(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate979(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate980(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1359(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1360(.a(gate394inter0), .b(s_116), .O(gate394inter1));
  and2  gate1361(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1362(.a(s_116), .O(gate394inter3));
  inv1  gate1363(.a(s_117), .O(gate394inter4));
  nand2 gate1364(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1365(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1366(.a(G8), .O(gate394inter7));
  inv1  gate1367(.a(G1057), .O(gate394inter8));
  nand2 gate1368(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1369(.a(s_117), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1370(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1371(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1372(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate981(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate982(.a(gate395inter0), .b(s_62), .O(gate395inter1));
  and2  gate983(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate984(.a(s_62), .O(gate395inter3));
  inv1  gate985(.a(s_63), .O(gate395inter4));
  nand2 gate986(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate987(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate988(.a(G9), .O(gate395inter7));
  inv1  gate989(.a(G1060), .O(gate395inter8));
  nand2 gate990(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate991(.a(s_63), .b(gate395inter3), .O(gate395inter10));
  nor2  gate992(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate993(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate994(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1079(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1080(.a(gate411inter0), .b(s_76), .O(gate411inter1));
  and2  gate1081(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1082(.a(s_76), .O(gate411inter3));
  inv1  gate1083(.a(s_77), .O(gate411inter4));
  nand2 gate1084(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1085(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1086(.a(G25), .O(gate411inter7));
  inv1  gate1087(.a(G1108), .O(gate411inter8));
  nand2 gate1088(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1089(.a(s_77), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1090(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1091(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1092(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1009(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1010(.a(gate415inter0), .b(s_66), .O(gate415inter1));
  and2  gate1011(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1012(.a(s_66), .O(gate415inter3));
  inv1  gate1013(.a(s_67), .O(gate415inter4));
  nand2 gate1014(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1015(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1016(.a(G29), .O(gate415inter7));
  inv1  gate1017(.a(G1120), .O(gate415inter8));
  nand2 gate1018(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1019(.a(s_67), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1020(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1021(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1022(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1149(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1150(.a(gate422inter0), .b(s_86), .O(gate422inter1));
  and2  gate1151(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1152(.a(s_86), .O(gate422inter3));
  inv1  gate1153(.a(s_87), .O(gate422inter4));
  nand2 gate1154(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1155(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1156(.a(G1039), .O(gate422inter7));
  inv1  gate1157(.a(G1135), .O(gate422inter8));
  nand2 gate1158(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1159(.a(s_87), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1160(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1161(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1162(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate953(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate954(.a(gate427inter0), .b(s_58), .O(gate427inter1));
  and2  gate955(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate956(.a(s_58), .O(gate427inter3));
  inv1  gate957(.a(s_59), .O(gate427inter4));
  nand2 gate958(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate959(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate960(.a(G5), .O(gate427inter7));
  inv1  gate961(.a(G1144), .O(gate427inter8));
  nand2 gate962(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate963(.a(s_59), .b(gate427inter3), .O(gate427inter10));
  nor2  gate964(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate965(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate966(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1541(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1542(.a(gate430inter0), .b(s_142), .O(gate430inter1));
  and2  gate1543(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1544(.a(s_142), .O(gate430inter3));
  inv1  gate1545(.a(s_143), .O(gate430inter4));
  nand2 gate1546(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1547(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1548(.a(G1051), .O(gate430inter7));
  inv1  gate1549(.a(G1147), .O(gate430inter8));
  nand2 gate1550(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1551(.a(s_143), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1552(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1553(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1554(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1555(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1556(.a(gate439inter0), .b(s_144), .O(gate439inter1));
  and2  gate1557(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1558(.a(s_144), .O(gate439inter3));
  inv1  gate1559(.a(s_145), .O(gate439inter4));
  nand2 gate1560(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1561(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1562(.a(G11), .O(gate439inter7));
  inv1  gate1563(.a(G1162), .O(gate439inter8));
  nand2 gate1564(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1565(.a(s_145), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1566(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1567(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1568(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1401(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1402(.a(gate444inter0), .b(s_122), .O(gate444inter1));
  and2  gate1403(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1404(.a(s_122), .O(gate444inter3));
  inv1  gate1405(.a(s_123), .O(gate444inter4));
  nand2 gate1406(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1407(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1408(.a(G1072), .O(gate444inter7));
  inv1  gate1409(.a(G1168), .O(gate444inter8));
  nand2 gate1410(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1411(.a(s_123), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1412(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1413(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1414(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1121(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1122(.a(gate446inter0), .b(s_82), .O(gate446inter1));
  and2  gate1123(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1124(.a(s_82), .O(gate446inter3));
  inv1  gate1125(.a(s_83), .O(gate446inter4));
  nand2 gate1126(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1127(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1128(.a(G1075), .O(gate446inter7));
  inv1  gate1129(.a(G1171), .O(gate446inter8));
  nand2 gate1130(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1131(.a(s_83), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1132(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1133(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1134(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1107(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1108(.a(gate448inter0), .b(s_80), .O(gate448inter1));
  and2  gate1109(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1110(.a(s_80), .O(gate448inter3));
  inv1  gate1111(.a(s_81), .O(gate448inter4));
  nand2 gate1112(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1113(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1114(.a(G1078), .O(gate448inter7));
  inv1  gate1115(.a(G1174), .O(gate448inter8));
  nand2 gate1116(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1117(.a(s_81), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1118(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1119(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1120(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1135(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1136(.a(gate456inter0), .b(s_84), .O(gate456inter1));
  and2  gate1137(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1138(.a(s_84), .O(gate456inter3));
  inv1  gate1139(.a(s_85), .O(gate456inter4));
  nand2 gate1140(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1141(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1142(.a(G1090), .O(gate456inter7));
  inv1  gate1143(.a(G1186), .O(gate456inter8));
  nand2 gate1144(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1145(.a(s_85), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1146(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1147(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1148(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1051(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1052(.a(gate457inter0), .b(s_72), .O(gate457inter1));
  and2  gate1053(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1054(.a(s_72), .O(gate457inter3));
  inv1  gate1055(.a(s_73), .O(gate457inter4));
  nand2 gate1056(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1057(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1058(.a(G20), .O(gate457inter7));
  inv1  gate1059(.a(G1189), .O(gate457inter8));
  nand2 gate1060(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1061(.a(s_73), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1062(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1063(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1064(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1527(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1528(.a(gate471inter0), .b(s_140), .O(gate471inter1));
  and2  gate1529(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1530(.a(s_140), .O(gate471inter3));
  inv1  gate1531(.a(s_141), .O(gate471inter4));
  nand2 gate1532(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1533(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1534(.a(G27), .O(gate471inter7));
  inv1  gate1535(.a(G1210), .O(gate471inter8));
  nand2 gate1536(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1537(.a(s_141), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1538(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1539(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1540(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate883(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate884(.a(gate477inter0), .b(s_48), .O(gate477inter1));
  and2  gate885(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate886(.a(s_48), .O(gate477inter3));
  inv1  gate887(.a(s_49), .O(gate477inter4));
  nand2 gate888(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate889(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate890(.a(G30), .O(gate477inter7));
  inv1  gate891(.a(G1219), .O(gate477inter8));
  nand2 gate892(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate893(.a(s_49), .b(gate477inter3), .O(gate477inter10));
  nor2  gate894(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate895(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate896(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1387(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1388(.a(gate478inter0), .b(s_120), .O(gate478inter1));
  and2  gate1389(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1390(.a(s_120), .O(gate478inter3));
  inv1  gate1391(.a(s_121), .O(gate478inter4));
  nand2 gate1392(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1393(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1394(.a(G1123), .O(gate478inter7));
  inv1  gate1395(.a(G1219), .O(gate478inter8));
  nand2 gate1396(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1397(.a(s_121), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1398(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1399(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1400(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1303(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1304(.a(gate487inter0), .b(s_108), .O(gate487inter1));
  and2  gate1305(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1306(.a(s_108), .O(gate487inter3));
  inv1  gate1307(.a(s_109), .O(gate487inter4));
  nand2 gate1308(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1309(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1310(.a(G1236), .O(gate487inter7));
  inv1  gate1311(.a(G1237), .O(gate487inter8));
  nand2 gate1312(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1313(.a(s_109), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1314(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1315(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1316(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1443(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1444(.a(gate495inter0), .b(s_128), .O(gate495inter1));
  and2  gate1445(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1446(.a(s_128), .O(gate495inter3));
  inv1  gate1447(.a(s_129), .O(gate495inter4));
  nand2 gate1448(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1449(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1450(.a(G1252), .O(gate495inter7));
  inv1  gate1451(.a(G1253), .O(gate495inter8));
  nand2 gate1452(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1453(.a(s_129), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1454(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1455(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1456(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate995(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate996(.a(gate501inter0), .b(s_64), .O(gate501inter1));
  and2  gate997(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate998(.a(s_64), .O(gate501inter3));
  inv1  gate999(.a(s_65), .O(gate501inter4));
  nand2 gate1000(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1001(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1002(.a(G1264), .O(gate501inter7));
  inv1  gate1003(.a(G1265), .O(gate501inter8));
  nand2 gate1004(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1005(.a(s_65), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1006(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1007(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1008(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1205(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1206(.a(gate509inter0), .b(s_94), .O(gate509inter1));
  and2  gate1207(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1208(.a(s_94), .O(gate509inter3));
  inv1  gate1209(.a(s_95), .O(gate509inter4));
  nand2 gate1210(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1211(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1212(.a(G1280), .O(gate509inter7));
  inv1  gate1213(.a(G1281), .O(gate509inter8));
  nand2 gate1214(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1215(.a(s_95), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1216(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1217(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1218(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule