module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate693(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate694(.a(gate19inter0), .b(s_76), .O(gate19inter1));
  and2  gate695(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate696(.a(s_76), .O(gate19inter3));
  inv1  gate697(.a(s_77), .O(gate19inter4));
  nand2 gate698(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate699(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate700(.a(N118), .O(gate19inter7));
  inv1  gate701(.a(N4), .O(gate19inter8));
  nand2 gate702(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate703(.a(s_77), .b(gate19inter3), .O(gate19inter10));
  nor2  gate704(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate705(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate706(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate637(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate638(.a(gate20inter0), .b(s_68), .O(gate20inter1));
  and2  gate639(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate640(.a(s_68), .O(gate20inter3));
  inv1  gate641(.a(s_69), .O(gate20inter4));
  nand2 gate642(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate643(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate644(.a(N8), .O(gate20inter7));
  inv1  gate645(.a(N119), .O(gate20inter8));
  nand2 gate646(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate647(.a(s_69), .b(gate20inter3), .O(gate20inter10));
  nor2  gate648(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate649(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate650(.a(gate20inter12), .b(gate20inter1), .O(N157));

  xor2  gate287(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate288(.a(gate21inter0), .b(s_18), .O(gate21inter1));
  and2  gate289(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate290(.a(s_18), .O(gate21inter3));
  inv1  gate291(.a(s_19), .O(gate21inter4));
  nand2 gate292(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate293(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate294(.a(N14), .O(gate21inter7));
  inv1  gate295(.a(N119), .O(gate21inter8));
  nand2 gate296(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate297(.a(s_19), .b(gate21inter3), .O(gate21inter10));
  nor2  gate298(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate299(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate300(.a(gate21inter12), .b(gate21inter1), .O(N158));

  xor2  gate721(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate722(.a(gate22inter0), .b(s_80), .O(gate22inter1));
  and2  gate723(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate724(.a(s_80), .O(gate22inter3));
  inv1  gate725(.a(s_81), .O(gate22inter4));
  nand2 gate726(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate727(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate728(.a(N122), .O(gate22inter7));
  inv1  gate729(.a(N17), .O(gate22inter8));
  nand2 gate730(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate731(.a(s_81), .b(gate22inter3), .O(gate22inter10));
  nor2  gate732(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate733(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate734(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );

  xor2  gate231(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate232(.a(gate25inter0), .b(s_10), .O(gate25inter1));
  and2  gate233(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate234(.a(s_10), .O(gate25inter3));
  inv1  gate235(.a(s_11), .O(gate25inter4));
  nand2 gate236(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate237(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate238(.a(N134), .O(gate25inter7));
  inv1  gate239(.a(N56), .O(gate25inter8));
  nand2 gate240(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate241(.a(s_11), .b(gate25inter3), .O(gate25inter10));
  nor2  gate242(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate243(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate244(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate651(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate652(.a(gate27inter0), .b(s_70), .O(gate27inter1));
  and2  gate653(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate654(.a(s_70), .O(gate27inter3));
  inv1  gate655(.a(s_71), .O(gate27inter4));
  nand2 gate656(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate657(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate658(.a(N142), .O(gate27inter7));
  inv1  gate659(.a(N82), .O(gate27inter8));
  nand2 gate660(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate661(.a(s_71), .b(gate27inter3), .O(gate27inter10));
  nor2  gate662(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate663(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate664(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate343(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate344(.a(gate30inter0), .b(s_26), .O(gate30inter1));
  and2  gate345(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate346(.a(s_26), .O(gate30inter3));
  inv1  gate347(.a(s_27), .O(gate30inter4));
  nand2 gate348(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate349(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate350(.a(N21), .O(gate30inter7));
  inv1  gate351(.a(N123), .O(gate30inter8));
  nand2 gate352(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate353(.a(s_27), .b(gate30inter3), .O(gate30inter10));
  nor2  gate354(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate355(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate356(.a(gate30inter12), .b(gate30inter1), .O(N183));

  xor2  gate483(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate484(.a(gate31inter0), .b(s_46), .O(gate31inter1));
  and2  gate485(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate486(.a(s_46), .O(gate31inter3));
  inv1  gate487(.a(s_47), .O(gate31inter4));
  nand2 gate488(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate489(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate490(.a(N27), .O(gate31inter7));
  inv1  gate491(.a(N123), .O(gate31inter8));
  nand2 gate492(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate493(.a(s_47), .b(gate31inter3), .O(gate31inter10));
  nor2  gate494(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate495(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate496(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );

  xor2  gate511(.a(N127), .b(N40), .O(gate33inter0));
  nand2 gate512(.a(gate33inter0), .b(s_50), .O(gate33inter1));
  and2  gate513(.a(N127), .b(N40), .O(gate33inter2));
  inv1  gate514(.a(s_50), .O(gate33inter3));
  inv1  gate515(.a(s_51), .O(gate33inter4));
  nand2 gate516(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate517(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate518(.a(N40), .O(gate33inter7));
  inv1  gate519(.a(N127), .O(gate33inter8));
  nand2 gate520(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate521(.a(s_51), .b(gate33inter3), .O(gate33inter10));
  nor2  gate522(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate523(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate524(.a(gate33inter12), .b(gate33inter1), .O(N186));

  xor2  gate371(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate372(.a(gate34inter0), .b(s_30), .O(gate34inter1));
  and2  gate373(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate374(.a(s_30), .O(gate34inter3));
  inv1  gate375(.a(s_31), .O(gate34inter4));
  nand2 gate376(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate377(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate378(.a(N47), .O(gate34inter7));
  inv1  gate379(.a(N131), .O(gate34inter8));
  nand2 gate380(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate381(.a(s_31), .b(gate34inter3), .O(gate34inter10));
  nor2  gate382(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate383(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate384(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate203(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate204(.a(gate35inter0), .b(s_6), .O(gate35inter1));
  and2  gate205(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate206(.a(s_6), .O(gate35inter3));
  inv1  gate207(.a(s_7), .O(gate35inter4));
  nand2 gate208(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate209(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate210(.a(N53), .O(gate35inter7));
  inv1  gate211(.a(N131), .O(gate35inter8));
  nand2 gate212(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate213(.a(s_7), .b(gate35inter3), .O(gate35inter10));
  nor2  gate214(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate215(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate216(.a(gate35inter12), .b(gate35inter1), .O(N188));

  xor2  gate623(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate624(.a(gate36inter0), .b(s_66), .O(gate36inter1));
  and2  gate625(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate626(.a(s_66), .O(gate36inter3));
  inv1  gate627(.a(s_67), .O(gate36inter4));
  nand2 gate628(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate629(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate630(.a(N60), .O(gate36inter7));
  inv1  gate631(.a(N135), .O(gate36inter8));
  nand2 gate632(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate633(.a(s_67), .b(gate36inter3), .O(gate36inter10));
  nor2  gate634(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate635(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate636(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate161(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate162(.a(gate41inter0), .b(s_0), .O(gate41inter1));
  and2  gate163(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate164(.a(s_0), .O(gate41inter3));
  inv1  gate165(.a(s_1), .O(gate41inter4));
  nand2 gate166(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate167(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate168(.a(N92), .O(gate41inter7));
  inv1  gate169(.a(N143), .O(gate41inter8));
  nand2 gate170(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate171(.a(s_1), .b(gate41inter3), .O(gate41inter10));
  nor2  gate172(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate173(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate174(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate357(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate358(.a(gate43inter0), .b(s_28), .O(gate43inter1));
  and2  gate359(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate360(.a(s_28), .O(gate43inter3));
  inv1  gate361(.a(s_29), .O(gate43inter4));
  nand2 gate362(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate363(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate364(.a(N105), .O(gate43inter7));
  inv1  gate365(.a(N147), .O(gate43inter8));
  nand2 gate366(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate367(.a(s_29), .b(gate43inter3), .O(gate43inter10));
  nor2  gate368(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate369(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate370(.a(gate43inter12), .b(gate43inter1), .O(N196));

  xor2  gate455(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate456(.a(gate44inter0), .b(s_42), .O(gate44inter1));
  and2  gate457(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate458(.a(s_42), .O(gate44inter3));
  inv1  gate459(.a(s_43), .O(gate44inter4));
  nand2 gate460(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate461(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate462(.a(N112), .O(gate44inter7));
  inv1  gate463(.a(N151), .O(gate44inter8));
  nand2 gate464(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate465(.a(s_43), .b(gate44inter3), .O(gate44inter10));
  nor2  gate466(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate467(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate468(.a(gate44inter12), .b(gate44inter1), .O(N197));
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate175(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate176(.a(gate52inter0), .b(s_2), .O(gate52inter1));
  and2  gate177(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate178(.a(s_2), .O(gate52inter3));
  inv1  gate179(.a(s_3), .O(gate52inter4));
  nand2 gate180(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate181(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate182(.a(N203), .O(gate52inter7));
  inv1  gate183(.a(N162), .O(gate52inter8));
  nand2 gate184(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate185(.a(s_3), .b(gate52inter3), .O(gate52inter10));
  nor2  gate186(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate187(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate188(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate245(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate246(.a(gate59inter0), .b(s_12), .O(gate59inter1));
  and2  gate247(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate248(.a(s_12), .O(gate59inter3));
  inv1  gate249(.a(s_13), .O(gate59inter4));
  nand2 gate250(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate251(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate252(.a(N203), .O(gate59inter7));
  inv1  gate253(.a(N177), .O(gate59inter8));
  nand2 gate254(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate255(.a(s_13), .b(gate59inter3), .O(gate59inter10));
  nor2  gate256(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate257(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate258(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate497(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate498(.a(gate62inter0), .b(s_48), .O(gate62inter1));
  and2  gate499(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate500(.a(s_48), .O(gate62inter3));
  inv1  gate501(.a(s_49), .O(gate62inter4));
  nand2 gate502(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate503(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate504(.a(N213), .O(gate62inter7));
  inv1  gate505(.a(N37), .O(gate62inter8));
  nand2 gate506(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate507(.a(s_49), .b(gate62inter3), .O(gate62inter10));
  nor2  gate508(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate509(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate510(.a(gate62inter12), .b(gate62inter1), .O(N254));
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );

  xor2  gate581(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate582(.a(gate66inter0), .b(s_60), .O(gate66inter1));
  and2  gate583(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate584(.a(s_60), .O(gate66inter3));
  inv1  gate585(.a(s_61), .O(gate66inter4));
  nand2 gate586(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate587(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate588(.a(N213), .O(gate66inter7));
  inv1  gate589(.a(N89), .O(gate66inter8));
  nand2 gate590(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate591(.a(s_61), .b(gate66inter3), .O(gate66inter10));
  nor2  gate592(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate593(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate594(.a(gate66inter12), .b(gate66inter1), .O(N258));

  xor2  gate301(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate302(.a(gate67inter0), .b(s_20), .O(gate67inter1));
  and2  gate303(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate304(.a(s_20), .O(gate67inter3));
  inv1  gate305(.a(s_21), .O(gate67inter4));
  nand2 gate306(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate307(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate308(.a(N213), .O(gate67inter7));
  inv1  gate309(.a(N102), .O(gate67inter8));
  nand2 gate310(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate311(.a(s_21), .b(gate67inter3), .O(gate67inter10));
  nor2  gate312(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate313(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate314(.a(gate67inter12), .b(gate67inter1), .O(N259));
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate399(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate400(.a(gate71inter0), .b(s_34), .O(gate71inter1));
  and2  gate401(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate402(.a(s_34), .O(gate71inter3));
  inv1  gate403(.a(s_35), .O(gate71inter4));
  nand2 gate404(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate405(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate406(.a(N230), .O(gate71inter7));
  inv1  gate407(.a(N185), .O(gate71inter8));
  nand2 gate408(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate409(.a(s_35), .b(gate71inter3), .O(gate71inter10));
  nor2  gate410(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate411(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate412(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );

  xor2  gate427(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate428(.a(gate74inter0), .b(s_38), .O(gate74inter1));
  and2  gate429(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate430(.a(s_38), .O(gate74inter3));
  inv1  gate431(.a(s_39), .O(gate74inter4));
  nand2 gate432(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate433(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate434(.a(N239), .O(gate74inter7));
  inv1  gate435(.a(N191), .O(gate74inter8));
  nand2 gate436(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate437(.a(s_39), .b(gate74inter3), .O(gate74inter10));
  nor2  gate438(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate439(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate440(.a(gate74inter12), .b(gate74inter1), .O(N276));

  xor2  gate259(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate260(.a(gate75inter0), .b(s_14), .O(gate75inter1));
  and2  gate261(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate262(.a(s_14), .O(gate75inter3));
  inv1  gate263(.a(s_15), .O(gate75inter4));
  nand2 gate264(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate265(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate266(.a(N243), .O(gate75inter7));
  inv1  gate267(.a(N193), .O(gate75inter8));
  nand2 gate268(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate269(.a(s_15), .b(gate75inter3), .O(gate75inter10));
  nor2  gate270(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate271(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate272(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate539(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate540(.a(gate78inter0), .b(s_54), .O(gate78inter1));
  and2  gate541(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate542(.a(s_54), .O(gate78inter3));
  inv1  gate543(.a(s_55), .O(gate78inter4));
  nand2 gate544(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate545(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate546(.a(N227), .O(gate78inter7));
  inv1  gate547(.a(N184), .O(gate78inter8));
  nand2 gate548(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate549(.a(s_55), .b(gate78inter3), .O(gate78inter10));
  nor2  gate550(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate551(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate552(.a(gate78inter12), .b(gate78inter1), .O(N288));

  xor2  gate609(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate610(.a(gate79inter0), .b(s_64), .O(gate79inter1));
  and2  gate611(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate612(.a(s_64), .O(gate79inter3));
  inv1  gate613(.a(s_65), .O(gate79inter4));
  nand2 gate614(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate615(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate616(.a(N230), .O(gate79inter7));
  inv1  gate617(.a(N186), .O(gate79inter8));
  nand2 gate618(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate619(.a(s_65), .b(gate79inter3), .O(gate79inter10));
  nor2  gate620(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate621(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate622(.a(gate79inter12), .b(gate79inter1), .O(N289));
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );

  xor2  gate385(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate386(.a(gate85inter0), .b(s_32), .O(gate85inter1));
  and2  gate387(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate388(.a(s_32), .O(gate85inter3));
  inv1  gate389(.a(s_33), .O(gate85inter4));
  nand2 gate390(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate391(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate392(.a(N251), .O(gate85inter7));
  inv1  gate393(.a(N198), .O(gate85inter8));
  nand2 gate394(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate395(.a(s_33), .b(gate85inter3), .O(gate85inter10));
  nor2  gate396(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate397(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate398(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );

  xor2  gate553(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate554(.a(gate102inter0), .b(s_56), .O(gate102inter1));
  and2  gate555(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate556(.a(s_56), .O(gate102inter3));
  inv1  gate557(.a(s_57), .O(gate102inter4));
  nand2 gate558(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate559(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate560(.a(N309), .O(gate102inter7));
  inv1  gate561(.a(N270), .O(gate102inter8));
  nand2 gate562(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate563(.a(s_57), .b(gate102inter3), .O(gate102inter10));
  nor2  gate564(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate565(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate566(.a(gate102inter12), .b(gate102inter1), .O(N333));

  xor2  gate189(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate190(.a(gate103inter0), .b(s_4), .O(gate103inter1));
  and2  gate191(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate192(.a(s_4), .O(gate103inter3));
  inv1  gate193(.a(s_5), .O(gate103inter4));
  nand2 gate194(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate195(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate196(.a(N8), .O(gate103inter7));
  inv1  gate197(.a(N319), .O(gate103inter8));
  nand2 gate198(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate199(.a(s_5), .b(gate103inter3), .O(gate103inter10));
  nor2  gate200(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate201(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate202(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate217(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate218(.a(gate105inter0), .b(s_8), .O(gate105inter1));
  and2  gate219(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate220(.a(s_8), .O(gate105inter3));
  inv1  gate221(.a(s_9), .O(gate105inter4));
  nand2 gate222(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate223(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate224(.a(N319), .O(gate105inter7));
  inv1  gate225(.a(N21), .O(gate105inter8));
  nand2 gate226(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate227(.a(s_9), .b(gate105inter3), .O(gate105inter10));
  nor2  gate228(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate229(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate230(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );

  xor2  gate441(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate442(.a(gate112inter0), .b(s_40), .O(gate112inter1));
  and2  gate443(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate444(.a(s_40), .O(gate112inter3));
  inv1  gate445(.a(s_41), .O(gate112inter4));
  nand2 gate446(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate447(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate448(.a(N309), .O(gate112inter7));
  inv1  gate449(.a(N285), .O(gate112inter8));
  nand2 gate450(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate451(.a(s_41), .b(gate112inter3), .O(gate112inter10));
  nor2  gate452(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate453(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate454(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate525(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate526(.a(gate115inter0), .b(s_52), .O(gate115inter1));
  and2  gate527(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate528(.a(s_52), .O(gate115inter3));
  inv1  gate529(.a(s_53), .O(gate115inter4));
  nand2 gate530(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate531(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate532(.a(N319), .O(gate115inter7));
  inv1  gate533(.a(N99), .O(gate115inter8));
  nand2 gate534(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate535(.a(s_53), .b(gate115inter3), .O(gate115inter10));
  nor2  gate536(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate537(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate538(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate567(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate568(.a(gate120inter0), .b(s_58), .O(gate120inter1));
  and2  gate569(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate570(.a(s_58), .O(gate120inter3));
  inv1  gate571(.a(s_59), .O(gate120inter4));
  nand2 gate572(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate573(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate574(.a(N333), .O(gate120inter7));
  inv1  gate575(.a(N303), .O(gate120inter8));
  nand2 gate576(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate577(.a(s_59), .b(gate120inter3), .O(gate120inter10));
  nor2  gate578(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate579(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate580(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );

  xor2  gate679(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate680(.a(gate122inter0), .b(s_74), .O(gate122inter1));
  and2  gate681(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate682(.a(s_74), .O(gate122inter3));
  inv1  gate683(.a(s_75), .O(gate122inter4));
  nand2 gate684(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate685(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate686(.a(N337), .O(gate122inter7));
  inv1  gate687(.a(N305), .O(gate122inter8));
  nand2 gate688(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate689(.a(s_75), .b(gate122inter3), .O(gate122inter10));
  nor2  gate690(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate691(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate692(.a(gate122inter12), .b(gate122inter1), .O(N353));

  xor2  gate469(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate470(.a(gate123inter0), .b(s_44), .O(gate123inter1));
  and2  gate471(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate472(.a(s_44), .O(gate123inter3));
  inv1  gate473(.a(s_45), .O(gate123inter4));
  nand2 gate474(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate475(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate476(.a(N339), .O(gate123inter7));
  inv1  gate477(.a(N306), .O(gate123inter8));
  nand2 gate478(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate479(.a(s_45), .b(gate123inter3), .O(gate123inter10));
  nor2  gate480(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate481(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate482(.a(gate123inter12), .b(gate123inter1), .O(N354));
nand2 gate124( .a(N341), .b(N307), .O(N355) );

  xor2  gate315(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate316(.a(gate125inter0), .b(s_22), .O(gate125inter1));
  and2  gate317(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate318(.a(s_22), .O(gate125inter3));
  inv1  gate319(.a(s_23), .O(gate125inter4));
  nand2 gate320(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate321(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate322(.a(N343), .O(gate125inter7));
  inv1  gate323(.a(N308), .O(gate125inter8));
  nand2 gate324(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate325(.a(s_23), .b(gate125inter3), .O(gate125inter10));
  nor2  gate326(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate327(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate328(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate329(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate330(.a(gate129inter0), .b(s_24), .O(gate129inter1));
  and2  gate331(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate332(.a(s_24), .O(gate129inter3));
  inv1  gate333(.a(s_25), .O(gate129inter4));
  nand2 gate334(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate335(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate336(.a(N14), .O(gate129inter7));
  inv1  gate337(.a(N360), .O(gate129inter8));
  nand2 gate338(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate339(.a(s_25), .b(gate129inter3), .O(gate129inter10));
  nor2  gate340(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate341(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate342(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate273(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate274(.a(gate131inter0), .b(s_16), .O(gate131inter1));
  and2  gate275(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate276(.a(s_16), .O(gate131inter3));
  inv1  gate277(.a(s_17), .O(gate131inter4));
  nand2 gate278(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate279(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate280(.a(N360), .O(gate131inter7));
  inv1  gate281(.a(N40), .O(gate131inter8));
  nand2 gate282(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate283(.a(s_17), .b(gate131inter3), .O(gate131inter10));
  nor2  gate284(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate285(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate286(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );

  xor2  gate665(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate666(.a(gate134inter0), .b(s_72), .O(gate134inter1));
  and2  gate667(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate668(.a(s_72), .O(gate134inter3));
  inv1  gate669(.a(s_73), .O(gate134inter4));
  nand2 gate670(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate671(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate672(.a(N360), .O(gate134inter7));
  inv1  gate673(.a(N79), .O(gate134inter8));
  nand2 gate674(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate675(.a(s_73), .b(gate134inter3), .O(gate134inter10));
  nor2  gate676(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate677(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate678(.a(gate134inter12), .b(gate134inter1), .O(N376));

  xor2  gate595(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate596(.a(gate135inter0), .b(s_62), .O(gate135inter1));
  and2  gate597(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate598(.a(s_62), .O(gate135inter3));
  inv1  gate599(.a(s_63), .O(gate135inter4));
  nand2 gate600(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate601(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate602(.a(N360), .O(gate135inter7));
  inv1  gate603(.a(N92), .O(gate135inter8));
  nand2 gate604(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate605(.a(s_63), .b(gate135inter3), .O(gate135inter10));
  nor2  gate606(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate607(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate608(.a(gate135inter12), .b(gate135inter1), .O(N377));

  xor2  gate413(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate414(.a(gate136inter0), .b(s_36), .O(gate136inter1));
  and2  gate415(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate416(.a(s_36), .O(gate136inter3));
  inv1  gate417(.a(s_37), .O(gate136inter4));
  nand2 gate418(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate419(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate420(.a(N360), .O(gate136inter7));
  inv1  gate421(.a(N105), .O(gate136inter8));
  nand2 gate422(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate423(.a(s_37), .b(gate136inter3), .O(gate136inter10));
  nor2  gate424(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate425(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate426(.a(gate136inter12), .b(gate136inter1), .O(N378));

  xor2  gate707(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate708(.a(gate137inter0), .b(s_78), .O(gate137inter1));
  and2  gate709(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate710(.a(s_78), .O(gate137inter3));
  inv1  gate711(.a(s_79), .O(gate137inter4));
  nand2 gate712(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate713(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate714(.a(N360), .O(gate137inter7));
  inv1  gate715(.a(N115), .O(gate137inter8));
  nand2 gate716(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate717(.a(s_79), .b(gate137inter3), .O(gate137inter10));
  nor2  gate718(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate719(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate720(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule