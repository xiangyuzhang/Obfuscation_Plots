module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1541(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1542(.a(gate9inter0), .b(s_142), .O(gate9inter1));
  and2  gate1543(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1544(.a(s_142), .O(gate9inter3));
  inv1  gate1545(.a(s_143), .O(gate9inter4));
  nand2 gate1546(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1547(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1548(.a(G1), .O(gate9inter7));
  inv1  gate1549(.a(G2), .O(gate9inter8));
  nand2 gate1550(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1551(.a(s_143), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1552(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1553(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1554(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1093(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1094(.a(gate11inter0), .b(s_78), .O(gate11inter1));
  and2  gate1095(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1096(.a(s_78), .O(gate11inter3));
  inv1  gate1097(.a(s_79), .O(gate11inter4));
  nand2 gate1098(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1099(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1100(.a(G5), .O(gate11inter7));
  inv1  gate1101(.a(G6), .O(gate11inter8));
  nand2 gate1102(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1103(.a(s_79), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1104(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1105(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1106(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1415(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1416(.a(gate13inter0), .b(s_124), .O(gate13inter1));
  and2  gate1417(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1418(.a(s_124), .O(gate13inter3));
  inv1  gate1419(.a(s_125), .O(gate13inter4));
  nand2 gate1420(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1421(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1422(.a(G9), .O(gate13inter7));
  inv1  gate1423(.a(G10), .O(gate13inter8));
  nand2 gate1424(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1425(.a(s_125), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1426(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1427(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1428(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate673(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate674(.a(gate15inter0), .b(s_18), .O(gate15inter1));
  and2  gate675(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate676(.a(s_18), .O(gate15inter3));
  inv1  gate677(.a(s_19), .O(gate15inter4));
  nand2 gate678(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate679(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate680(.a(G13), .O(gate15inter7));
  inv1  gate681(.a(G14), .O(gate15inter8));
  nand2 gate682(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate683(.a(s_19), .b(gate15inter3), .O(gate15inter10));
  nor2  gate684(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate685(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate686(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate729(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate730(.a(gate22inter0), .b(s_26), .O(gate22inter1));
  and2  gate731(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate732(.a(s_26), .O(gate22inter3));
  inv1  gate733(.a(s_27), .O(gate22inter4));
  nand2 gate734(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate735(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate736(.a(G27), .O(gate22inter7));
  inv1  gate737(.a(G28), .O(gate22inter8));
  nand2 gate738(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate739(.a(s_27), .b(gate22inter3), .O(gate22inter10));
  nor2  gate740(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate741(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate742(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1555(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1556(.a(gate26inter0), .b(s_144), .O(gate26inter1));
  and2  gate1557(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1558(.a(s_144), .O(gate26inter3));
  inv1  gate1559(.a(s_145), .O(gate26inter4));
  nand2 gate1560(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1561(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1562(.a(G9), .O(gate26inter7));
  inv1  gate1563(.a(G13), .O(gate26inter8));
  nand2 gate1564(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1565(.a(s_145), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1566(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1567(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1568(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate799(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate800(.a(gate32inter0), .b(s_36), .O(gate32inter1));
  and2  gate801(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate802(.a(s_36), .O(gate32inter3));
  inv1  gate803(.a(s_37), .O(gate32inter4));
  nand2 gate804(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate805(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate806(.a(G12), .O(gate32inter7));
  inv1  gate807(.a(G16), .O(gate32inter8));
  nand2 gate808(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate809(.a(s_37), .b(gate32inter3), .O(gate32inter10));
  nor2  gate810(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate811(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate812(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1023(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1024(.a(gate35inter0), .b(s_68), .O(gate35inter1));
  and2  gate1025(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1026(.a(s_68), .O(gate35inter3));
  inv1  gate1027(.a(s_69), .O(gate35inter4));
  nand2 gate1028(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1029(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1030(.a(G18), .O(gate35inter7));
  inv1  gate1031(.a(G22), .O(gate35inter8));
  nand2 gate1032(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1033(.a(s_69), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1034(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1035(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1036(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1457(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1458(.a(gate42inter0), .b(s_130), .O(gate42inter1));
  and2  gate1459(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1460(.a(s_130), .O(gate42inter3));
  inv1  gate1461(.a(s_131), .O(gate42inter4));
  nand2 gate1462(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1463(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1464(.a(G2), .O(gate42inter7));
  inv1  gate1465(.a(G266), .O(gate42inter8));
  nand2 gate1466(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1467(.a(s_131), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1468(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1469(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1470(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate813(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate814(.a(gate43inter0), .b(s_38), .O(gate43inter1));
  and2  gate815(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate816(.a(s_38), .O(gate43inter3));
  inv1  gate817(.a(s_39), .O(gate43inter4));
  nand2 gate818(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate819(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate820(.a(G3), .O(gate43inter7));
  inv1  gate821(.a(G269), .O(gate43inter8));
  nand2 gate822(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate823(.a(s_39), .b(gate43inter3), .O(gate43inter10));
  nor2  gate824(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate825(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate826(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate911(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate912(.a(gate57inter0), .b(s_52), .O(gate57inter1));
  and2  gate913(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate914(.a(s_52), .O(gate57inter3));
  inv1  gate915(.a(s_53), .O(gate57inter4));
  nand2 gate916(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate917(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate918(.a(G17), .O(gate57inter7));
  inv1  gate919(.a(G290), .O(gate57inter8));
  nand2 gate920(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate921(.a(s_53), .b(gate57inter3), .O(gate57inter10));
  nor2  gate922(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate923(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate924(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1191(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1192(.a(gate59inter0), .b(s_92), .O(gate59inter1));
  and2  gate1193(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1194(.a(s_92), .O(gate59inter3));
  inv1  gate1195(.a(s_93), .O(gate59inter4));
  nand2 gate1196(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1197(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1198(.a(G19), .O(gate59inter7));
  inv1  gate1199(.a(G293), .O(gate59inter8));
  nand2 gate1200(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1201(.a(s_93), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1202(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1203(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1204(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate953(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate954(.a(gate62inter0), .b(s_58), .O(gate62inter1));
  and2  gate955(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate956(.a(s_58), .O(gate62inter3));
  inv1  gate957(.a(s_59), .O(gate62inter4));
  nand2 gate958(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate959(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate960(.a(G22), .O(gate62inter7));
  inv1  gate961(.a(G296), .O(gate62inter8));
  nand2 gate962(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate963(.a(s_59), .b(gate62inter3), .O(gate62inter10));
  nor2  gate964(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate965(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate966(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate967(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate968(.a(gate64inter0), .b(s_60), .O(gate64inter1));
  and2  gate969(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate970(.a(s_60), .O(gate64inter3));
  inv1  gate971(.a(s_61), .O(gate64inter4));
  nand2 gate972(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate973(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate974(.a(G24), .O(gate64inter7));
  inv1  gate975(.a(G299), .O(gate64inter8));
  nand2 gate976(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate977(.a(s_61), .b(gate64inter3), .O(gate64inter10));
  nor2  gate978(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate979(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate980(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1443(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1444(.a(gate68inter0), .b(s_128), .O(gate68inter1));
  and2  gate1445(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1446(.a(s_128), .O(gate68inter3));
  inv1  gate1447(.a(s_129), .O(gate68inter4));
  nand2 gate1448(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1449(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1450(.a(G28), .O(gate68inter7));
  inv1  gate1451(.a(G305), .O(gate68inter8));
  nand2 gate1452(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1453(.a(s_129), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1454(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1455(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1456(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1569(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1570(.a(gate74inter0), .b(s_146), .O(gate74inter1));
  and2  gate1571(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1572(.a(s_146), .O(gate74inter3));
  inv1  gate1573(.a(s_147), .O(gate74inter4));
  nand2 gate1574(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1575(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1576(.a(G5), .O(gate74inter7));
  inv1  gate1577(.a(G314), .O(gate74inter8));
  nand2 gate1578(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1579(.a(s_147), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1580(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1581(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1582(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1583(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1584(.a(gate78inter0), .b(s_148), .O(gate78inter1));
  and2  gate1585(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1586(.a(s_148), .O(gate78inter3));
  inv1  gate1587(.a(s_149), .O(gate78inter4));
  nand2 gate1588(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1589(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1590(.a(G6), .O(gate78inter7));
  inv1  gate1591(.a(G320), .O(gate78inter8));
  nand2 gate1592(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1593(.a(s_149), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1594(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1595(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1596(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate743(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate744(.a(gate80inter0), .b(s_28), .O(gate80inter1));
  and2  gate745(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate746(.a(s_28), .O(gate80inter3));
  inv1  gate747(.a(s_29), .O(gate80inter4));
  nand2 gate748(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate749(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate750(.a(G14), .O(gate80inter7));
  inv1  gate751(.a(G323), .O(gate80inter8));
  nand2 gate752(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate753(.a(s_29), .b(gate80inter3), .O(gate80inter10));
  nor2  gate754(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate755(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate756(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1079(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1080(.a(gate81inter0), .b(s_76), .O(gate81inter1));
  and2  gate1081(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1082(.a(s_76), .O(gate81inter3));
  inv1  gate1083(.a(s_77), .O(gate81inter4));
  nand2 gate1084(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1085(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1086(.a(G3), .O(gate81inter7));
  inv1  gate1087(.a(G326), .O(gate81inter8));
  nand2 gate1088(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1089(.a(s_77), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1090(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1091(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1092(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1345(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1346(.a(gate88inter0), .b(s_114), .O(gate88inter1));
  and2  gate1347(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1348(.a(s_114), .O(gate88inter3));
  inv1  gate1349(.a(s_115), .O(gate88inter4));
  nand2 gate1350(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1351(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1352(.a(G16), .O(gate88inter7));
  inv1  gate1353(.a(G335), .O(gate88inter8));
  nand2 gate1354(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1355(.a(s_115), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1356(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1357(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1358(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate687(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate688(.a(gate94inter0), .b(s_20), .O(gate94inter1));
  and2  gate689(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate690(.a(s_20), .O(gate94inter3));
  inv1  gate691(.a(s_21), .O(gate94inter4));
  nand2 gate692(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate693(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate694(.a(G22), .O(gate94inter7));
  inv1  gate695(.a(G344), .O(gate94inter8));
  nand2 gate696(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate697(.a(s_21), .b(gate94inter3), .O(gate94inter10));
  nor2  gate698(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate699(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate700(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate631(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate632(.a(gate96inter0), .b(s_12), .O(gate96inter1));
  and2  gate633(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate634(.a(s_12), .O(gate96inter3));
  inv1  gate635(.a(s_13), .O(gate96inter4));
  nand2 gate636(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate637(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate638(.a(G30), .O(gate96inter7));
  inv1  gate639(.a(G347), .O(gate96inter8));
  nand2 gate640(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate641(.a(s_13), .b(gate96inter3), .O(gate96inter10));
  nor2  gate642(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate643(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate644(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate645(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate646(.a(gate102inter0), .b(s_14), .O(gate102inter1));
  and2  gate647(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate648(.a(s_14), .O(gate102inter3));
  inv1  gate649(.a(s_15), .O(gate102inter4));
  nand2 gate650(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate651(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate652(.a(G24), .O(gate102inter7));
  inv1  gate653(.a(G356), .O(gate102inter8));
  nand2 gate654(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate655(.a(s_15), .b(gate102inter3), .O(gate102inter10));
  nor2  gate656(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate657(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate658(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate715(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate716(.a(gate109inter0), .b(s_24), .O(gate109inter1));
  and2  gate717(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate718(.a(s_24), .O(gate109inter3));
  inv1  gate719(.a(s_25), .O(gate109inter4));
  nand2 gate720(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate721(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate722(.a(G370), .O(gate109inter7));
  inv1  gate723(.a(G371), .O(gate109inter8));
  nand2 gate724(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate725(.a(s_25), .b(gate109inter3), .O(gate109inter10));
  nor2  gate726(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate727(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate728(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1177(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1178(.a(gate117inter0), .b(s_90), .O(gate117inter1));
  and2  gate1179(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1180(.a(s_90), .O(gate117inter3));
  inv1  gate1181(.a(s_91), .O(gate117inter4));
  nand2 gate1182(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1183(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1184(.a(G386), .O(gate117inter7));
  inv1  gate1185(.a(G387), .O(gate117inter8));
  nand2 gate1186(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1187(.a(s_91), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1188(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1189(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1190(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate981(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate982(.a(gate125inter0), .b(s_62), .O(gate125inter1));
  and2  gate983(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate984(.a(s_62), .O(gate125inter3));
  inv1  gate985(.a(s_63), .O(gate125inter4));
  nand2 gate986(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate987(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate988(.a(G402), .O(gate125inter7));
  inv1  gate989(.a(G403), .O(gate125inter8));
  nand2 gate990(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate991(.a(s_63), .b(gate125inter3), .O(gate125inter10));
  nor2  gate992(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate993(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate994(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1331(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1332(.a(gate135inter0), .b(s_112), .O(gate135inter1));
  and2  gate1333(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1334(.a(s_112), .O(gate135inter3));
  inv1  gate1335(.a(s_113), .O(gate135inter4));
  nand2 gate1336(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1337(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1338(.a(G422), .O(gate135inter7));
  inv1  gate1339(.a(G423), .O(gate135inter8));
  nand2 gate1340(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1341(.a(s_113), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1342(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1343(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1344(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate575(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate576(.a(gate138inter0), .b(s_4), .O(gate138inter1));
  and2  gate577(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate578(.a(s_4), .O(gate138inter3));
  inv1  gate579(.a(s_5), .O(gate138inter4));
  nand2 gate580(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate581(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate582(.a(G432), .O(gate138inter7));
  inv1  gate583(.a(G435), .O(gate138inter8));
  nand2 gate584(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate585(.a(s_5), .b(gate138inter3), .O(gate138inter10));
  nor2  gate586(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate587(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate588(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1065(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1066(.a(gate139inter0), .b(s_74), .O(gate139inter1));
  and2  gate1067(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1068(.a(s_74), .O(gate139inter3));
  inv1  gate1069(.a(s_75), .O(gate139inter4));
  nand2 gate1070(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1071(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1072(.a(G438), .O(gate139inter7));
  inv1  gate1073(.a(G441), .O(gate139inter8));
  nand2 gate1074(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1075(.a(s_75), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1076(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1077(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1078(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1275(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1276(.a(gate143inter0), .b(s_104), .O(gate143inter1));
  and2  gate1277(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1278(.a(s_104), .O(gate143inter3));
  inv1  gate1279(.a(s_105), .O(gate143inter4));
  nand2 gate1280(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1281(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1282(.a(G462), .O(gate143inter7));
  inv1  gate1283(.a(G465), .O(gate143inter8));
  nand2 gate1284(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1285(.a(s_105), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1286(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1287(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1288(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1317(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1318(.a(gate154inter0), .b(s_110), .O(gate154inter1));
  and2  gate1319(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1320(.a(s_110), .O(gate154inter3));
  inv1  gate1321(.a(s_111), .O(gate154inter4));
  nand2 gate1322(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1323(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1324(.a(G429), .O(gate154inter7));
  inv1  gate1325(.a(G522), .O(gate154inter8));
  nand2 gate1326(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1327(.a(s_111), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1328(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1329(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1330(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1387(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1388(.a(gate158inter0), .b(s_120), .O(gate158inter1));
  and2  gate1389(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1390(.a(s_120), .O(gate158inter3));
  inv1  gate1391(.a(s_121), .O(gate158inter4));
  nand2 gate1392(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1393(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1394(.a(G441), .O(gate158inter7));
  inv1  gate1395(.a(G528), .O(gate158inter8));
  nand2 gate1396(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1397(.a(s_121), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1398(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1399(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1400(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1163(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1164(.a(gate162inter0), .b(s_88), .O(gate162inter1));
  and2  gate1165(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1166(.a(s_88), .O(gate162inter3));
  inv1  gate1167(.a(s_89), .O(gate162inter4));
  nand2 gate1168(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1169(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1170(.a(G453), .O(gate162inter7));
  inv1  gate1171(.a(G534), .O(gate162inter8));
  nand2 gate1172(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1173(.a(s_89), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1174(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1175(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1176(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1499(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1500(.a(gate164inter0), .b(s_136), .O(gate164inter1));
  and2  gate1501(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1502(.a(s_136), .O(gate164inter3));
  inv1  gate1503(.a(s_137), .O(gate164inter4));
  nand2 gate1504(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1505(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1506(.a(G459), .O(gate164inter7));
  inv1  gate1507(.a(G537), .O(gate164inter8));
  nand2 gate1508(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1509(.a(s_137), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1510(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1511(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1512(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1205(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1206(.a(gate171inter0), .b(s_94), .O(gate171inter1));
  and2  gate1207(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1208(.a(s_94), .O(gate171inter3));
  inv1  gate1209(.a(s_95), .O(gate171inter4));
  nand2 gate1210(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1211(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1212(.a(G480), .O(gate171inter7));
  inv1  gate1213(.a(G549), .O(gate171inter8));
  nand2 gate1214(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1215(.a(s_95), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1216(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1217(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1218(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate547(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate548(.a(gate174inter0), .b(s_0), .O(gate174inter1));
  and2  gate549(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate550(.a(s_0), .O(gate174inter3));
  inv1  gate551(.a(s_1), .O(gate174inter4));
  nand2 gate552(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate553(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate554(.a(G489), .O(gate174inter7));
  inv1  gate555(.a(G552), .O(gate174inter8));
  nand2 gate556(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate557(.a(s_1), .b(gate174inter3), .O(gate174inter10));
  nor2  gate558(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate559(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate560(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1513(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1514(.a(gate175inter0), .b(s_138), .O(gate175inter1));
  and2  gate1515(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1516(.a(s_138), .O(gate175inter3));
  inv1  gate1517(.a(s_139), .O(gate175inter4));
  nand2 gate1518(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1519(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1520(.a(G492), .O(gate175inter7));
  inv1  gate1521(.a(G555), .O(gate175inter8));
  nand2 gate1522(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1523(.a(s_139), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1524(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1525(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1526(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate617(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate618(.a(gate190inter0), .b(s_10), .O(gate190inter1));
  and2  gate619(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate620(.a(s_10), .O(gate190inter3));
  inv1  gate621(.a(s_11), .O(gate190inter4));
  nand2 gate622(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate623(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate624(.a(G580), .O(gate190inter7));
  inv1  gate625(.a(G581), .O(gate190inter8));
  nand2 gate626(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate627(.a(s_11), .b(gate190inter3), .O(gate190inter10));
  nor2  gate628(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate629(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate630(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate701(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate702(.a(gate192inter0), .b(s_22), .O(gate192inter1));
  and2  gate703(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate704(.a(s_22), .O(gate192inter3));
  inv1  gate705(.a(s_23), .O(gate192inter4));
  nand2 gate706(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate707(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate708(.a(G584), .O(gate192inter7));
  inv1  gate709(.a(G585), .O(gate192inter8));
  nand2 gate710(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate711(.a(s_23), .b(gate192inter3), .O(gate192inter10));
  nor2  gate712(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate713(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate714(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1037(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1038(.a(gate193inter0), .b(s_70), .O(gate193inter1));
  and2  gate1039(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1040(.a(s_70), .O(gate193inter3));
  inv1  gate1041(.a(s_71), .O(gate193inter4));
  nand2 gate1042(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1043(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1044(.a(G586), .O(gate193inter7));
  inv1  gate1045(.a(G587), .O(gate193inter8));
  nand2 gate1046(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1047(.a(s_71), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1048(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1049(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1050(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1597(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1598(.a(gate197inter0), .b(s_150), .O(gate197inter1));
  and2  gate1599(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1600(.a(s_150), .O(gate197inter3));
  inv1  gate1601(.a(s_151), .O(gate197inter4));
  nand2 gate1602(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1603(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1604(.a(G594), .O(gate197inter7));
  inv1  gate1605(.a(G595), .O(gate197inter8));
  nand2 gate1606(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1607(.a(s_151), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1608(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1609(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1610(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate561(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate562(.a(gate204inter0), .b(s_2), .O(gate204inter1));
  and2  gate563(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate564(.a(s_2), .O(gate204inter3));
  inv1  gate565(.a(s_3), .O(gate204inter4));
  nand2 gate566(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate567(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate568(.a(G607), .O(gate204inter7));
  inv1  gate569(.a(G617), .O(gate204inter8));
  nand2 gate570(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate571(.a(s_3), .b(gate204inter3), .O(gate204inter10));
  nor2  gate572(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate573(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate574(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate995(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate996(.a(gate205inter0), .b(s_64), .O(gate205inter1));
  and2  gate997(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate998(.a(s_64), .O(gate205inter3));
  inv1  gate999(.a(s_65), .O(gate205inter4));
  nand2 gate1000(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1001(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1002(.a(G622), .O(gate205inter7));
  inv1  gate1003(.a(G627), .O(gate205inter8));
  nand2 gate1004(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1005(.a(s_65), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1006(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1007(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1008(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1247(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1248(.a(gate211inter0), .b(s_100), .O(gate211inter1));
  and2  gate1249(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1250(.a(s_100), .O(gate211inter3));
  inv1  gate1251(.a(s_101), .O(gate211inter4));
  nand2 gate1252(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1253(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1254(.a(G612), .O(gate211inter7));
  inv1  gate1255(.a(G669), .O(gate211inter8));
  nand2 gate1256(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1257(.a(s_101), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1258(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1259(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1260(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1135(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1136(.a(gate219inter0), .b(s_84), .O(gate219inter1));
  and2  gate1137(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1138(.a(s_84), .O(gate219inter3));
  inv1  gate1139(.a(s_85), .O(gate219inter4));
  nand2 gate1140(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1141(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1142(.a(G632), .O(gate219inter7));
  inv1  gate1143(.a(G681), .O(gate219inter8));
  nand2 gate1144(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1145(.a(s_85), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1146(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1147(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1148(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1485(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1486(.a(gate224inter0), .b(s_134), .O(gate224inter1));
  and2  gate1487(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1488(.a(s_134), .O(gate224inter3));
  inv1  gate1489(.a(s_135), .O(gate224inter4));
  nand2 gate1490(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1491(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1492(.a(G637), .O(gate224inter7));
  inv1  gate1493(.a(G687), .O(gate224inter8));
  nand2 gate1494(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1495(.a(s_135), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1496(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1497(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1498(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate589(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate590(.a(gate226inter0), .b(s_6), .O(gate226inter1));
  and2  gate591(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate592(.a(s_6), .O(gate226inter3));
  inv1  gate593(.a(s_7), .O(gate226inter4));
  nand2 gate594(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate595(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate596(.a(G692), .O(gate226inter7));
  inv1  gate597(.a(G693), .O(gate226inter8));
  nand2 gate598(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate599(.a(s_7), .b(gate226inter3), .O(gate226inter10));
  nor2  gate600(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate601(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate602(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1303(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1304(.a(gate231inter0), .b(s_108), .O(gate231inter1));
  and2  gate1305(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1306(.a(s_108), .O(gate231inter3));
  inv1  gate1307(.a(s_109), .O(gate231inter4));
  nand2 gate1308(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1309(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1310(.a(G702), .O(gate231inter7));
  inv1  gate1311(.a(G703), .O(gate231inter8));
  nand2 gate1312(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1313(.a(s_109), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1314(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1315(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1316(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1121(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1122(.a(gate234inter0), .b(s_82), .O(gate234inter1));
  and2  gate1123(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1124(.a(s_82), .O(gate234inter3));
  inv1  gate1125(.a(s_83), .O(gate234inter4));
  nand2 gate1126(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1127(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1128(.a(G245), .O(gate234inter7));
  inv1  gate1129(.a(G721), .O(gate234inter8));
  nand2 gate1130(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1131(.a(s_83), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1132(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1133(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1134(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1233(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1234(.a(gate235inter0), .b(s_98), .O(gate235inter1));
  and2  gate1235(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1236(.a(s_98), .O(gate235inter3));
  inv1  gate1237(.a(s_99), .O(gate235inter4));
  nand2 gate1238(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1239(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1240(.a(G248), .O(gate235inter7));
  inv1  gate1241(.a(G724), .O(gate235inter8));
  nand2 gate1242(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1243(.a(s_99), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1244(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1245(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1246(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate771(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate772(.a(gate237inter0), .b(s_32), .O(gate237inter1));
  and2  gate773(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate774(.a(s_32), .O(gate237inter3));
  inv1  gate775(.a(s_33), .O(gate237inter4));
  nand2 gate776(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate777(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate778(.a(G254), .O(gate237inter7));
  inv1  gate779(.a(G706), .O(gate237inter8));
  nand2 gate780(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate781(.a(s_33), .b(gate237inter3), .O(gate237inter10));
  nor2  gate782(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate783(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate784(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate925(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate926(.a(gate239inter0), .b(s_54), .O(gate239inter1));
  and2  gate927(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate928(.a(s_54), .O(gate239inter3));
  inv1  gate929(.a(s_55), .O(gate239inter4));
  nand2 gate930(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate931(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate932(.a(G260), .O(gate239inter7));
  inv1  gate933(.a(G712), .O(gate239inter8));
  nand2 gate934(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate935(.a(s_55), .b(gate239inter3), .O(gate239inter10));
  nor2  gate936(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate937(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate938(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate827(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate828(.a(gate244inter0), .b(s_40), .O(gate244inter1));
  and2  gate829(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate830(.a(s_40), .O(gate244inter3));
  inv1  gate831(.a(s_41), .O(gate244inter4));
  nand2 gate832(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate833(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate834(.a(G721), .O(gate244inter7));
  inv1  gate835(.a(G733), .O(gate244inter8));
  nand2 gate836(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate837(.a(s_41), .b(gate244inter3), .O(gate244inter10));
  nor2  gate838(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate839(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate840(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1527(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1528(.a(gate249inter0), .b(s_140), .O(gate249inter1));
  and2  gate1529(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1530(.a(s_140), .O(gate249inter3));
  inv1  gate1531(.a(s_141), .O(gate249inter4));
  nand2 gate1532(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1533(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1534(.a(G254), .O(gate249inter7));
  inv1  gate1535(.a(G742), .O(gate249inter8));
  nand2 gate1536(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1537(.a(s_141), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1538(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1539(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1540(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate603(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate604(.a(gate257inter0), .b(s_8), .O(gate257inter1));
  and2  gate605(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate606(.a(s_8), .O(gate257inter3));
  inv1  gate607(.a(s_9), .O(gate257inter4));
  nand2 gate608(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate609(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate610(.a(G754), .O(gate257inter7));
  inv1  gate611(.a(G755), .O(gate257inter8));
  nand2 gate612(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate613(.a(s_9), .b(gate257inter3), .O(gate257inter10));
  nor2  gate614(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate615(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate616(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate869(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate870(.a(gate259inter0), .b(s_46), .O(gate259inter1));
  and2  gate871(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate872(.a(s_46), .O(gate259inter3));
  inv1  gate873(.a(s_47), .O(gate259inter4));
  nand2 gate874(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate875(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate876(.a(G758), .O(gate259inter7));
  inv1  gate877(.a(G759), .O(gate259inter8));
  nand2 gate878(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate879(.a(s_47), .b(gate259inter3), .O(gate259inter10));
  nor2  gate880(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate881(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate882(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1471(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1472(.a(gate262inter0), .b(s_132), .O(gate262inter1));
  and2  gate1473(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1474(.a(s_132), .O(gate262inter3));
  inv1  gate1475(.a(s_133), .O(gate262inter4));
  nand2 gate1476(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1477(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1478(.a(G764), .O(gate262inter7));
  inv1  gate1479(.a(G765), .O(gate262inter8));
  nand2 gate1480(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1481(.a(s_133), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1482(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1483(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1484(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate785(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate786(.a(gate263inter0), .b(s_34), .O(gate263inter1));
  and2  gate787(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate788(.a(s_34), .O(gate263inter3));
  inv1  gate789(.a(s_35), .O(gate263inter4));
  nand2 gate790(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate791(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate792(.a(G766), .O(gate263inter7));
  inv1  gate793(.a(G767), .O(gate263inter8));
  nand2 gate794(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate795(.a(s_35), .b(gate263inter3), .O(gate263inter10));
  nor2  gate796(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate797(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate798(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate841(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate842(.a(gate266inter0), .b(s_42), .O(gate266inter1));
  and2  gate843(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate844(.a(s_42), .O(gate266inter3));
  inv1  gate845(.a(s_43), .O(gate266inter4));
  nand2 gate846(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate847(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate848(.a(G645), .O(gate266inter7));
  inv1  gate849(.a(G773), .O(gate266inter8));
  nand2 gate850(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate851(.a(s_43), .b(gate266inter3), .O(gate266inter10));
  nor2  gate852(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate853(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate854(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1401(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1402(.a(gate270inter0), .b(s_122), .O(gate270inter1));
  and2  gate1403(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1404(.a(s_122), .O(gate270inter3));
  inv1  gate1405(.a(s_123), .O(gate270inter4));
  nand2 gate1406(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1407(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1408(.a(G657), .O(gate270inter7));
  inv1  gate1409(.a(G785), .O(gate270inter8));
  nand2 gate1410(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1411(.a(s_123), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1412(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1413(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1414(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate897(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate898(.a(gate274inter0), .b(s_50), .O(gate274inter1));
  and2  gate899(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate900(.a(s_50), .O(gate274inter3));
  inv1  gate901(.a(s_51), .O(gate274inter4));
  nand2 gate902(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate903(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate904(.a(G770), .O(gate274inter7));
  inv1  gate905(.a(G794), .O(gate274inter8));
  nand2 gate906(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate907(.a(s_51), .b(gate274inter3), .O(gate274inter10));
  nor2  gate908(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate909(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate910(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1359(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1360(.a(gate285inter0), .b(s_116), .O(gate285inter1));
  and2  gate1361(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1362(.a(s_116), .O(gate285inter3));
  inv1  gate1363(.a(s_117), .O(gate285inter4));
  nand2 gate1364(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1365(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1366(.a(G660), .O(gate285inter7));
  inv1  gate1367(.a(G812), .O(gate285inter8));
  nand2 gate1368(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1369(.a(s_117), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1370(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1371(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1372(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate659(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate660(.a(gate291inter0), .b(s_16), .O(gate291inter1));
  and2  gate661(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate662(.a(s_16), .O(gate291inter3));
  inv1  gate663(.a(s_17), .O(gate291inter4));
  nand2 gate664(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate665(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate666(.a(G822), .O(gate291inter7));
  inv1  gate667(.a(G823), .O(gate291inter8));
  nand2 gate668(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate669(.a(s_17), .b(gate291inter3), .O(gate291inter10));
  nor2  gate670(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate671(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate672(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1009(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1010(.a(gate394inter0), .b(s_66), .O(gate394inter1));
  and2  gate1011(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1012(.a(s_66), .O(gate394inter3));
  inv1  gate1013(.a(s_67), .O(gate394inter4));
  nand2 gate1014(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1015(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1016(.a(G8), .O(gate394inter7));
  inv1  gate1017(.a(G1057), .O(gate394inter8));
  nand2 gate1018(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1019(.a(s_67), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1020(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1021(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1022(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1373(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1374(.a(gate408inter0), .b(s_118), .O(gate408inter1));
  and2  gate1375(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1376(.a(s_118), .O(gate408inter3));
  inv1  gate1377(.a(s_119), .O(gate408inter4));
  nand2 gate1378(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1379(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1380(.a(G22), .O(gate408inter7));
  inv1  gate1381(.a(G1099), .O(gate408inter8));
  nand2 gate1382(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1383(.a(s_119), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1384(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1385(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1386(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1051(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1052(.a(gate410inter0), .b(s_72), .O(gate410inter1));
  and2  gate1053(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1054(.a(s_72), .O(gate410inter3));
  inv1  gate1055(.a(s_73), .O(gate410inter4));
  nand2 gate1056(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1057(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1058(.a(G24), .O(gate410inter7));
  inv1  gate1059(.a(G1105), .O(gate410inter8));
  nand2 gate1060(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1061(.a(s_73), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1062(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1063(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1064(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1149(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1150(.a(gate411inter0), .b(s_86), .O(gate411inter1));
  and2  gate1151(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1152(.a(s_86), .O(gate411inter3));
  inv1  gate1153(.a(s_87), .O(gate411inter4));
  nand2 gate1154(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1155(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1156(.a(G25), .O(gate411inter7));
  inv1  gate1157(.a(G1108), .O(gate411inter8));
  nand2 gate1158(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1159(.a(s_87), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1160(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1161(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1162(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate883(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate884(.a(gate413inter0), .b(s_48), .O(gate413inter1));
  and2  gate885(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate886(.a(s_48), .O(gate413inter3));
  inv1  gate887(.a(s_49), .O(gate413inter4));
  nand2 gate888(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate889(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate890(.a(G27), .O(gate413inter7));
  inv1  gate891(.a(G1114), .O(gate413inter8));
  nand2 gate892(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate893(.a(s_49), .b(gate413inter3), .O(gate413inter10));
  nor2  gate894(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate895(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate896(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1289(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1290(.a(gate419inter0), .b(s_106), .O(gate419inter1));
  and2  gate1291(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1292(.a(s_106), .O(gate419inter3));
  inv1  gate1293(.a(s_107), .O(gate419inter4));
  nand2 gate1294(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1295(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1296(.a(G1), .O(gate419inter7));
  inv1  gate1297(.a(G1132), .O(gate419inter8));
  nand2 gate1298(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1299(.a(s_107), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1300(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1301(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1302(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1261(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1262(.a(gate428inter0), .b(s_102), .O(gate428inter1));
  and2  gate1263(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1264(.a(s_102), .O(gate428inter3));
  inv1  gate1265(.a(s_103), .O(gate428inter4));
  nand2 gate1266(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1267(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1268(.a(G1048), .O(gate428inter7));
  inv1  gate1269(.a(G1144), .O(gate428inter8));
  nand2 gate1270(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1271(.a(s_103), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1272(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1273(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1274(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1219(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1220(.a(gate437inter0), .b(s_96), .O(gate437inter1));
  and2  gate1221(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1222(.a(s_96), .O(gate437inter3));
  inv1  gate1223(.a(s_97), .O(gate437inter4));
  nand2 gate1224(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1225(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1226(.a(G10), .O(gate437inter7));
  inv1  gate1227(.a(G1159), .O(gate437inter8));
  nand2 gate1228(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1229(.a(s_97), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1230(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1231(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1232(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate757(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate758(.a(gate441inter0), .b(s_30), .O(gate441inter1));
  and2  gate759(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate760(.a(s_30), .O(gate441inter3));
  inv1  gate761(.a(s_31), .O(gate441inter4));
  nand2 gate762(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate763(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate764(.a(G12), .O(gate441inter7));
  inv1  gate765(.a(G1165), .O(gate441inter8));
  nand2 gate766(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate767(.a(s_31), .b(gate441inter3), .O(gate441inter10));
  nor2  gate768(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate769(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate770(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate855(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate856(.a(gate456inter0), .b(s_44), .O(gate456inter1));
  and2  gate857(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate858(.a(s_44), .O(gate456inter3));
  inv1  gate859(.a(s_45), .O(gate456inter4));
  nand2 gate860(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate861(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate862(.a(G1090), .O(gate456inter7));
  inv1  gate863(.a(G1186), .O(gate456inter8));
  nand2 gate864(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate865(.a(s_45), .b(gate456inter3), .O(gate456inter10));
  nor2  gate866(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate867(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate868(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate939(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate940(.a(gate509inter0), .b(s_56), .O(gate509inter1));
  and2  gate941(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate942(.a(s_56), .O(gate509inter3));
  inv1  gate943(.a(s_57), .O(gate509inter4));
  nand2 gate944(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate945(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate946(.a(G1280), .O(gate509inter7));
  inv1  gate947(.a(G1281), .O(gate509inter8));
  nand2 gate948(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate949(.a(s_57), .b(gate509inter3), .O(gate509inter10));
  nor2  gate950(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate951(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate952(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1429(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1430(.a(gate512inter0), .b(s_126), .O(gate512inter1));
  and2  gate1431(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1432(.a(s_126), .O(gate512inter3));
  inv1  gate1433(.a(s_127), .O(gate512inter4));
  nand2 gate1434(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1435(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1436(.a(G1286), .O(gate512inter7));
  inv1  gate1437(.a(G1287), .O(gate512inter8));
  nand2 gate1438(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1439(.a(s_127), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1440(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1441(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1442(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1107(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1108(.a(gate513inter0), .b(s_80), .O(gate513inter1));
  and2  gate1109(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1110(.a(s_80), .O(gate513inter3));
  inv1  gate1111(.a(s_81), .O(gate513inter4));
  nand2 gate1112(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1113(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1114(.a(G1288), .O(gate513inter7));
  inv1  gate1115(.a(G1289), .O(gate513inter8));
  nand2 gate1116(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1117(.a(s_81), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1118(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1119(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1120(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule