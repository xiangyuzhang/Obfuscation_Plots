module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1443(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1444(.a(gate13inter0), .b(s_128), .O(gate13inter1));
  and2  gate1445(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1446(.a(s_128), .O(gate13inter3));
  inv1  gate1447(.a(s_129), .O(gate13inter4));
  nand2 gate1448(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1449(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1450(.a(G9), .O(gate13inter7));
  inv1  gate1451(.a(G10), .O(gate13inter8));
  nand2 gate1452(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1453(.a(s_129), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1454(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1455(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1456(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1499(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1500(.a(gate17inter0), .b(s_136), .O(gate17inter1));
  and2  gate1501(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1502(.a(s_136), .O(gate17inter3));
  inv1  gate1503(.a(s_137), .O(gate17inter4));
  nand2 gate1504(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1505(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1506(.a(G17), .O(gate17inter7));
  inv1  gate1507(.a(G18), .O(gate17inter8));
  nand2 gate1508(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1509(.a(s_137), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1510(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1511(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1512(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1205(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1206(.a(gate21inter0), .b(s_94), .O(gate21inter1));
  and2  gate1207(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1208(.a(s_94), .O(gate21inter3));
  inv1  gate1209(.a(s_95), .O(gate21inter4));
  nand2 gate1210(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1211(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1212(.a(G25), .O(gate21inter7));
  inv1  gate1213(.a(G26), .O(gate21inter8));
  nand2 gate1214(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1215(.a(s_95), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1216(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1217(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1218(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1121(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1122(.a(gate23inter0), .b(s_82), .O(gate23inter1));
  and2  gate1123(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1124(.a(s_82), .O(gate23inter3));
  inv1  gate1125(.a(s_83), .O(gate23inter4));
  nand2 gate1126(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1127(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1128(.a(G29), .O(gate23inter7));
  inv1  gate1129(.a(G30), .O(gate23inter8));
  nand2 gate1130(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1131(.a(s_83), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1132(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1133(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1134(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate883(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate884(.a(gate25inter0), .b(s_48), .O(gate25inter1));
  and2  gate885(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate886(.a(s_48), .O(gate25inter3));
  inv1  gate887(.a(s_49), .O(gate25inter4));
  nand2 gate888(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate889(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate890(.a(G1), .O(gate25inter7));
  inv1  gate891(.a(G5), .O(gate25inter8));
  nand2 gate892(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate893(.a(s_49), .b(gate25inter3), .O(gate25inter10));
  nor2  gate894(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate895(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate896(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate981(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate982(.a(gate32inter0), .b(s_62), .O(gate32inter1));
  and2  gate983(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate984(.a(s_62), .O(gate32inter3));
  inv1  gate985(.a(s_63), .O(gate32inter4));
  nand2 gate986(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate987(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate988(.a(G12), .O(gate32inter7));
  inv1  gate989(.a(G16), .O(gate32inter8));
  nand2 gate990(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate991(.a(s_63), .b(gate32inter3), .O(gate32inter10));
  nor2  gate992(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate993(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate994(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1583(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1584(.a(gate41inter0), .b(s_148), .O(gate41inter1));
  and2  gate1585(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1586(.a(s_148), .O(gate41inter3));
  inv1  gate1587(.a(s_149), .O(gate41inter4));
  nand2 gate1588(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1589(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1590(.a(G1), .O(gate41inter7));
  inv1  gate1591(.a(G266), .O(gate41inter8));
  nand2 gate1592(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1593(.a(s_149), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1594(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1595(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1596(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1177(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1178(.a(gate48inter0), .b(s_90), .O(gate48inter1));
  and2  gate1179(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1180(.a(s_90), .O(gate48inter3));
  inv1  gate1181(.a(s_91), .O(gate48inter4));
  nand2 gate1182(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1183(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1184(.a(G8), .O(gate48inter7));
  inv1  gate1185(.a(G275), .O(gate48inter8));
  nand2 gate1186(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1187(.a(s_91), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1188(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1189(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1190(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1541(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1542(.a(gate51inter0), .b(s_142), .O(gate51inter1));
  and2  gate1543(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1544(.a(s_142), .O(gate51inter3));
  inv1  gate1545(.a(s_143), .O(gate51inter4));
  nand2 gate1546(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1547(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1548(.a(G11), .O(gate51inter7));
  inv1  gate1549(.a(G281), .O(gate51inter8));
  nand2 gate1550(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1551(.a(s_143), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1552(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1553(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1554(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1331(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1332(.a(gate54inter0), .b(s_112), .O(gate54inter1));
  and2  gate1333(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1334(.a(s_112), .O(gate54inter3));
  inv1  gate1335(.a(s_113), .O(gate54inter4));
  nand2 gate1336(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1337(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1338(.a(G14), .O(gate54inter7));
  inv1  gate1339(.a(G284), .O(gate54inter8));
  nand2 gate1340(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1341(.a(s_113), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1342(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1343(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1344(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate813(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate814(.a(gate58inter0), .b(s_38), .O(gate58inter1));
  and2  gate815(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate816(.a(s_38), .O(gate58inter3));
  inv1  gate817(.a(s_39), .O(gate58inter4));
  nand2 gate818(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate819(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate820(.a(G18), .O(gate58inter7));
  inv1  gate821(.a(G290), .O(gate58inter8));
  nand2 gate822(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate823(.a(s_39), .b(gate58inter3), .O(gate58inter10));
  nor2  gate824(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate825(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate826(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate687(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate688(.a(gate59inter0), .b(s_20), .O(gate59inter1));
  and2  gate689(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate690(.a(s_20), .O(gate59inter3));
  inv1  gate691(.a(s_21), .O(gate59inter4));
  nand2 gate692(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate693(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate694(.a(G19), .O(gate59inter7));
  inv1  gate695(.a(G293), .O(gate59inter8));
  nand2 gate696(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate697(.a(s_21), .b(gate59inter3), .O(gate59inter10));
  nor2  gate698(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate699(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate700(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1415(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1416(.a(gate61inter0), .b(s_124), .O(gate61inter1));
  and2  gate1417(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1418(.a(s_124), .O(gate61inter3));
  inv1  gate1419(.a(s_125), .O(gate61inter4));
  nand2 gate1420(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1421(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1422(.a(G21), .O(gate61inter7));
  inv1  gate1423(.a(G296), .O(gate61inter8));
  nand2 gate1424(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1425(.a(s_125), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1426(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1427(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1428(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate841(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate842(.a(gate68inter0), .b(s_42), .O(gate68inter1));
  and2  gate843(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate844(.a(s_42), .O(gate68inter3));
  inv1  gate845(.a(s_43), .O(gate68inter4));
  nand2 gate846(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate847(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate848(.a(G28), .O(gate68inter7));
  inv1  gate849(.a(G305), .O(gate68inter8));
  nand2 gate850(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate851(.a(s_43), .b(gate68inter3), .O(gate68inter10));
  nor2  gate852(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate853(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate854(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1303(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1304(.a(gate72inter0), .b(s_108), .O(gate72inter1));
  and2  gate1305(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1306(.a(s_108), .O(gate72inter3));
  inv1  gate1307(.a(s_109), .O(gate72inter4));
  nand2 gate1308(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1309(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1310(.a(G32), .O(gate72inter7));
  inv1  gate1311(.a(G311), .O(gate72inter8));
  nand2 gate1312(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1313(.a(s_109), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1314(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1315(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1316(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1023(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1024(.a(gate84inter0), .b(s_68), .O(gate84inter1));
  and2  gate1025(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1026(.a(s_68), .O(gate84inter3));
  inv1  gate1027(.a(s_69), .O(gate84inter4));
  nand2 gate1028(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1029(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1030(.a(G15), .O(gate84inter7));
  inv1  gate1031(.a(G329), .O(gate84inter8));
  nand2 gate1032(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1033(.a(s_69), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1034(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1035(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1036(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate561(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate562(.a(gate88inter0), .b(s_2), .O(gate88inter1));
  and2  gate563(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate564(.a(s_2), .O(gate88inter3));
  inv1  gate565(.a(s_3), .O(gate88inter4));
  nand2 gate566(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate567(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate568(.a(G16), .O(gate88inter7));
  inv1  gate569(.a(G335), .O(gate88inter8));
  nand2 gate570(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate571(.a(s_3), .b(gate88inter3), .O(gate88inter10));
  nor2  gate572(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate573(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate574(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1247(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1248(.a(gate92inter0), .b(s_100), .O(gate92inter1));
  and2  gate1249(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1250(.a(s_100), .O(gate92inter3));
  inv1  gate1251(.a(s_101), .O(gate92inter4));
  nand2 gate1252(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1253(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1254(.a(G29), .O(gate92inter7));
  inv1  gate1255(.a(G341), .O(gate92inter8));
  nand2 gate1256(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1257(.a(s_101), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1258(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1259(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1260(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate575(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate576(.a(gate93inter0), .b(s_4), .O(gate93inter1));
  and2  gate577(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate578(.a(s_4), .O(gate93inter3));
  inv1  gate579(.a(s_5), .O(gate93inter4));
  nand2 gate580(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate581(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate582(.a(G18), .O(gate93inter7));
  inv1  gate583(.a(G344), .O(gate93inter8));
  nand2 gate584(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate585(.a(s_5), .b(gate93inter3), .O(gate93inter10));
  nor2  gate586(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate587(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate588(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1065(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1066(.a(gate97inter0), .b(s_74), .O(gate97inter1));
  and2  gate1067(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1068(.a(s_74), .O(gate97inter3));
  inv1  gate1069(.a(s_75), .O(gate97inter4));
  nand2 gate1070(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1071(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1072(.a(G19), .O(gate97inter7));
  inv1  gate1073(.a(G350), .O(gate97inter8));
  nand2 gate1074(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1075(.a(s_75), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1076(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1077(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1078(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate869(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate870(.a(gate101inter0), .b(s_46), .O(gate101inter1));
  and2  gate871(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate872(.a(s_46), .O(gate101inter3));
  inv1  gate873(.a(s_47), .O(gate101inter4));
  nand2 gate874(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate875(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate876(.a(G20), .O(gate101inter7));
  inv1  gate877(.a(G356), .O(gate101inter8));
  nand2 gate878(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate879(.a(s_47), .b(gate101inter3), .O(gate101inter10));
  nor2  gate880(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate881(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate882(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1527(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1528(.a(gate104inter0), .b(s_140), .O(gate104inter1));
  and2  gate1529(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1530(.a(s_140), .O(gate104inter3));
  inv1  gate1531(.a(s_141), .O(gate104inter4));
  nand2 gate1532(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1533(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1534(.a(G32), .O(gate104inter7));
  inv1  gate1535(.a(G359), .O(gate104inter8));
  nand2 gate1536(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1537(.a(s_141), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1538(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1539(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1540(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1051(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1052(.a(gate105inter0), .b(s_72), .O(gate105inter1));
  and2  gate1053(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1054(.a(s_72), .O(gate105inter3));
  inv1  gate1055(.a(s_73), .O(gate105inter4));
  nand2 gate1056(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1057(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1058(.a(G362), .O(gate105inter7));
  inv1  gate1059(.a(G363), .O(gate105inter8));
  nand2 gate1060(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1061(.a(s_73), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1062(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1063(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1064(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate939(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate940(.a(gate118inter0), .b(s_56), .O(gate118inter1));
  and2  gate941(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate942(.a(s_56), .O(gate118inter3));
  inv1  gate943(.a(s_57), .O(gate118inter4));
  nand2 gate944(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate945(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate946(.a(G388), .O(gate118inter7));
  inv1  gate947(.a(G389), .O(gate118inter8));
  nand2 gate948(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate949(.a(s_57), .b(gate118inter3), .O(gate118inter10));
  nor2  gate950(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate951(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate952(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1093(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1094(.a(gate120inter0), .b(s_78), .O(gate120inter1));
  and2  gate1095(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1096(.a(s_78), .O(gate120inter3));
  inv1  gate1097(.a(s_79), .O(gate120inter4));
  nand2 gate1098(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1099(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1100(.a(G392), .O(gate120inter7));
  inv1  gate1101(.a(G393), .O(gate120inter8));
  nand2 gate1102(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1103(.a(s_79), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1104(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1105(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1106(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate967(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate968(.a(gate123inter0), .b(s_60), .O(gate123inter1));
  and2  gate969(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate970(.a(s_60), .O(gate123inter3));
  inv1  gate971(.a(s_61), .O(gate123inter4));
  nand2 gate972(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate973(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate974(.a(G398), .O(gate123inter7));
  inv1  gate975(.a(G399), .O(gate123inter8));
  nand2 gate976(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate977(.a(s_61), .b(gate123inter3), .O(gate123inter10));
  nor2  gate978(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate979(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate980(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate645(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate646(.a(gate136inter0), .b(s_14), .O(gate136inter1));
  and2  gate647(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate648(.a(s_14), .O(gate136inter3));
  inv1  gate649(.a(s_15), .O(gate136inter4));
  nand2 gate650(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate651(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate652(.a(G424), .O(gate136inter7));
  inv1  gate653(.a(G425), .O(gate136inter8));
  nand2 gate654(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate655(.a(s_15), .b(gate136inter3), .O(gate136inter10));
  nor2  gate656(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate657(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate658(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate729(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate730(.a(gate157inter0), .b(s_26), .O(gate157inter1));
  and2  gate731(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate732(.a(s_26), .O(gate157inter3));
  inv1  gate733(.a(s_27), .O(gate157inter4));
  nand2 gate734(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate735(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate736(.a(G438), .O(gate157inter7));
  inv1  gate737(.a(G528), .O(gate157inter8));
  nand2 gate738(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate739(.a(s_27), .b(gate157inter3), .O(gate157inter10));
  nor2  gate740(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate741(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate742(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate855(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate856(.a(gate159inter0), .b(s_44), .O(gate159inter1));
  and2  gate857(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate858(.a(s_44), .O(gate159inter3));
  inv1  gate859(.a(s_45), .O(gate159inter4));
  nand2 gate860(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate861(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate862(.a(G444), .O(gate159inter7));
  inv1  gate863(.a(G531), .O(gate159inter8));
  nand2 gate864(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate865(.a(s_45), .b(gate159inter3), .O(gate159inter10));
  nor2  gate866(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate867(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate868(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate953(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate954(.a(gate162inter0), .b(s_58), .O(gate162inter1));
  and2  gate955(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate956(.a(s_58), .O(gate162inter3));
  inv1  gate957(.a(s_59), .O(gate162inter4));
  nand2 gate958(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate959(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate960(.a(G453), .O(gate162inter7));
  inv1  gate961(.a(G534), .O(gate162inter8));
  nand2 gate962(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate963(.a(s_59), .b(gate162inter3), .O(gate162inter10));
  nor2  gate964(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate965(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate966(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1261(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1262(.a(gate169inter0), .b(s_102), .O(gate169inter1));
  and2  gate1263(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1264(.a(s_102), .O(gate169inter3));
  inv1  gate1265(.a(s_103), .O(gate169inter4));
  nand2 gate1266(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1267(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1268(.a(G474), .O(gate169inter7));
  inv1  gate1269(.a(G546), .O(gate169inter8));
  nand2 gate1270(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1271(.a(s_103), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1272(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1273(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1274(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1163(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1164(.a(gate170inter0), .b(s_88), .O(gate170inter1));
  and2  gate1165(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1166(.a(s_88), .O(gate170inter3));
  inv1  gate1167(.a(s_89), .O(gate170inter4));
  nand2 gate1168(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1169(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1170(.a(G477), .O(gate170inter7));
  inv1  gate1171(.a(G546), .O(gate170inter8));
  nand2 gate1172(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1173(.a(s_89), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1174(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1175(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1176(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1009(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1010(.a(gate186inter0), .b(s_66), .O(gate186inter1));
  and2  gate1011(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1012(.a(s_66), .O(gate186inter3));
  inv1  gate1013(.a(s_67), .O(gate186inter4));
  nand2 gate1014(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1015(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1016(.a(G572), .O(gate186inter7));
  inv1  gate1017(.a(G573), .O(gate186inter8));
  nand2 gate1018(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1019(.a(s_67), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1020(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1021(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1022(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1555(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1556(.a(gate187inter0), .b(s_144), .O(gate187inter1));
  and2  gate1557(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1558(.a(s_144), .O(gate187inter3));
  inv1  gate1559(.a(s_145), .O(gate187inter4));
  nand2 gate1560(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1561(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1562(.a(G574), .O(gate187inter7));
  inv1  gate1563(.a(G575), .O(gate187inter8));
  nand2 gate1564(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1565(.a(s_145), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1566(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1567(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1568(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate589(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate590(.a(gate192inter0), .b(s_6), .O(gate192inter1));
  and2  gate591(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate592(.a(s_6), .O(gate192inter3));
  inv1  gate593(.a(s_7), .O(gate192inter4));
  nand2 gate594(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate595(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate596(.a(G584), .O(gate192inter7));
  inv1  gate597(.a(G585), .O(gate192inter8));
  nand2 gate598(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate599(.a(s_7), .b(gate192inter3), .O(gate192inter10));
  nor2  gate600(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate601(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate602(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1471(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1472(.a(gate194inter0), .b(s_132), .O(gate194inter1));
  and2  gate1473(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1474(.a(s_132), .O(gate194inter3));
  inv1  gate1475(.a(s_133), .O(gate194inter4));
  nand2 gate1476(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1477(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1478(.a(G588), .O(gate194inter7));
  inv1  gate1479(.a(G589), .O(gate194inter8));
  nand2 gate1480(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1481(.a(s_133), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1482(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1483(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1484(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate659(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate660(.a(gate199inter0), .b(s_16), .O(gate199inter1));
  and2  gate661(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate662(.a(s_16), .O(gate199inter3));
  inv1  gate663(.a(s_17), .O(gate199inter4));
  nand2 gate664(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate665(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate666(.a(G598), .O(gate199inter7));
  inv1  gate667(.a(G599), .O(gate199inter8));
  nand2 gate668(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate669(.a(s_17), .b(gate199inter3), .O(gate199inter10));
  nor2  gate670(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate671(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate672(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate617(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate618(.a(gate202inter0), .b(s_10), .O(gate202inter1));
  and2  gate619(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate620(.a(s_10), .O(gate202inter3));
  inv1  gate621(.a(s_11), .O(gate202inter4));
  nand2 gate622(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate623(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate624(.a(G612), .O(gate202inter7));
  inv1  gate625(.a(G617), .O(gate202inter8));
  nand2 gate626(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate627(.a(s_11), .b(gate202inter3), .O(gate202inter10));
  nor2  gate628(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate629(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate630(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate771(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate772(.a(gate203inter0), .b(s_32), .O(gate203inter1));
  and2  gate773(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate774(.a(s_32), .O(gate203inter3));
  inv1  gate775(.a(s_33), .O(gate203inter4));
  nand2 gate776(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate777(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate778(.a(G602), .O(gate203inter7));
  inv1  gate779(.a(G612), .O(gate203inter8));
  nand2 gate780(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate781(.a(s_33), .b(gate203inter3), .O(gate203inter10));
  nor2  gate782(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate783(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate784(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate925(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate926(.a(gate204inter0), .b(s_54), .O(gate204inter1));
  and2  gate927(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate928(.a(s_54), .O(gate204inter3));
  inv1  gate929(.a(s_55), .O(gate204inter4));
  nand2 gate930(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate931(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate932(.a(G607), .O(gate204inter7));
  inv1  gate933(.a(G617), .O(gate204inter8));
  nand2 gate934(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate935(.a(s_55), .b(gate204inter3), .O(gate204inter10));
  nor2  gate936(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate937(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate938(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate897(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate898(.a(gate206inter0), .b(s_50), .O(gate206inter1));
  and2  gate899(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate900(.a(s_50), .O(gate206inter3));
  inv1  gate901(.a(s_51), .O(gate206inter4));
  nand2 gate902(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate903(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate904(.a(G632), .O(gate206inter7));
  inv1  gate905(.a(G637), .O(gate206inter8));
  nand2 gate906(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate907(.a(s_51), .b(gate206inter3), .O(gate206inter10));
  nor2  gate908(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate909(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate910(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1569(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1570(.a(gate207inter0), .b(s_146), .O(gate207inter1));
  and2  gate1571(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1572(.a(s_146), .O(gate207inter3));
  inv1  gate1573(.a(s_147), .O(gate207inter4));
  nand2 gate1574(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1575(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1576(.a(G622), .O(gate207inter7));
  inv1  gate1577(.a(G632), .O(gate207inter8));
  nand2 gate1578(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1579(.a(s_147), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1580(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1581(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1582(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1387(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1388(.a(gate213inter0), .b(s_120), .O(gate213inter1));
  and2  gate1389(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1390(.a(s_120), .O(gate213inter3));
  inv1  gate1391(.a(s_121), .O(gate213inter4));
  nand2 gate1392(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1393(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1394(.a(G602), .O(gate213inter7));
  inv1  gate1395(.a(G672), .O(gate213inter8));
  nand2 gate1396(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1397(.a(s_121), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1398(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1399(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1400(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate827(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate828(.a(gate219inter0), .b(s_40), .O(gate219inter1));
  and2  gate829(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate830(.a(s_40), .O(gate219inter3));
  inv1  gate831(.a(s_41), .O(gate219inter4));
  nand2 gate832(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate833(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate834(.a(G632), .O(gate219inter7));
  inv1  gate835(.a(G681), .O(gate219inter8));
  nand2 gate836(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate837(.a(s_41), .b(gate219inter3), .O(gate219inter10));
  nor2  gate838(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate839(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate840(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1219(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1220(.a(gate228inter0), .b(s_96), .O(gate228inter1));
  and2  gate1221(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1222(.a(s_96), .O(gate228inter3));
  inv1  gate1223(.a(s_97), .O(gate228inter4));
  nand2 gate1224(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1225(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1226(.a(G696), .O(gate228inter7));
  inv1  gate1227(.a(G697), .O(gate228inter8));
  nand2 gate1228(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1229(.a(s_97), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1230(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1231(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1232(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1289(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1290(.a(gate238inter0), .b(s_106), .O(gate238inter1));
  and2  gate1291(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1292(.a(s_106), .O(gate238inter3));
  inv1  gate1293(.a(s_107), .O(gate238inter4));
  nand2 gate1294(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1295(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1296(.a(G257), .O(gate238inter7));
  inv1  gate1297(.a(G709), .O(gate238inter8));
  nand2 gate1298(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1299(.a(s_107), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1300(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1301(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1302(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1107(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1108(.a(gate243inter0), .b(s_80), .O(gate243inter1));
  and2  gate1109(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1110(.a(s_80), .O(gate243inter3));
  inv1  gate1111(.a(s_81), .O(gate243inter4));
  nand2 gate1112(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1113(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1114(.a(G245), .O(gate243inter7));
  inv1  gate1115(.a(G733), .O(gate243inter8));
  nand2 gate1116(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1117(.a(s_81), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1118(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1119(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1120(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate673(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate674(.a(gate245inter0), .b(s_18), .O(gate245inter1));
  and2  gate675(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate676(.a(s_18), .O(gate245inter3));
  inv1  gate677(.a(s_19), .O(gate245inter4));
  nand2 gate678(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate679(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate680(.a(G248), .O(gate245inter7));
  inv1  gate681(.a(G736), .O(gate245inter8));
  nand2 gate682(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate683(.a(s_19), .b(gate245inter3), .O(gate245inter10));
  nor2  gate684(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate685(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate686(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate603(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate604(.a(gate255inter0), .b(s_8), .O(gate255inter1));
  and2  gate605(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate606(.a(s_8), .O(gate255inter3));
  inv1  gate607(.a(s_9), .O(gate255inter4));
  nand2 gate608(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate609(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate610(.a(G263), .O(gate255inter7));
  inv1  gate611(.a(G751), .O(gate255inter8));
  nand2 gate612(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate613(.a(s_9), .b(gate255inter3), .O(gate255inter10));
  nor2  gate614(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate615(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate616(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1359(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1360(.a(gate276inter0), .b(s_116), .O(gate276inter1));
  and2  gate1361(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1362(.a(s_116), .O(gate276inter3));
  inv1  gate1363(.a(s_117), .O(gate276inter4));
  nand2 gate1364(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1365(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1366(.a(G773), .O(gate276inter7));
  inv1  gate1367(.a(G797), .O(gate276inter8));
  nand2 gate1368(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1369(.a(s_117), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1370(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1371(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1372(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1135(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1136(.a(gate277inter0), .b(s_84), .O(gate277inter1));
  and2  gate1137(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1138(.a(s_84), .O(gate277inter3));
  inv1  gate1139(.a(s_85), .O(gate277inter4));
  nand2 gate1140(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1141(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1142(.a(G648), .O(gate277inter7));
  inv1  gate1143(.a(G800), .O(gate277inter8));
  nand2 gate1144(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1145(.a(s_85), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1146(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1147(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1148(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1233(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1234(.a(gate282inter0), .b(s_98), .O(gate282inter1));
  and2  gate1235(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1236(.a(s_98), .O(gate282inter3));
  inv1  gate1237(.a(s_99), .O(gate282inter4));
  nand2 gate1238(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1239(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1240(.a(G782), .O(gate282inter7));
  inv1  gate1241(.a(G806), .O(gate282inter8));
  nand2 gate1242(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1243(.a(s_99), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1244(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1245(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1246(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate701(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate702(.a(gate284inter0), .b(s_22), .O(gate284inter1));
  and2  gate703(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate704(.a(s_22), .O(gate284inter3));
  inv1  gate705(.a(s_23), .O(gate284inter4));
  nand2 gate706(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate707(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate708(.a(G785), .O(gate284inter7));
  inv1  gate709(.a(G809), .O(gate284inter8));
  nand2 gate710(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate711(.a(s_23), .b(gate284inter3), .O(gate284inter10));
  nor2  gate712(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate713(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate714(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1275(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1276(.a(gate286inter0), .b(s_104), .O(gate286inter1));
  and2  gate1277(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1278(.a(s_104), .O(gate286inter3));
  inv1  gate1279(.a(s_105), .O(gate286inter4));
  nand2 gate1280(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1281(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1282(.a(G788), .O(gate286inter7));
  inv1  gate1283(.a(G812), .O(gate286inter8));
  nand2 gate1284(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1285(.a(s_105), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1286(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1287(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1288(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1345(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1346(.a(gate287inter0), .b(s_114), .O(gate287inter1));
  and2  gate1347(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1348(.a(s_114), .O(gate287inter3));
  inv1  gate1349(.a(s_115), .O(gate287inter4));
  nand2 gate1350(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1351(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1352(.a(G663), .O(gate287inter7));
  inv1  gate1353(.a(G815), .O(gate287inter8));
  nand2 gate1354(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1355(.a(s_115), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1356(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1357(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1358(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1373(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1374(.a(gate288inter0), .b(s_118), .O(gate288inter1));
  and2  gate1375(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1376(.a(s_118), .O(gate288inter3));
  inv1  gate1377(.a(s_119), .O(gate288inter4));
  nand2 gate1378(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1379(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1380(.a(G791), .O(gate288inter7));
  inv1  gate1381(.a(G815), .O(gate288inter8));
  nand2 gate1382(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1383(.a(s_119), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1384(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1385(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1386(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate757(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate758(.a(gate293inter0), .b(s_30), .O(gate293inter1));
  and2  gate759(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate760(.a(s_30), .O(gate293inter3));
  inv1  gate761(.a(s_31), .O(gate293inter4));
  nand2 gate762(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate763(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate764(.a(G828), .O(gate293inter7));
  inv1  gate765(.a(G829), .O(gate293inter8));
  nand2 gate766(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate767(.a(s_31), .b(gate293inter3), .O(gate293inter10));
  nor2  gate768(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate769(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate770(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1191(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1192(.a(gate296inter0), .b(s_92), .O(gate296inter1));
  and2  gate1193(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1194(.a(s_92), .O(gate296inter3));
  inv1  gate1195(.a(s_93), .O(gate296inter4));
  nand2 gate1196(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1197(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1198(.a(G826), .O(gate296inter7));
  inv1  gate1199(.a(G827), .O(gate296inter8));
  nand2 gate1200(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1201(.a(s_93), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1202(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1203(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1204(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1037(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1038(.a(gate387inter0), .b(s_70), .O(gate387inter1));
  and2  gate1039(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1040(.a(s_70), .O(gate387inter3));
  inv1  gate1041(.a(s_71), .O(gate387inter4));
  nand2 gate1042(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1043(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1044(.a(G1), .O(gate387inter7));
  inv1  gate1045(.a(G1036), .O(gate387inter8));
  nand2 gate1046(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1047(.a(s_71), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1048(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1049(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1050(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate785(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate786(.a(gate389inter0), .b(s_34), .O(gate389inter1));
  and2  gate787(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate788(.a(s_34), .O(gate389inter3));
  inv1  gate789(.a(s_35), .O(gate389inter4));
  nand2 gate790(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate791(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate792(.a(G3), .O(gate389inter7));
  inv1  gate793(.a(G1042), .O(gate389inter8));
  nand2 gate794(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate795(.a(s_35), .b(gate389inter3), .O(gate389inter10));
  nor2  gate796(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate797(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate798(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1457(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1458(.a(gate406inter0), .b(s_130), .O(gate406inter1));
  and2  gate1459(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1460(.a(s_130), .O(gate406inter3));
  inv1  gate1461(.a(s_131), .O(gate406inter4));
  nand2 gate1462(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1463(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1464(.a(G20), .O(gate406inter7));
  inv1  gate1465(.a(G1093), .O(gate406inter8));
  nand2 gate1466(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1467(.a(s_131), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1468(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1469(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1470(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1317(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1318(.a(gate412inter0), .b(s_110), .O(gate412inter1));
  and2  gate1319(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1320(.a(s_110), .O(gate412inter3));
  inv1  gate1321(.a(s_111), .O(gate412inter4));
  nand2 gate1322(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1323(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1324(.a(G26), .O(gate412inter7));
  inv1  gate1325(.a(G1111), .O(gate412inter8));
  nand2 gate1326(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1327(.a(s_111), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1328(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1329(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1330(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1429(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1430(.a(gate420inter0), .b(s_126), .O(gate420inter1));
  and2  gate1431(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1432(.a(s_126), .O(gate420inter3));
  inv1  gate1433(.a(s_127), .O(gate420inter4));
  nand2 gate1434(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1435(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1436(.a(G1036), .O(gate420inter7));
  inv1  gate1437(.a(G1132), .O(gate420inter8));
  nand2 gate1438(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1439(.a(s_127), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1440(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1441(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1442(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate547(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate548(.a(gate421inter0), .b(s_0), .O(gate421inter1));
  and2  gate549(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate550(.a(s_0), .O(gate421inter3));
  inv1  gate551(.a(s_1), .O(gate421inter4));
  nand2 gate552(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate553(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate554(.a(G2), .O(gate421inter7));
  inv1  gate555(.a(G1135), .O(gate421inter8));
  nand2 gate556(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate557(.a(s_1), .b(gate421inter3), .O(gate421inter10));
  nor2  gate558(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate559(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate560(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1513(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1514(.a(gate463inter0), .b(s_138), .O(gate463inter1));
  and2  gate1515(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1516(.a(s_138), .O(gate463inter3));
  inv1  gate1517(.a(s_139), .O(gate463inter4));
  nand2 gate1518(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1519(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1520(.a(G23), .O(gate463inter7));
  inv1  gate1521(.a(G1198), .O(gate463inter8));
  nand2 gate1522(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1523(.a(s_139), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1524(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1525(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1526(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1401(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1402(.a(gate465inter0), .b(s_122), .O(gate465inter1));
  and2  gate1403(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1404(.a(s_122), .O(gate465inter3));
  inv1  gate1405(.a(s_123), .O(gate465inter4));
  nand2 gate1406(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1407(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1408(.a(G24), .O(gate465inter7));
  inv1  gate1409(.a(G1201), .O(gate465inter8));
  nand2 gate1410(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1411(.a(s_123), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1412(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1413(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1414(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate995(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate996(.a(gate469inter0), .b(s_64), .O(gate469inter1));
  and2  gate997(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate998(.a(s_64), .O(gate469inter3));
  inv1  gate999(.a(s_65), .O(gate469inter4));
  nand2 gate1000(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1001(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1002(.a(G26), .O(gate469inter7));
  inv1  gate1003(.a(G1207), .O(gate469inter8));
  nand2 gate1004(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1005(.a(s_65), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1006(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1007(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1008(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate715(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate716(.a(gate472inter0), .b(s_24), .O(gate472inter1));
  and2  gate717(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate718(.a(s_24), .O(gate472inter3));
  inv1  gate719(.a(s_25), .O(gate472inter4));
  nand2 gate720(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate721(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate722(.a(G1114), .O(gate472inter7));
  inv1  gate723(.a(G1210), .O(gate472inter8));
  nand2 gate724(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate725(.a(s_25), .b(gate472inter3), .O(gate472inter10));
  nor2  gate726(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate727(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate728(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1079(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1080(.a(gate478inter0), .b(s_76), .O(gate478inter1));
  and2  gate1081(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1082(.a(s_76), .O(gate478inter3));
  inv1  gate1083(.a(s_77), .O(gate478inter4));
  nand2 gate1084(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1085(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1086(.a(G1123), .O(gate478inter7));
  inv1  gate1087(.a(G1219), .O(gate478inter8));
  nand2 gate1088(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1089(.a(s_77), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1090(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1091(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1092(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1149(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1150(.a(gate482inter0), .b(s_86), .O(gate482inter1));
  and2  gate1151(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1152(.a(s_86), .O(gate482inter3));
  inv1  gate1153(.a(s_87), .O(gate482inter4));
  nand2 gate1154(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1155(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1156(.a(G1129), .O(gate482inter7));
  inv1  gate1157(.a(G1225), .O(gate482inter8));
  nand2 gate1158(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1159(.a(s_87), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1160(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1161(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1162(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate911(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate912(.a(gate493inter0), .b(s_52), .O(gate493inter1));
  and2  gate913(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate914(.a(s_52), .O(gate493inter3));
  inv1  gate915(.a(s_53), .O(gate493inter4));
  nand2 gate916(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate917(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate918(.a(G1248), .O(gate493inter7));
  inv1  gate919(.a(G1249), .O(gate493inter8));
  nand2 gate920(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate921(.a(s_53), .b(gate493inter3), .O(gate493inter10));
  nor2  gate922(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate923(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate924(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1485(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1486(.a(gate502inter0), .b(s_134), .O(gate502inter1));
  and2  gate1487(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1488(.a(s_134), .O(gate502inter3));
  inv1  gate1489(.a(s_135), .O(gate502inter4));
  nand2 gate1490(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1491(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1492(.a(G1266), .O(gate502inter7));
  inv1  gate1493(.a(G1267), .O(gate502inter8));
  nand2 gate1494(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1495(.a(s_135), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1496(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1497(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1498(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1597(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1598(.a(gate503inter0), .b(s_150), .O(gate503inter1));
  and2  gate1599(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1600(.a(s_150), .O(gate503inter3));
  inv1  gate1601(.a(s_151), .O(gate503inter4));
  nand2 gate1602(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1603(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1604(.a(G1268), .O(gate503inter7));
  inv1  gate1605(.a(G1269), .O(gate503inter8));
  nand2 gate1606(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1607(.a(s_151), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1608(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1609(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1610(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate799(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate800(.a(gate504inter0), .b(s_36), .O(gate504inter1));
  and2  gate801(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate802(.a(s_36), .O(gate504inter3));
  inv1  gate803(.a(s_37), .O(gate504inter4));
  nand2 gate804(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate805(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate806(.a(G1270), .O(gate504inter7));
  inv1  gate807(.a(G1271), .O(gate504inter8));
  nand2 gate808(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate809(.a(s_37), .b(gate504inter3), .O(gate504inter10));
  nor2  gate810(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate811(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate812(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate743(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate744(.a(gate507inter0), .b(s_28), .O(gate507inter1));
  and2  gate745(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate746(.a(s_28), .O(gate507inter3));
  inv1  gate747(.a(s_29), .O(gate507inter4));
  nand2 gate748(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate749(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate750(.a(G1276), .O(gate507inter7));
  inv1  gate751(.a(G1277), .O(gate507inter8));
  nand2 gate752(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate753(.a(s_29), .b(gate507inter3), .O(gate507inter10));
  nor2  gate754(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate755(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate756(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate631(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate632(.a(gate510inter0), .b(s_12), .O(gate510inter1));
  and2  gate633(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate634(.a(s_12), .O(gate510inter3));
  inv1  gate635(.a(s_13), .O(gate510inter4));
  nand2 gate636(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate637(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate638(.a(G1282), .O(gate510inter7));
  inv1  gate639(.a(G1283), .O(gate510inter8));
  nand2 gate640(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate641(.a(s_13), .b(gate510inter3), .O(gate510inter10));
  nor2  gate642(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate643(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate644(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule