module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate497(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate498(.a(gate22inter0), .b(s_48), .O(gate22inter1));
  and2  gate499(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate500(.a(s_48), .O(gate22inter3));
  inv1  gate501(.a(s_49), .O(gate22inter4));
  nand2 gate502(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate503(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate504(.a(N122), .O(gate22inter7));
  inv1  gate505(.a(N17), .O(gate22inter8));
  nand2 gate506(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate507(.a(s_49), .b(gate22inter3), .O(gate22inter10));
  nor2  gate508(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate509(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate510(.a(gate22inter12), .b(gate22inter1), .O(N159));

  xor2  gate455(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate456(.a(gate23inter0), .b(s_42), .O(gate23inter1));
  and2  gate457(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate458(.a(s_42), .O(gate23inter3));
  inv1  gate459(.a(s_43), .O(gate23inter4));
  nand2 gate460(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate461(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate462(.a(N126), .O(gate23inter7));
  inv1  gate463(.a(N30), .O(gate23inter8));
  nand2 gate464(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate465(.a(s_43), .b(gate23inter3), .O(gate23inter10));
  nor2  gate466(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate467(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate468(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate189(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate190(.a(gate30inter0), .b(s_4), .O(gate30inter1));
  and2  gate191(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate192(.a(s_4), .O(gate30inter3));
  inv1  gate193(.a(s_5), .O(gate30inter4));
  nand2 gate194(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate195(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate196(.a(N21), .O(gate30inter7));
  inv1  gate197(.a(N123), .O(gate30inter8));
  nand2 gate198(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate199(.a(s_5), .b(gate30inter3), .O(gate30inter10));
  nor2  gate200(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate201(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate202(.a(gate30inter12), .b(gate30inter1), .O(N183));

  xor2  gate273(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate274(.a(gate31inter0), .b(s_16), .O(gate31inter1));
  and2  gate275(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate276(.a(s_16), .O(gate31inter3));
  inv1  gate277(.a(s_17), .O(gate31inter4));
  nand2 gate278(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate279(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate280(.a(N27), .O(gate31inter7));
  inv1  gate281(.a(N123), .O(gate31inter8));
  nand2 gate282(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate283(.a(s_17), .b(gate31inter3), .O(gate31inter10));
  nor2  gate284(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate285(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate286(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate413(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate414(.a(gate37inter0), .b(s_36), .O(gate37inter1));
  and2  gate415(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate416(.a(s_36), .O(gate37inter3));
  inv1  gate417(.a(s_37), .O(gate37inter4));
  nand2 gate418(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate419(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate420(.a(N66), .O(gate37inter7));
  inv1  gate421(.a(N135), .O(gate37inter8));
  nand2 gate422(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate423(.a(s_37), .b(gate37inter3), .O(gate37inter10));
  nor2  gate424(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate425(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate426(.a(gate37inter12), .b(gate37inter1), .O(N190));
nor2 gate38( .a(N73), .b(N139), .O(N191) );

  xor2  gate469(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate470(.a(gate39inter0), .b(s_44), .O(gate39inter1));
  and2  gate471(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate472(.a(s_44), .O(gate39inter3));
  inv1  gate473(.a(s_45), .O(gate39inter4));
  nand2 gate474(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate475(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate476(.a(N79), .O(gate39inter7));
  inv1  gate477(.a(N139), .O(gate39inter8));
  nand2 gate478(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate479(.a(s_45), .b(gate39inter3), .O(gate39inter10));
  nor2  gate480(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate481(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate482(.a(gate39inter12), .b(gate39inter1), .O(N192));
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate343(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate344(.a(gate41inter0), .b(s_26), .O(gate41inter1));
  and2  gate345(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate346(.a(s_26), .O(gate41inter3));
  inv1  gate347(.a(s_27), .O(gate41inter4));
  nand2 gate348(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate349(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate350(.a(N92), .O(gate41inter7));
  inv1  gate351(.a(N143), .O(gate41inter8));
  nand2 gate352(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate353(.a(s_27), .b(gate41inter3), .O(gate41inter10));
  nor2  gate354(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate355(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate356(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate301(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate302(.a(gate60inter0), .b(s_20), .O(gate60inter1));
  and2  gate303(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate304(.a(s_20), .O(gate60inter3));
  inv1  gate305(.a(s_21), .O(gate60inter4));
  nand2 gate306(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate307(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate308(.a(N213), .O(gate60inter7));
  inv1  gate309(.a(N24), .O(gate60inter8));
  nand2 gate310(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate311(.a(s_21), .b(gate60inter3), .O(gate60inter10));
  nor2  gate312(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate313(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate314(.a(gate60inter12), .b(gate60inter1), .O(N250));
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );

  xor2  gate175(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate176(.a(gate63inter0), .b(s_2), .O(gate63inter1));
  and2  gate177(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate178(.a(s_2), .O(gate63inter3));
  inv1  gate179(.a(s_3), .O(gate63inter4));
  nand2 gate180(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate181(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate182(.a(N213), .O(gate63inter7));
  inv1  gate183(.a(N50), .O(gate63inter8));
  nand2 gate184(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate185(.a(s_3), .b(gate63inter3), .O(gate63inter10));
  nor2  gate186(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate187(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate188(.a(gate63inter12), .b(gate63inter1), .O(N255));
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate511(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate512(.a(gate65inter0), .b(s_50), .O(gate65inter1));
  and2  gate513(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate514(.a(s_50), .O(gate65inter3));
  inv1  gate515(.a(s_51), .O(gate65inter4));
  nand2 gate516(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate517(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate518(.a(N213), .O(gate65inter7));
  inv1  gate519(.a(N76), .O(gate65inter8));
  nand2 gate520(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate521(.a(s_51), .b(gate65inter3), .O(gate65inter10));
  nor2  gate522(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate523(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate524(.a(gate65inter12), .b(gate65inter1), .O(N257));

  xor2  gate203(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate204(.a(gate66inter0), .b(s_6), .O(gate66inter1));
  and2  gate205(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate206(.a(s_6), .O(gate66inter3));
  inv1  gate207(.a(s_7), .O(gate66inter4));
  nand2 gate208(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate209(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate210(.a(N213), .O(gate66inter7));
  inv1  gate211(.a(N89), .O(gate66inter8));
  nand2 gate212(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate213(.a(s_7), .b(gate66inter3), .O(gate66inter10));
  nor2  gate214(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate215(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate216(.a(gate66inter12), .b(gate66inter1), .O(N258));
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate161(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate162(.a(gate75inter0), .b(s_0), .O(gate75inter1));
  and2  gate163(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate164(.a(s_0), .O(gate75inter3));
  inv1  gate165(.a(s_1), .O(gate75inter4));
  nand2 gate166(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate167(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate168(.a(N243), .O(gate75inter7));
  inv1  gate169(.a(N193), .O(gate75inter8));
  nand2 gate170(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate171(.a(s_1), .b(gate75inter3), .O(gate75inter10));
  nor2  gate172(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate173(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate174(.a(gate75inter12), .b(gate75inter1), .O(N279));

  xor2  gate441(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate442(.a(gate76inter0), .b(s_40), .O(gate76inter1));
  and2  gate443(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate444(.a(s_40), .O(gate76inter3));
  inv1  gate445(.a(s_41), .O(gate76inter4));
  nand2 gate446(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate447(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate448(.a(N247), .O(gate76inter7));
  inv1  gate449(.a(N195), .O(gate76inter8));
  nand2 gate450(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate451(.a(s_41), .b(gate76inter3), .O(gate76inter10));
  nor2  gate452(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate453(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate454(.a(gate76inter12), .b(gate76inter1), .O(N282));
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate231(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate232(.a(gate80inter0), .b(s_10), .O(gate80inter1));
  and2  gate233(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate234(.a(s_10), .O(gate80inter3));
  inv1  gate235(.a(s_11), .O(gate80inter4));
  nand2 gate236(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate237(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate238(.a(N233), .O(gate80inter7));
  inv1  gate239(.a(N188), .O(gate80inter8));
  nand2 gate240(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate241(.a(s_11), .b(gate80inter3), .O(gate80inter10));
  nor2  gate242(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate243(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate244(.a(gate80inter12), .b(gate80inter1), .O(N290));

  xor2  gate357(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate358(.a(gate81inter0), .b(s_28), .O(gate81inter1));
  and2  gate359(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate360(.a(s_28), .O(gate81inter3));
  inv1  gate361(.a(s_29), .O(gate81inter4));
  nand2 gate362(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate363(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate364(.a(N236), .O(gate81inter7));
  inv1  gate365(.a(N190), .O(gate81inter8));
  nand2 gate366(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate367(.a(s_29), .b(gate81inter3), .O(gate81inter10));
  nor2  gate368(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate369(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate370(.a(gate81inter12), .b(gate81inter1), .O(N291));
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );

  xor2  gate483(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate484(.a(gate85inter0), .b(s_46), .O(gate85inter1));
  and2  gate485(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate486(.a(s_46), .O(gate85inter3));
  inv1  gate487(.a(s_47), .O(gate85inter4));
  nand2 gate488(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate489(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate490(.a(N251), .O(gate85inter7));
  inv1  gate491(.a(N198), .O(gate85inter8));
  nand2 gate492(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate493(.a(s_47), .b(gate85inter3), .O(gate85inter10));
  nor2  gate494(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate495(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate496(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate385(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate386(.a(gate99inter0), .b(s_32), .O(gate99inter1));
  and2  gate387(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate388(.a(s_32), .O(gate99inter3));
  inv1  gate389(.a(s_33), .O(gate99inter4));
  nand2 gate390(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate391(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate392(.a(N309), .O(gate99inter7));
  inv1  gate393(.a(N260), .O(gate99inter8));
  nand2 gate394(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate395(.a(s_33), .b(gate99inter3), .O(gate99inter10));
  nor2  gate396(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate397(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate398(.a(gate99inter12), .b(gate99inter1), .O(N330));
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );

  xor2  gate399(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate400(.a(gate104inter0), .b(s_34), .O(gate104inter1));
  and2  gate401(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate402(.a(s_34), .O(gate104inter3));
  inv1  gate403(.a(s_35), .O(gate104inter4));
  nand2 gate404(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate405(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate406(.a(N309), .O(gate104inter7));
  inv1  gate407(.a(N273), .O(gate104inter8));
  nand2 gate408(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate409(.a(s_35), .b(gate104inter3), .O(gate104inter10));
  nor2  gate410(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate411(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate412(.a(gate104inter12), .b(gate104inter1), .O(N335));
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate287(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate288(.a(gate110inter0), .b(s_18), .O(gate110inter1));
  and2  gate289(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate290(.a(s_18), .O(gate110inter3));
  inv1  gate291(.a(s_19), .O(gate110inter4));
  nand2 gate292(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate293(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate294(.a(N309), .O(gate110inter7));
  inv1  gate295(.a(N282), .O(gate110inter8));
  nand2 gate296(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate297(.a(s_19), .b(gate110inter3), .O(gate110inter10));
  nor2  gate298(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate299(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate300(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate427(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate428(.a(gate113inter0), .b(s_38), .O(gate113inter1));
  and2  gate429(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate430(.a(s_38), .O(gate113inter3));
  inv1  gate431(.a(s_39), .O(gate113inter4));
  nand2 gate432(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate433(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate434(.a(N319), .O(gate113inter7));
  inv1  gate435(.a(N73), .O(gate113inter8));
  nand2 gate436(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate437(.a(s_39), .b(gate113inter3), .O(gate113inter10));
  nor2  gate438(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate439(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate440(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );

  xor2  gate245(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate246(.a(gate116inter0), .b(s_12), .O(gate116inter1));
  and2  gate247(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate248(.a(s_12), .O(gate116inter3));
  inv1  gate249(.a(s_13), .O(gate116inter4));
  nand2 gate250(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate251(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate252(.a(N319), .O(gate116inter7));
  inv1  gate253(.a(N112), .O(gate116inter8));
  nand2 gate254(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate255(.a(s_13), .b(gate116inter3), .O(gate116inter10));
  nor2  gate256(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate257(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate258(.a(gate116inter12), .b(gate116inter1), .O(N347));
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate371(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate372(.a(gate118inter0), .b(s_30), .O(gate118inter1));
  and2  gate373(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate374(.a(s_30), .O(gate118inter3));
  inv1  gate375(.a(s_31), .O(gate118inter4));
  nand2 gate376(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate377(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate378(.a(N331), .O(gate118inter7));
  inv1  gate379(.a(N301), .O(gate118inter8));
  nand2 gate380(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate381(.a(s_31), .b(gate118inter3), .O(gate118inter10));
  nor2  gate382(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate383(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate384(.a(gate118inter12), .b(gate118inter1), .O(N349));

  xor2  gate259(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate260(.a(gate119inter0), .b(s_14), .O(gate119inter1));
  and2  gate261(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate262(.a(s_14), .O(gate119inter3));
  inv1  gate263(.a(s_15), .O(gate119inter4));
  nand2 gate264(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate265(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate266(.a(N332), .O(gate119inter7));
  inv1  gate267(.a(N302), .O(gate119inter8));
  nand2 gate268(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate269(.a(s_15), .b(gate119inter3), .O(gate119inter10));
  nor2  gate270(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate271(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate272(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate315(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate316(.a(gate121inter0), .b(s_22), .O(gate121inter1));
  and2  gate317(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate318(.a(s_22), .O(gate121inter3));
  inv1  gate319(.a(s_23), .O(gate121inter4));
  nand2 gate320(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate321(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate322(.a(N335), .O(gate121inter7));
  inv1  gate323(.a(N304), .O(gate121inter8));
  nand2 gate324(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate325(.a(s_23), .b(gate121inter3), .O(gate121inter10));
  nor2  gate326(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate327(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate328(.a(gate121inter12), .b(gate121inter1), .O(N352));
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );

  xor2  gate329(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate330(.a(gate124inter0), .b(s_24), .O(gate124inter1));
  and2  gate331(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate332(.a(s_24), .O(gate124inter3));
  inv1  gate333(.a(s_25), .O(gate124inter4));
  nand2 gate334(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate335(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate336(.a(N341), .O(gate124inter7));
  inv1  gate337(.a(N307), .O(gate124inter8));
  nand2 gate338(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate339(.a(s_25), .b(gate124inter3), .O(gate124inter10));
  nor2  gate340(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate341(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate342(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate217(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate218(.a(gate136inter0), .b(s_8), .O(gate136inter1));
  and2  gate219(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate220(.a(s_8), .O(gate136inter3));
  inv1  gate221(.a(s_9), .O(gate136inter4));
  nand2 gate222(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate223(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate224(.a(N360), .O(gate136inter7));
  inv1  gate225(.a(N105), .O(gate136inter8));
  nand2 gate226(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate227(.a(s_9), .b(gate136inter3), .O(gate136inter10));
  nor2  gate228(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate229(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate230(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule