module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate883(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate884(.a(gate9inter0), .b(s_48), .O(gate9inter1));
  and2  gate885(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate886(.a(s_48), .O(gate9inter3));
  inv1  gate887(.a(s_49), .O(gate9inter4));
  nand2 gate888(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate889(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate890(.a(G1), .O(gate9inter7));
  inv1  gate891(.a(G2), .O(gate9inter8));
  nand2 gate892(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate893(.a(s_49), .b(gate9inter3), .O(gate9inter10));
  nor2  gate894(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate895(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate896(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1177(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1178(.a(gate11inter0), .b(s_90), .O(gate11inter1));
  and2  gate1179(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1180(.a(s_90), .O(gate11inter3));
  inv1  gate1181(.a(s_91), .O(gate11inter4));
  nand2 gate1182(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1183(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1184(.a(G5), .O(gate11inter7));
  inv1  gate1185(.a(G6), .O(gate11inter8));
  nand2 gate1186(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1187(.a(s_91), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1188(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1189(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1190(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2017(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2018(.a(gate13inter0), .b(s_210), .O(gate13inter1));
  and2  gate2019(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2020(.a(s_210), .O(gate13inter3));
  inv1  gate2021(.a(s_211), .O(gate13inter4));
  nand2 gate2022(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2023(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2024(.a(G9), .O(gate13inter7));
  inv1  gate2025(.a(G10), .O(gate13inter8));
  nand2 gate2026(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2027(.a(s_211), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2028(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2029(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2030(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1807(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1808(.a(gate14inter0), .b(s_180), .O(gate14inter1));
  and2  gate1809(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1810(.a(s_180), .O(gate14inter3));
  inv1  gate1811(.a(s_181), .O(gate14inter4));
  nand2 gate1812(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1813(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1814(.a(G11), .O(gate14inter7));
  inv1  gate1815(.a(G12), .O(gate14inter8));
  nand2 gate1816(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1817(.a(s_181), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1818(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1819(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1820(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1975(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1976(.a(gate28inter0), .b(s_204), .O(gate28inter1));
  and2  gate1977(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1978(.a(s_204), .O(gate28inter3));
  inv1  gate1979(.a(s_205), .O(gate28inter4));
  nand2 gate1980(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1981(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1982(.a(G10), .O(gate28inter7));
  inv1  gate1983(.a(G14), .O(gate28inter8));
  nand2 gate1984(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1985(.a(s_205), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1986(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1987(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1988(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1695(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1696(.a(gate31inter0), .b(s_164), .O(gate31inter1));
  and2  gate1697(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1698(.a(s_164), .O(gate31inter3));
  inv1  gate1699(.a(s_165), .O(gate31inter4));
  nand2 gate1700(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1701(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1702(.a(G4), .O(gate31inter7));
  inv1  gate1703(.a(G8), .O(gate31inter8));
  nand2 gate1704(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1705(.a(s_165), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1706(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1707(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1708(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1233(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1234(.a(gate34inter0), .b(s_98), .O(gate34inter1));
  and2  gate1235(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1236(.a(s_98), .O(gate34inter3));
  inv1  gate1237(.a(s_99), .O(gate34inter4));
  nand2 gate1238(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1239(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1240(.a(G25), .O(gate34inter7));
  inv1  gate1241(.a(G29), .O(gate34inter8));
  nand2 gate1242(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1243(.a(s_99), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1244(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1245(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1246(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2045(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2046(.a(gate36inter0), .b(s_214), .O(gate36inter1));
  and2  gate2047(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2048(.a(s_214), .O(gate36inter3));
  inv1  gate2049(.a(s_215), .O(gate36inter4));
  nand2 gate2050(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2051(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2052(.a(G26), .O(gate36inter7));
  inv1  gate2053(.a(G30), .O(gate36inter8));
  nand2 gate2054(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2055(.a(s_215), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2056(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2057(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2058(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate799(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate800(.a(gate38inter0), .b(s_36), .O(gate38inter1));
  and2  gate801(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate802(.a(s_36), .O(gate38inter3));
  inv1  gate803(.a(s_37), .O(gate38inter4));
  nand2 gate804(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate805(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate806(.a(G27), .O(gate38inter7));
  inv1  gate807(.a(G31), .O(gate38inter8));
  nand2 gate808(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate809(.a(s_37), .b(gate38inter3), .O(gate38inter10));
  nor2  gate810(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate811(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate812(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1107(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1108(.a(gate43inter0), .b(s_80), .O(gate43inter1));
  and2  gate1109(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1110(.a(s_80), .O(gate43inter3));
  inv1  gate1111(.a(s_81), .O(gate43inter4));
  nand2 gate1112(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1113(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1114(.a(G3), .O(gate43inter7));
  inv1  gate1115(.a(G269), .O(gate43inter8));
  nand2 gate1116(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1117(.a(s_81), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1118(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1119(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1120(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate631(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate632(.a(gate45inter0), .b(s_12), .O(gate45inter1));
  and2  gate633(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate634(.a(s_12), .O(gate45inter3));
  inv1  gate635(.a(s_13), .O(gate45inter4));
  nand2 gate636(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate637(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate638(.a(G5), .O(gate45inter7));
  inv1  gate639(.a(G272), .O(gate45inter8));
  nand2 gate640(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate641(.a(s_13), .b(gate45inter3), .O(gate45inter10));
  nor2  gate642(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate643(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate644(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate603(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate604(.a(gate47inter0), .b(s_8), .O(gate47inter1));
  and2  gate605(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate606(.a(s_8), .O(gate47inter3));
  inv1  gate607(.a(s_9), .O(gate47inter4));
  nand2 gate608(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate609(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate610(.a(G7), .O(gate47inter7));
  inv1  gate611(.a(G275), .O(gate47inter8));
  nand2 gate612(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate613(.a(s_9), .b(gate47inter3), .O(gate47inter10));
  nor2  gate614(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate615(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate616(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2087(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2088(.a(gate59inter0), .b(s_220), .O(gate59inter1));
  and2  gate2089(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2090(.a(s_220), .O(gate59inter3));
  inv1  gate2091(.a(s_221), .O(gate59inter4));
  nand2 gate2092(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2093(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2094(.a(G19), .O(gate59inter7));
  inv1  gate2095(.a(G293), .O(gate59inter8));
  nand2 gate2096(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2097(.a(s_221), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2098(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2099(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2100(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate2185(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2186(.a(gate60inter0), .b(s_234), .O(gate60inter1));
  and2  gate2187(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2188(.a(s_234), .O(gate60inter3));
  inv1  gate2189(.a(s_235), .O(gate60inter4));
  nand2 gate2190(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2191(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2192(.a(G20), .O(gate60inter7));
  inv1  gate2193(.a(G293), .O(gate60inter8));
  nand2 gate2194(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2195(.a(s_235), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2196(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2197(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2198(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate897(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate898(.a(gate63inter0), .b(s_50), .O(gate63inter1));
  and2  gate899(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate900(.a(s_50), .O(gate63inter3));
  inv1  gate901(.a(s_51), .O(gate63inter4));
  nand2 gate902(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate903(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate904(.a(G23), .O(gate63inter7));
  inv1  gate905(.a(G299), .O(gate63inter8));
  nand2 gate906(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate907(.a(s_51), .b(gate63inter3), .O(gate63inter10));
  nor2  gate908(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate909(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate910(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1037(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1038(.a(gate64inter0), .b(s_70), .O(gate64inter1));
  and2  gate1039(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1040(.a(s_70), .O(gate64inter3));
  inv1  gate1041(.a(s_71), .O(gate64inter4));
  nand2 gate1042(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1043(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1044(.a(G24), .O(gate64inter7));
  inv1  gate1045(.a(G299), .O(gate64inter8));
  nand2 gate1046(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1047(.a(s_71), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1048(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1049(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1050(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1149(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1150(.a(gate66inter0), .b(s_86), .O(gate66inter1));
  and2  gate1151(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1152(.a(s_86), .O(gate66inter3));
  inv1  gate1153(.a(s_87), .O(gate66inter4));
  nand2 gate1154(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1155(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1156(.a(G26), .O(gate66inter7));
  inv1  gate1157(.a(G302), .O(gate66inter8));
  nand2 gate1158(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1159(.a(s_87), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1160(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1161(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1162(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1023(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1024(.a(gate69inter0), .b(s_68), .O(gate69inter1));
  and2  gate1025(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1026(.a(s_68), .O(gate69inter3));
  inv1  gate1027(.a(s_69), .O(gate69inter4));
  nand2 gate1028(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1029(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1030(.a(G29), .O(gate69inter7));
  inv1  gate1031(.a(G308), .O(gate69inter8));
  nand2 gate1032(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1033(.a(s_69), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1034(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1035(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1036(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2115(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2116(.a(gate77inter0), .b(s_224), .O(gate77inter1));
  and2  gate2117(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2118(.a(s_224), .O(gate77inter3));
  inv1  gate2119(.a(s_225), .O(gate77inter4));
  nand2 gate2120(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2121(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2122(.a(G2), .O(gate77inter7));
  inv1  gate2123(.a(G320), .O(gate77inter8));
  nand2 gate2124(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2125(.a(s_225), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2126(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2127(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2128(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1905(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1906(.a(gate80inter0), .b(s_194), .O(gate80inter1));
  and2  gate1907(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1908(.a(s_194), .O(gate80inter3));
  inv1  gate1909(.a(s_195), .O(gate80inter4));
  nand2 gate1910(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1911(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1912(.a(G14), .O(gate80inter7));
  inv1  gate1913(.a(G323), .O(gate80inter8));
  nand2 gate1914(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1915(.a(s_195), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1916(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1917(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1918(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2227(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2228(.a(gate81inter0), .b(s_240), .O(gate81inter1));
  and2  gate2229(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2230(.a(s_240), .O(gate81inter3));
  inv1  gate2231(.a(s_241), .O(gate81inter4));
  nand2 gate2232(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2233(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2234(.a(G3), .O(gate81inter7));
  inv1  gate2235(.a(G326), .O(gate81inter8));
  nand2 gate2236(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2237(.a(s_241), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2238(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2239(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2240(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate617(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate618(.a(gate87inter0), .b(s_10), .O(gate87inter1));
  and2  gate619(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate620(.a(s_10), .O(gate87inter3));
  inv1  gate621(.a(s_11), .O(gate87inter4));
  nand2 gate622(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate623(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate624(.a(G12), .O(gate87inter7));
  inv1  gate625(.a(G335), .O(gate87inter8));
  nand2 gate626(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate627(.a(s_11), .b(gate87inter3), .O(gate87inter10));
  nor2  gate628(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate629(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate630(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1737(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1738(.a(gate88inter0), .b(s_170), .O(gate88inter1));
  and2  gate1739(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1740(.a(s_170), .O(gate88inter3));
  inv1  gate1741(.a(s_171), .O(gate88inter4));
  nand2 gate1742(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1743(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1744(.a(G16), .O(gate88inter7));
  inv1  gate1745(.a(G335), .O(gate88inter8));
  nand2 gate1746(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1747(.a(s_171), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1748(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1749(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1750(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2073(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2074(.a(gate89inter0), .b(s_218), .O(gate89inter1));
  and2  gate2075(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2076(.a(s_218), .O(gate89inter3));
  inv1  gate2077(.a(s_219), .O(gate89inter4));
  nand2 gate2078(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2079(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2080(.a(G17), .O(gate89inter7));
  inv1  gate2081(.a(G338), .O(gate89inter8));
  nand2 gate2082(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2083(.a(s_219), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2084(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2085(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2086(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1989(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1990(.a(gate91inter0), .b(s_206), .O(gate91inter1));
  and2  gate1991(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1992(.a(s_206), .O(gate91inter3));
  inv1  gate1993(.a(s_207), .O(gate91inter4));
  nand2 gate1994(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1995(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1996(.a(G25), .O(gate91inter7));
  inv1  gate1997(.a(G341), .O(gate91inter8));
  nand2 gate1998(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1999(.a(s_207), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2000(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2001(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2002(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1471(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1472(.a(gate92inter0), .b(s_132), .O(gate92inter1));
  and2  gate1473(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1474(.a(s_132), .O(gate92inter3));
  inv1  gate1475(.a(s_133), .O(gate92inter4));
  nand2 gate1476(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1477(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1478(.a(G29), .O(gate92inter7));
  inv1  gate1479(.a(G341), .O(gate92inter8));
  nand2 gate1480(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1481(.a(s_133), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1482(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1483(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1484(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1205(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1206(.a(gate93inter0), .b(s_94), .O(gate93inter1));
  and2  gate1207(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1208(.a(s_94), .O(gate93inter3));
  inv1  gate1209(.a(s_95), .O(gate93inter4));
  nand2 gate1210(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1211(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1212(.a(G18), .O(gate93inter7));
  inv1  gate1213(.a(G344), .O(gate93inter8));
  nand2 gate1214(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1215(.a(s_95), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1216(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1217(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1218(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1555(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1556(.a(gate96inter0), .b(s_144), .O(gate96inter1));
  and2  gate1557(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1558(.a(s_144), .O(gate96inter3));
  inv1  gate1559(.a(s_145), .O(gate96inter4));
  nand2 gate1560(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1561(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1562(.a(G30), .O(gate96inter7));
  inv1  gate1563(.a(G347), .O(gate96inter8));
  nand2 gate1564(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1565(.a(s_145), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1566(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1567(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1568(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate729(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate730(.a(gate99inter0), .b(s_26), .O(gate99inter1));
  and2  gate731(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate732(.a(s_26), .O(gate99inter3));
  inv1  gate733(.a(s_27), .O(gate99inter4));
  nand2 gate734(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate735(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate736(.a(G27), .O(gate99inter7));
  inv1  gate737(.a(G353), .O(gate99inter8));
  nand2 gate738(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate739(.a(s_27), .b(gate99inter3), .O(gate99inter10));
  nor2  gate740(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate741(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate742(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate911(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate912(.a(gate118inter0), .b(s_52), .O(gate118inter1));
  and2  gate913(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate914(.a(s_52), .O(gate118inter3));
  inv1  gate915(.a(s_53), .O(gate118inter4));
  nand2 gate916(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate917(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate918(.a(G388), .O(gate118inter7));
  inv1  gate919(.a(G389), .O(gate118inter8));
  nand2 gate920(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate921(.a(s_53), .b(gate118inter3), .O(gate118inter10));
  nor2  gate922(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate923(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate924(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1009(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1010(.a(gate126inter0), .b(s_66), .O(gate126inter1));
  and2  gate1011(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1012(.a(s_66), .O(gate126inter3));
  inv1  gate1013(.a(s_67), .O(gate126inter4));
  nand2 gate1014(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1015(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1016(.a(G404), .O(gate126inter7));
  inv1  gate1017(.a(G405), .O(gate126inter8));
  nand2 gate1018(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1019(.a(s_67), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1020(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1021(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1022(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1275(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1276(.a(gate129inter0), .b(s_104), .O(gate129inter1));
  and2  gate1277(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1278(.a(s_104), .O(gate129inter3));
  inv1  gate1279(.a(s_105), .O(gate129inter4));
  nand2 gate1280(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1281(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1282(.a(G410), .O(gate129inter7));
  inv1  gate1283(.a(G411), .O(gate129inter8));
  nand2 gate1284(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1285(.a(s_105), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1286(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1287(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1288(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate981(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate982(.a(gate131inter0), .b(s_62), .O(gate131inter1));
  and2  gate983(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate984(.a(s_62), .O(gate131inter3));
  inv1  gate985(.a(s_63), .O(gate131inter4));
  nand2 gate986(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate987(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate988(.a(G414), .O(gate131inter7));
  inv1  gate989(.a(G415), .O(gate131inter8));
  nand2 gate990(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate991(.a(s_63), .b(gate131inter3), .O(gate131inter10));
  nor2  gate992(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate993(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate994(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate715(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate716(.a(gate133inter0), .b(s_24), .O(gate133inter1));
  and2  gate717(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate718(.a(s_24), .O(gate133inter3));
  inv1  gate719(.a(s_25), .O(gate133inter4));
  nand2 gate720(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate721(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate722(.a(G418), .O(gate133inter7));
  inv1  gate723(.a(G419), .O(gate133inter8));
  nand2 gate724(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate725(.a(s_25), .b(gate133inter3), .O(gate133inter10));
  nor2  gate726(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate727(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate728(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1569(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1570(.a(gate134inter0), .b(s_146), .O(gate134inter1));
  and2  gate1571(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1572(.a(s_146), .O(gate134inter3));
  inv1  gate1573(.a(s_147), .O(gate134inter4));
  nand2 gate1574(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1575(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1576(.a(G420), .O(gate134inter7));
  inv1  gate1577(.a(G421), .O(gate134inter8));
  nand2 gate1578(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1579(.a(s_147), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1580(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1581(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1582(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2143(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2144(.a(gate135inter0), .b(s_228), .O(gate135inter1));
  and2  gate2145(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2146(.a(s_228), .O(gate135inter3));
  inv1  gate2147(.a(s_229), .O(gate135inter4));
  nand2 gate2148(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2149(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2150(.a(G422), .O(gate135inter7));
  inv1  gate2151(.a(G423), .O(gate135inter8));
  nand2 gate2152(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2153(.a(s_229), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2154(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2155(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2156(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate967(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate968(.a(gate141inter0), .b(s_60), .O(gate141inter1));
  and2  gate969(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate970(.a(s_60), .O(gate141inter3));
  inv1  gate971(.a(s_61), .O(gate141inter4));
  nand2 gate972(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate973(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate974(.a(G450), .O(gate141inter7));
  inv1  gate975(.a(G453), .O(gate141inter8));
  nand2 gate976(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate977(.a(s_61), .b(gate141inter3), .O(gate141inter10));
  nor2  gate978(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate979(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate980(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate925(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate926(.a(gate142inter0), .b(s_54), .O(gate142inter1));
  and2  gate927(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate928(.a(s_54), .O(gate142inter3));
  inv1  gate929(.a(s_55), .O(gate142inter4));
  nand2 gate930(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate931(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate932(.a(G456), .O(gate142inter7));
  inv1  gate933(.a(G459), .O(gate142inter8));
  nand2 gate934(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate935(.a(s_55), .b(gate142inter3), .O(gate142inter10));
  nor2  gate936(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate937(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate938(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1317(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1318(.a(gate147inter0), .b(s_110), .O(gate147inter1));
  and2  gate1319(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1320(.a(s_110), .O(gate147inter3));
  inv1  gate1321(.a(s_111), .O(gate147inter4));
  nand2 gate1322(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1323(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1324(.a(G486), .O(gate147inter7));
  inv1  gate1325(.a(G489), .O(gate147inter8));
  nand2 gate1326(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1327(.a(s_111), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1328(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1329(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1330(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1191(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1192(.a(gate148inter0), .b(s_92), .O(gate148inter1));
  and2  gate1193(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1194(.a(s_92), .O(gate148inter3));
  inv1  gate1195(.a(s_93), .O(gate148inter4));
  nand2 gate1196(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1197(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1198(.a(G492), .O(gate148inter7));
  inv1  gate1199(.a(G495), .O(gate148inter8));
  nand2 gate1200(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1201(.a(s_93), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1202(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1203(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1204(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate2171(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2172(.a(gate149inter0), .b(s_232), .O(gate149inter1));
  and2  gate2173(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2174(.a(s_232), .O(gate149inter3));
  inv1  gate2175(.a(s_233), .O(gate149inter4));
  nand2 gate2176(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2177(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2178(.a(G498), .O(gate149inter7));
  inv1  gate2179(.a(G501), .O(gate149inter8));
  nand2 gate2180(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2181(.a(s_233), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2182(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2183(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2184(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1051(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1052(.a(gate152inter0), .b(s_72), .O(gate152inter1));
  and2  gate1053(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1054(.a(s_72), .O(gate152inter3));
  inv1  gate1055(.a(s_73), .O(gate152inter4));
  nand2 gate1056(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1057(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1058(.a(G516), .O(gate152inter7));
  inv1  gate1059(.a(G519), .O(gate152inter8));
  nand2 gate1060(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1061(.a(s_73), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1062(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1063(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1064(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate813(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate814(.a(gate159inter0), .b(s_38), .O(gate159inter1));
  and2  gate815(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate816(.a(s_38), .O(gate159inter3));
  inv1  gate817(.a(s_39), .O(gate159inter4));
  nand2 gate818(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate819(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate820(.a(G444), .O(gate159inter7));
  inv1  gate821(.a(G531), .O(gate159inter8));
  nand2 gate822(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate823(.a(s_39), .b(gate159inter3), .O(gate159inter10));
  nor2  gate824(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate825(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate826(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1429(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1430(.a(gate161inter0), .b(s_126), .O(gate161inter1));
  and2  gate1431(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1432(.a(s_126), .O(gate161inter3));
  inv1  gate1433(.a(s_127), .O(gate161inter4));
  nand2 gate1434(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1435(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1436(.a(G450), .O(gate161inter7));
  inv1  gate1437(.a(G534), .O(gate161inter8));
  nand2 gate1438(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1439(.a(s_127), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1440(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1441(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1442(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1387(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1388(.a(gate162inter0), .b(s_120), .O(gate162inter1));
  and2  gate1389(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1390(.a(s_120), .O(gate162inter3));
  inv1  gate1391(.a(s_121), .O(gate162inter4));
  nand2 gate1392(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1393(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1394(.a(G453), .O(gate162inter7));
  inv1  gate1395(.a(G534), .O(gate162inter8));
  nand2 gate1396(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1397(.a(s_121), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1398(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1399(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1400(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate1247(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1248(.a(gate163inter0), .b(s_100), .O(gate163inter1));
  and2  gate1249(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1250(.a(s_100), .O(gate163inter3));
  inv1  gate1251(.a(s_101), .O(gate163inter4));
  nand2 gate1252(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1253(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1254(.a(G456), .O(gate163inter7));
  inv1  gate1255(.a(G537), .O(gate163inter8));
  nand2 gate1256(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1257(.a(s_101), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1258(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1259(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1260(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2101(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2102(.a(gate165inter0), .b(s_222), .O(gate165inter1));
  and2  gate2103(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2104(.a(s_222), .O(gate165inter3));
  inv1  gate2105(.a(s_223), .O(gate165inter4));
  nand2 gate2106(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2107(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2108(.a(G462), .O(gate165inter7));
  inv1  gate2109(.a(G540), .O(gate165inter8));
  nand2 gate2110(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2111(.a(s_223), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2112(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2113(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2114(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate953(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate954(.a(gate166inter0), .b(s_58), .O(gate166inter1));
  and2  gate955(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate956(.a(s_58), .O(gate166inter3));
  inv1  gate957(.a(s_59), .O(gate166inter4));
  nand2 gate958(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate959(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate960(.a(G465), .O(gate166inter7));
  inv1  gate961(.a(G540), .O(gate166inter8));
  nand2 gate962(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate963(.a(s_59), .b(gate166inter3), .O(gate166inter10));
  nor2  gate964(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate965(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate966(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1079(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1080(.a(gate169inter0), .b(s_76), .O(gate169inter1));
  and2  gate1081(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1082(.a(s_76), .O(gate169inter3));
  inv1  gate1083(.a(s_77), .O(gate169inter4));
  nand2 gate1084(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1085(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1086(.a(G474), .O(gate169inter7));
  inv1  gate1087(.a(G546), .O(gate169inter8));
  nand2 gate1088(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1089(.a(s_77), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1090(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1091(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1092(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1359(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1360(.a(gate173inter0), .b(s_116), .O(gate173inter1));
  and2  gate1361(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1362(.a(s_116), .O(gate173inter3));
  inv1  gate1363(.a(s_117), .O(gate173inter4));
  nand2 gate1364(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1365(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1366(.a(G486), .O(gate173inter7));
  inv1  gate1367(.a(G552), .O(gate173inter8));
  nand2 gate1368(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1369(.a(s_117), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1370(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1371(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1372(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1597(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1598(.a(gate175inter0), .b(s_150), .O(gate175inter1));
  and2  gate1599(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1600(.a(s_150), .O(gate175inter3));
  inv1  gate1601(.a(s_151), .O(gate175inter4));
  nand2 gate1602(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1603(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1604(.a(G492), .O(gate175inter7));
  inv1  gate1605(.a(G555), .O(gate175inter8));
  nand2 gate1606(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1607(.a(s_151), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1608(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1609(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1610(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1345(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1346(.a(gate186inter0), .b(s_114), .O(gate186inter1));
  and2  gate1347(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1348(.a(s_114), .O(gate186inter3));
  inv1  gate1349(.a(s_115), .O(gate186inter4));
  nand2 gate1350(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1351(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1352(.a(G572), .O(gate186inter7));
  inv1  gate1353(.a(G573), .O(gate186inter8));
  nand2 gate1354(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1355(.a(s_115), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1356(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1357(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1358(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1135(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1136(.a(gate189inter0), .b(s_84), .O(gate189inter1));
  and2  gate1137(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1138(.a(s_84), .O(gate189inter3));
  inv1  gate1139(.a(s_85), .O(gate189inter4));
  nand2 gate1140(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1141(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1142(.a(G578), .O(gate189inter7));
  inv1  gate1143(.a(G579), .O(gate189inter8));
  nand2 gate1144(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1145(.a(s_85), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1146(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1147(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1148(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate575(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate576(.a(gate190inter0), .b(s_4), .O(gate190inter1));
  and2  gate577(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate578(.a(s_4), .O(gate190inter3));
  inv1  gate579(.a(s_5), .O(gate190inter4));
  nand2 gate580(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate581(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate582(.a(G580), .O(gate190inter7));
  inv1  gate583(.a(G581), .O(gate190inter8));
  nand2 gate584(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate585(.a(s_5), .b(gate190inter3), .O(gate190inter10));
  nor2  gate586(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate587(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate588(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1709(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1710(.a(gate197inter0), .b(s_166), .O(gate197inter1));
  and2  gate1711(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1712(.a(s_166), .O(gate197inter3));
  inv1  gate1713(.a(s_167), .O(gate197inter4));
  nand2 gate1714(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1715(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1716(.a(G594), .O(gate197inter7));
  inv1  gate1717(.a(G595), .O(gate197inter8));
  nand2 gate1718(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1719(.a(s_167), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1720(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1721(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1722(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1961(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1962(.a(gate198inter0), .b(s_202), .O(gate198inter1));
  and2  gate1963(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1964(.a(s_202), .O(gate198inter3));
  inv1  gate1965(.a(s_203), .O(gate198inter4));
  nand2 gate1966(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1967(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1968(.a(G596), .O(gate198inter7));
  inv1  gate1969(.a(G597), .O(gate198inter8));
  nand2 gate1970(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1971(.a(s_203), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1972(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1973(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1974(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1835(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1836(.a(gate199inter0), .b(s_184), .O(gate199inter1));
  and2  gate1837(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1838(.a(s_184), .O(gate199inter3));
  inv1  gate1839(.a(s_185), .O(gate199inter4));
  nand2 gate1840(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1841(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1842(.a(G598), .O(gate199inter7));
  inv1  gate1843(.a(G599), .O(gate199inter8));
  nand2 gate1844(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1845(.a(s_185), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1846(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1847(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1848(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1289(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1290(.a(gate207inter0), .b(s_106), .O(gate207inter1));
  and2  gate1291(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1292(.a(s_106), .O(gate207inter3));
  inv1  gate1293(.a(s_107), .O(gate207inter4));
  nand2 gate1294(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1295(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1296(.a(G622), .O(gate207inter7));
  inv1  gate1297(.a(G632), .O(gate207inter8));
  nand2 gate1298(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1299(.a(s_107), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1300(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1301(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1302(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2003(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2004(.a(gate214inter0), .b(s_208), .O(gate214inter1));
  and2  gate2005(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2006(.a(s_208), .O(gate214inter3));
  inv1  gate2007(.a(s_209), .O(gate214inter4));
  nand2 gate2008(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2009(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2010(.a(G612), .O(gate214inter7));
  inv1  gate2011(.a(G672), .O(gate214inter8));
  nand2 gate2012(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2013(.a(s_209), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2014(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2015(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2016(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1485(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1486(.a(gate217inter0), .b(s_134), .O(gate217inter1));
  and2  gate1487(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1488(.a(s_134), .O(gate217inter3));
  inv1  gate1489(.a(s_135), .O(gate217inter4));
  nand2 gate1490(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1491(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1492(.a(G622), .O(gate217inter7));
  inv1  gate1493(.a(G678), .O(gate217inter8));
  nand2 gate1494(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1495(.a(s_135), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1496(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1497(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1498(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate687(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate688(.a(gate220inter0), .b(s_20), .O(gate220inter1));
  and2  gate689(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate690(.a(s_20), .O(gate220inter3));
  inv1  gate691(.a(s_21), .O(gate220inter4));
  nand2 gate692(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate693(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate694(.a(G637), .O(gate220inter7));
  inv1  gate695(.a(G681), .O(gate220inter8));
  nand2 gate696(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate697(.a(s_21), .b(gate220inter3), .O(gate220inter10));
  nor2  gate698(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate699(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate700(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1667(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1668(.a(gate221inter0), .b(s_160), .O(gate221inter1));
  and2  gate1669(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1670(.a(s_160), .O(gate221inter3));
  inv1  gate1671(.a(s_161), .O(gate221inter4));
  nand2 gate1672(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1673(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1674(.a(G622), .O(gate221inter7));
  inv1  gate1675(.a(G684), .O(gate221inter8));
  nand2 gate1676(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1677(.a(s_161), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1678(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1679(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1680(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate561(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate562(.a(gate227inter0), .b(s_2), .O(gate227inter1));
  and2  gate563(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate564(.a(s_2), .O(gate227inter3));
  inv1  gate565(.a(s_3), .O(gate227inter4));
  nand2 gate566(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate567(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate568(.a(G694), .O(gate227inter7));
  inv1  gate569(.a(G695), .O(gate227inter8));
  nand2 gate570(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate571(.a(s_3), .b(gate227inter3), .O(gate227inter10));
  nor2  gate572(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate573(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate574(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate2213(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2214(.a(gate228inter0), .b(s_238), .O(gate228inter1));
  and2  gate2215(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2216(.a(s_238), .O(gate228inter3));
  inv1  gate2217(.a(s_239), .O(gate228inter4));
  nand2 gate2218(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2219(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2220(.a(G696), .O(gate228inter7));
  inv1  gate2221(.a(G697), .O(gate228inter8));
  nand2 gate2222(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2223(.a(s_239), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2224(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2225(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2226(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate547(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate548(.a(gate229inter0), .b(s_0), .O(gate229inter1));
  and2  gate549(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate550(.a(s_0), .O(gate229inter3));
  inv1  gate551(.a(s_1), .O(gate229inter4));
  nand2 gate552(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate553(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate554(.a(G698), .O(gate229inter7));
  inv1  gate555(.a(G699), .O(gate229inter8));
  nand2 gate556(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate557(.a(s_1), .b(gate229inter3), .O(gate229inter10));
  nor2  gate558(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate559(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate560(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1401(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1402(.a(gate233inter0), .b(s_122), .O(gate233inter1));
  and2  gate1403(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1404(.a(s_122), .O(gate233inter3));
  inv1  gate1405(.a(s_123), .O(gate233inter4));
  nand2 gate1406(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1407(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1408(.a(G242), .O(gate233inter7));
  inv1  gate1409(.a(G718), .O(gate233inter8));
  nand2 gate1410(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1411(.a(s_123), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1412(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1413(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1414(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1541(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1542(.a(gate234inter0), .b(s_142), .O(gate234inter1));
  and2  gate1543(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1544(.a(s_142), .O(gate234inter3));
  inv1  gate1545(.a(s_143), .O(gate234inter4));
  nand2 gate1546(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1547(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1548(.a(G245), .O(gate234inter7));
  inv1  gate1549(.a(G721), .O(gate234inter8));
  nand2 gate1550(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1551(.a(s_143), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1552(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1553(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1554(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1751(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1752(.a(gate236inter0), .b(s_172), .O(gate236inter1));
  and2  gate1753(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1754(.a(s_172), .O(gate236inter3));
  inv1  gate1755(.a(s_173), .O(gate236inter4));
  nand2 gate1756(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1757(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1758(.a(G251), .O(gate236inter7));
  inv1  gate1759(.a(G727), .O(gate236inter8));
  nand2 gate1760(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1761(.a(s_173), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1762(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1763(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1764(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate869(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate870(.a(gate238inter0), .b(s_46), .O(gate238inter1));
  and2  gate871(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate872(.a(s_46), .O(gate238inter3));
  inv1  gate873(.a(s_47), .O(gate238inter4));
  nand2 gate874(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate875(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate876(.a(G257), .O(gate238inter7));
  inv1  gate877(.a(G709), .O(gate238inter8));
  nand2 gate878(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate879(.a(s_47), .b(gate238inter3), .O(gate238inter10));
  nor2  gate880(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate881(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate882(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1261(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1262(.a(gate239inter0), .b(s_102), .O(gate239inter1));
  and2  gate1263(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1264(.a(s_102), .O(gate239inter3));
  inv1  gate1265(.a(s_103), .O(gate239inter4));
  nand2 gate1266(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1267(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1268(.a(G260), .O(gate239inter7));
  inv1  gate1269(.a(G712), .O(gate239inter8));
  nand2 gate1270(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1271(.a(s_103), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1272(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1273(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1274(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1639(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1640(.a(gate266inter0), .b(s_156), .O(gate266inter1));
  and2  gate1641(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1642(.a(s_156), .O(gate266inter3));
  inv1  gate1643(.a(s_157), .O(gate266inter4));
  nand2 gate1644(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1645(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1646(.a(G645), .O(gate266inter7));
  inv1  gate1647(.a(G773), .O(gate266inter8));
  nand2 gate1648(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1649(.a(s_157), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1650(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1651(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1652(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1765(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1766(.a(gate269inter0), .b(s_174), .O(gate269inter1));
  and2  gate1767(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1768(.a(s_174), .O(gate269inter3));
  inv1  gate1769(.a(s_175), .O(gate269inter4));
  nand2 gate1770(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1771(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1772(.a(G654), .O(gate269inter7));
  inv1  gate1773(.a(G782), .O(gate269inter8));
  nand2 gate1774(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1775(.a(s_175), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1776(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1777(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1778(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate1849(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1850(.a(gate270inter0), .b(s_186), .O(gate270inter1));
  and2  gate1851(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1852(.a(s_186), .O(gate270inter3));
  inv1  gate1853(.a(s_187), .O(gate270inter4));
  nand2 gate1854(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1855(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1856(.a(G657), .O(gate270inter7));
  inv1  gate1857(.a(G785), .O(gate270inter8));
  nand2 gate1858(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1859(.a(s_187), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1860(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1861(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1862(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1891(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1892(.a(gate274inter0), .b(s_192), .O(gate274inter1));
  and2  gate1893(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1894(.a(s_192), .O(gate274inter3));
  inv1  gate1895(.a(s_193), .O(gate274inter4));
  nand2 gate1896(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1897(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1898(.a(G770), .O(gate274inter7));
  inv1  gate1899(.a(G794), .O(gate274inter8));
  nand2 gate1900(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1901(.a(s_193), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1902(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1903(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1904(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1611(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1612(.a(gate276inter0), .b(s_152), .O(gate276inter1));
  and2  gate1613(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1614(.a(s_152), .O(gate276inter3));
  inv1  gate1615(.a(s_153), .O(gate276inter4));
  nand2 gate1616(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1617(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1618(.a(G773), .O(gate276inter7));
  inv1  gate1619(.a(G797), .O(gate276inter8));
  nand2 gate1620(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1621(.a(s_153), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1622(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1623(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1624(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate589(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate590(.a(gate277inter0), .b(s_6), .O(gate277inter1));
  and2  gate591(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate592(.a(s_6), .O(gate277inter3));
  inv1  gate593(.a(s_7), .O(gate277inter4));
  nand2 gate594(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate595(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate596(.a(G648), .O(gate277inter7));
  inv1  gate597(.a(G800), .O(gate277inter8));
  nand2 gate598(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate599(.a(s_7), .b(gate277inter3), .O(gate277inter10));
  nor2  gate600(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate601(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate602(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1121(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1122(.a(gate278inter0), .b(s_82), .O(gate278inter1));
  and2  gate1123(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1124(.a(s_82), .O(gate278inter3));
  inv1  gate1125(.a(s_83), .O(gate278inter4));
  nand2 gate1126(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1127(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1128(.a(G776), .O(gate278inter7));
  inv1  gate1129(.a(G800), .O(gate278inter8));
  nand2 gate1130(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1131(.a(s_83), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1132(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1133(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1134(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2157(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2158(.a(gate280inter0), .b(s_230), .O(gate280inter1));
  and2  gate2159(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2160(.a(s_230), .O(gate280inter3));
  inv1  gate2161(.a(s_231), .O(gate280inter4));
  nand2 gate2162(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2163(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2164(.a(G779), .O(gate280inter7));
  inv1  gate2165(.a(G803), .O(gate280inter8));
  nand2 gate2166(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2167(.a(s_231), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2168(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2169(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2170(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1723(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1724(.a(gate284inter0), .b(s_168), .O(gate284inter1));
  and2  gate1725(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1726(.a(s_168), .O(gate284inter3));
  inv1  gate1727(.a(s_169), .O(gate284inter4));
  nand2 gate1728(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1729(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1730(.a(G785), .O(gate284inter7));
  inv1  gate1731(.a(G809), .O(gate284inter8));
  nand2 gate1732(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1733(.a(s_169), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1734(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1735(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1736(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1513(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1514(.a(gate286inter0), .b(s_138), .O(gate286inter1));
  and2  gate1515(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1516(.a(s_138), .O(gate286inter3));
  inv1  gate1517(.a(s_139), .O(gate286inter4));
  nand2 gate1518(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1519(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1520(.a(G788), .O(gate286inter7));
  inv1  gate1521(.a(G812), .O(gate286inter8));
  nand2 gate1522(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1523(.a(s_139), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1524(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1525(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1526(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1163(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1164(.a(gate287inter0), .b(s_88), .O(gate287inter1));
  and2  gate1165(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1166(.a(s_88), .O(gate287inter3));
  inv1  gate1167(.a(s_89), .O(gate287inter4));
  nand2 gate1168(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1169(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1170(.a(G663), .O(gate287inter7));
  inv1  gate1171(.a(G815), .O(gate287inter8));
  nand2 gate1172(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1173(.a(s_89), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1174(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1175(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1176(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate785(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate786(.a(gate288inter0), .b(s_34), .O(gate288inter1));
  and2  gate787(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate788(.a(s_34), .O(gate288inter3));
  inv1  gate789(.a(s_35), .O(gate288inter4));
  nand2 gate790(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate791(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate792(.a(G791), .O(gate288inter7));
  inv1  gate793(.a(G815), .O(gate288inter8));
  nand2 gate794(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate795(.a(s_35), .b(gate288inter3), .O(gate288inter10));
  nor2  gate796(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate797(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate798(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate939(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate940(.a(gate293inter0), .b(s_56), .O(gate293inter1));
  and2  gate941(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate942(.a(s_56), .O(gate293inter3));
  inv1  gate943(.a(s_57), .O(gate293inter4));
  nand2 gate944(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate945(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate946(.a(G828), .O(gate293inter7));
  inv1  gate947(.a(G829), .O(gate293inter8));
  nand2 gate948(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate949(.a(s_57), .b(gate293inter3), .O(gate293inter10));
  nor2  gate950(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate951(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate952(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate757(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate758(.a(gate295inter0), .b(s_30), .O(gate295inter1));
  and2  gate759(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate760(.a(s_30), .O(gate295inter3));
  inv1  gate761(.a(s_31), .O(gate295inter4));
  nand2 gate762(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate763(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate764(.a(G830), .O(gate295inter7));
  inv1  gate765(.a(G831), .O(gate295inter8));
  nand2 gate766(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate767(.a(s_31), .b(gate295inter3), .O(gate295inter10));
  nor2  gate768(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate769(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate770(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1681(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1682(.a(gate388inter0), .b(s_162), .O(gate388inter1));
  and2  gate1683(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1684(.a(s_162), .O(gate388inter3));
  inv1  gate1685(.a(s_163), .O(gate388inter4));
  nand2 gate1686(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1687(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1688(.a(G2), .O(gate388inter7));
  inv1  gate1689(.a(G1039), .O(gate388inter8));
  nand2 gate1690(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1691(.a(s_163), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1692(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1693(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1694(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1219(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1220(.a(gate390inter0), .b(s_96), .O(gate390inter1));
  and2  gate1221(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1222(.a(s_96), .O(gate390inter3));
  inv1  gate1223(.a(s_97), .O(gate390inter4));
  nand2 gate1224(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1225(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1226(.a(G4), .O(gate390inter7));
  inv1  gate1227(.a(G1045), .O(gate390inter8));
  nand2 gate1228(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1229(.a(s_97), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1230(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1231(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1232(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1093(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1094(.a(gate392inter0), .b(s_78), .O(gate392inter1));
  and2  gate1095(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1096(.a(s_78), .O(gate392inter3));
  inv1  gate1097(.a(s_79), .O(gate392inter4));
  nand2 gate1098(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1099(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1100(.a(G6), .O(gate392inter7));
  inv1  gate1101(.a(G1051), .O(gate392inter8));
  nand2 gate1102(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1103(.a(s_79), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1104(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1105(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1106(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1919(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1920(.a(gate395inter0), .b(s_196), .O(gate395inter1));
  and2  gate1921(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1922(.a(s_196), .O(gate395inter3));
  inv1  gate1923(.a(s_197), .O(gate395inter4));
  nand2 gate1924(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1925(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1926(.a(G9), .O(gate395inter7));
  inv1  gate1927(.a(G1060), .O(gate395inter8));
  nand2 gate1928(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1929(.a(s_197), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1930(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1931(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1932(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1583(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1584(.a(gate397inter0), .b(s_148), .O(gate397inter1));
  and2  gate1585(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1586(.a(s_148), .O(gate397inter3));
  inv1  gate1587(.a(s_149), .O(gate397inter4));
  nand2 gate1588(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1589(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1590(.a(G11), .O(gate397inter7));
  inv1  gate1591(.a(G1066), .O(gate397inter8));
  nand2 gate1592(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1593(.a(s_149), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1594(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1595(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1596(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1527(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1528(.a(gate401inter0), .b(s_140), .O(gate401inter1));
  and2  gate1529(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1530(.a(s_140), .O(gate401inter3));
  inv1  gate1531(.a(s_141), .O(gate401inter4));
  nand2 gate1532(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1533(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1534(.a(G15), .O(gate401inter7));
  inv1  gate1535(.a(G1078), .O(gate401inter8));
  nand2 gate1536(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1537(.a(s_141), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1538(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1539(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1540(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1457(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1458(.a(gate405inter0), .b(s_130), .O(gate405inter1));
  and2  gate1459(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1460(.a(s_130), .O(gate405inter3));
  inv1  gate1461(.a(s_131), .O(gate405inter4));
  nand2 gate1462(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1463(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1464(.a(G19), .O(gate405inter7));
  inv1  gate1465(.a(G1090), .O(gate405inter8));
  nand2 gate1466(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1467(.a(s_131), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1468(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1469(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1470(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1443(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1444(.a(gate407inter0), .b(s_128), .O(gate407inter1));
  and2  gate1445(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1446(.a(s_128), .O(gate407inter3));
  inv1  gate1447(.a(s_129), .O(gate407inter4));
  nand2 gate1448(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1449(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1450(.a(G21), .O(gate407inter7));
  inv1  gate1451(.a(G1096), .O(gate407inter8));
  nand2 gate1452(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1453(.a(s_129), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1454(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1455(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1456(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate995(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate996(.a(gate413inter0), .b(s_64), .O(gate413inter1));
  and2  gate997(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate998(.a(s_64), .O(gate413inter3));
  inv1  gate999(.a(s_65), .O(gate413inter4));
  nand2 gate1000(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1001(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1002(.a(G27), .O(gate413inter7));
  inv1  gate1003(.a(G1114), .O(gate413inter8));
  nand2 gate1004(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1005(.a(s_65), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1006(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1007(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1008(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate841(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate842(.a(gate414inter0), .b(s_42), .O(gate414inter1));
  and2  gate843(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate844(.a(s_42), .O(gate414inter3));
  inv1  gate845(.a(s_43), .O(gate414inter4));
  nand2 gate846(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate847(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate848(.a(G28), .O(gate414inter7));
  inv1  gate849(.a(G1117), .O(gate414inter8));
  nand2 gate850(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate851(.a(s_43), .b(gate414inter3), .O(gate414inter10));
  nor2  gate852(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate853(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate854(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1821(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1822(.a(gate417inter0), .b(s_182), .O(gate417inter1));
  and2  gate1823(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1824(.a(s_182), .O(gate417inter3));
  inv1  gate1825(.a(s_183), .O(gate417inter4));
  nand2 gate1826(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1827(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1828(.a(G31), .O(gate417inter7));
  inv1  gate1829(.a(G1126), .O(gate417inter8));
  nand2 gate1830(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1831(.a(s_183), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1832(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1833(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1834(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2199(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2200(.a(gate420inter0), .b(s_236), .O(gate420inter1));
  and2  gate2201(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2202(.a(s_236), .O(gate420inter3));
  inv1  gate2203(.a(s_237), .O(gate420inter4));
  nand2 gate2204(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2205(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2206(.a(G1036), .O(gate420inter7));
  inv1  gate2207(.a(G1132), .O(gate420inter8));
  nand2 gate2208(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2209(.a(s_237), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2210(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2211(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2212(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2059(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2060(.a(gate425inter0), .b(s_216), .O(gate425inter1));
  and2  gate2061(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2062(.a(s_216), .O(gate425inter3));
  inv1  gate2063(.a(s_217), .O(gate425inter4));
  nand2 gate2064(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2065(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2066(.a(G4), .O(gate425inter7));
  inv1  gate2067(.a(G1141), .O(gate425inter8));
  nand2 gate2068(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2069(.a(s_217), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2070(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2071(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2072(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate673(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate674(.a(gate436inter0), .b(s_18), .O(gate436inter1));
  and2  gate675(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate676(.a(s_18), .O(gate436inter3));
  inv1  gate677(.a(s_19), .O(gate436inter4));
  nand2 gate678(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate679(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate680(.a(G1060), .O(gate436inter7));
  inv1  gate681(.a(G1156), .O(gate436inter8));
  nand2 gate682(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate683(.a(s_19), .b(gate436inter3), .O(gate436inter10));
  nor2  gate684(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate685(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate686(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1331(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1332(.a(gate437inter0), .b(s_112), .O(gate437inter1));
  and2  gate1333(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1334(.a(s_112), .O(gate437inter3));
  inv1  gate1335(.a(s_113), .O(gate437inter4));
  nand2 gate1336(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1337(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1338(.a(G10), .O(gate437inter7));
  inv1  gate1339(.a(G1159), .O(gate437inter8));
  nand2 gate1340(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1341(.a(s_113), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1342(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1343(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1344(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1877(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1878(.a(gate443inter0), .b(s_190), .O(gate443inter1));
  and2  gate1879(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1880(.a(s_190), .O(gate443inter3));
  inv1  gate1881(.a(s_191), .O(gate443inter4));
  nand2 gate1882(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1883(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1884(.a(G13), .O(gate443inter7));
  inv1  gate1885(.a(G1168), .O(gate443inter8));
  nand2 gate1886(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1887(.a(s_191), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1888(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1889(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1890(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1947(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1948(.a(gate453inter0), .b(s_200), .O(gate453inter1));
  and2  gate1949(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1950(.a(s_200), .O(gate453inter3));
  inv1  gate1951(.a(s_201), .O(gate453inter4));
  nand2 gate1952(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1953(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1954(.a(G18), .O(gate453inter7));
  inv1  gate1955(.a(G1183), .O(gate453inter8));
  nand2 gate1956(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1957(.a(s_201), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1958(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1959(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1960(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate855(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate856(.a(gate459inter0), .b(s_44), .O(gate459inter1));
  and2  gate857(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate858(.a(s_44), .O(gate459inter3));
  inv1  gate859(.a(s_45), .O(gate459inter4));
  nand2 gate860(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate861(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate862(.a(G21), .O(gate459inter7));
  inv1  gate863(.a(G1192), .O(gate459inter8));
  nand2 gate864(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate865(.a(s_45), .b(gate459inter3), .O(gate459inter10));
  nor2  gate866(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate867(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate868(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate645(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate646(.a(gate460inter0), .b(s_14), .O(gate460inter1));
  and2  gate647(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate648(.a(s_14), .O(gate460inter3));
  inv1  gate649(.a(s_15), .O(gate460inter4));
  nand2 gate650(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate651(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate652(.a(G1096), .O(gate460inter7));
  inv1  gate653(.a(G1192), .O(gate460inter8));
  nand2 gate654(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate655(.a(s_15), .b(gate460inter3), .O(gate460inter10));
  nor2  gate656(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate657(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate658(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1065(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1066(.a(gate463inter0), .b(s_74), .O(gate463inter1));
  and2  gate1067(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1068(.a(s_74), .O(gate463inter3));
  inv1  gate1069(.a(s_75), .O(gate463inter4));
  nand2 gate1070(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1071(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1072(.a(G23), .O(gate463inter7));
  inv1  gate1073(.a(G1198), .O(gate463inter8));
  nand2 gate1074(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1075(.a(s_75), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1076(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1077(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1078(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2031(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2032(.a(gate465inter0), .b(s_212), .O(gate465inter1));
  and2  gate2033(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2034(.a(s_212), .O(gate465inter3));
  inv1  gate2035(.a(s_213), .O(gate465inter4));
  nand2 gate2036(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2037(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2038(.a(G24), .O(gate465inter7));
  inv1  gate2039(.a(G1201), .O(gate465inter8));
  nand2 gate2040(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2041(.a(s_213), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2042(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2043(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2044(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1625(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1626(.a(gate466inter0), .b(s_154), .O(gate466inter1));
  and2  gate1627(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1628(.a(s_154), .O(gate466inter3));
  inv1  gate1629(.a(s_155), .O(gate466inter4));
  nand2 gate1630(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1631(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1632(.a(G1105), .O(gate466inter7));
  inv1  gate1633(.a(G1201), .O(gate466inter8));
  nand2 gate1634(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1635(.a(s_155), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1636(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1637(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1638(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1863(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1864(.a(gate469inter0), .b(s_188), .O(gate469inter1));
  and2  gate1865(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1866(.a(s_188), .O(gate469inter3));
  inv1  gate1867(.a(s_189), .O(gate469inter4));
  nand2 gate1868(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1869(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1870(.a(G26), .O(gate469inter7));
  inv1  gate1871(.a(G1207), .O(gate469inter8));
  nand2 gate1872(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1873(.a(s_189), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1874(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1875(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1876(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2129(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2130(.a(gate471inter0), .b(s_226), .O(gate471inter1));
  and2  gate2131(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2132(.a(s_226), .O(gate471inter3));
  inv1  gate2133(.a(s_227), .O(gate471inter4));
  nand2 gate2134(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2135(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2136(.a(G27), .O(gate471inter7));
  inv1  gate2137(.a(G1210), .O(gate471inter8));
  nand2 gate2138(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2139(.a(s_227), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2140(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2141(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2142(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate743(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate744(.a(gate473inter0), .b(s_28), .O(gate473inter1));
  and2  gate745(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate746(.a(s_28), .O(gate473inter3));
  inv1  gate747(.a(s_29), .O(gate473inter4));
  nand2 gate748(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate749(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate750(.a(G28), .O(gate473inter7));
  inv1  gate751(.a(G1213), .O(gate473inter8));
  nand2 gate752(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate753(.a(s_29), .b(gate473inter3), .O(gate473inter10));
  nor2  gate754(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate755(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate756(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1793(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1794(.a(gate476inter0), .b(s_178), .O(gate476inter1));
  and2  gate1795(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1796(.a(s_178), .O(gate476inter3));
  inv1  gate1797(.a(s_179), .O(gate476inter4));
  nand2 gate1798(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1799(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1800(.a(G1120), .O(gate476inter7));
  inv1  gate1801(.a(G1216), .O(gate476inter8));
  nand2 gate1802(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1803(.a(s_179), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1804(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1805(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1806(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1373(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1374(.a(gate483inter0), .b(s_118), .O(gate483inter1));
  and2  gate1375(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1376(.a(s_118), .O(gate483inter3));
  inv1  gate1377(.a(s_119), .O(gate483inter4));
  nand2 gate1378(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1379(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1380(.a(G1228), .O(gate483inter7));
  inv1  gate1381(.a(G1229), .O(gate483inter8));
  nand2 gate1382(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1383(.a(s_119), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1384(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1385(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1386(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1499(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1500(.a(gate491inter0), .b(s_136), .O(gate491inter1));
  and2  gate1501(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1502(.a(s_136), .O(gate491inter3));
  inv1  gate1503(.a(s_137), .O(gate491inter4));
  nand2 gate1504(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1505(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1506(.a(G1244), .O(gate491inter7));
  inv1  gate1507(.a(G1245), .O(gate491inter8));
  nand2 gate1508(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1509(.a(s_137), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1510(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1511(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1512(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate771(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate772(.a(gate495inter0), .b(s_32), .O(gate495inter1));
  and2  gate773(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate774(.a(s_32), .O(gate495inter3));
  inv1  gate775(.a(s_33), .O(gate495inter4));
  nand2 gate776(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate777(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate778(.a(G1252), .O(gate495inter7));
  inv1  gate779(.a(G1253), .O(gate495inter8));
  nand2 gate780(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate781(.a(s_33), .b(gate495inter3), .O(gate495inter10));
  nor2  gate782(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate783(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate784(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1779(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1780(.a(gate499inter0), .b(s_176), .O(gate499inter1));
  and2  gate1781(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1782(.a(s_176), .O(gate499inter3));
  inv1  gate1783(.a(s_177), .O(gate499inter4));
  nand2 gate1784(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1785(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1786(.a(G1260), .O(gate499inter7));
  inv1  gate1787(.a(G1261), .O(gate499inter8));
  nand2 gate1788(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1789(.a(s_177), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1790(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1791(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1792(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1933(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1934(.a(gate500inter0), .b(s_198), .O(gate500inter1));
  and2  gate1935(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1936(.a(s_198), .O(gate500inter3));
  inv1  gate1937(.a(s_199), .O(gate500inter4));
  nand2 gate1938(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1939(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1940(.a(G1262), .O(gate500inter7));
  inv1  gate1941(.a(G1263), .O(gate500inter8));
  nand2 gate1942(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1943(.a(s_199), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1944(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1945(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1946(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1653(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1654(.a(gate501inter0), .b(s_158), .O(gate501inter1));
  and2  gate1655(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1656(.a(s_158), .O(gate501inter3));
  inv1  gate1657(.a(s_159), .O(gate501inter4));
  nand2 gate1658(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1659(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1660(.a(G1264), .O(gate501inter7));
  inv1  gate1661(.a(G1265), .O(gate501inter8));
  nand2 gate1662(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1663(.a(s_159), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1664(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1665(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1666(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate827(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate828(.a(gate502inter0), .b(s_40), .O(gate502inter1));
  and2  gate829(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate830(.a(s_40), .O(gate502inter3));
  inv1  gate831(.a(s_41), .O(gate502inter4));
  nand2 gate832(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate833(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate834(.a(G1266), .O(gate502inter7));
  inv1  gate835(.a(G1267), .O(gate502inter8));
  nand2 gate836(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate837(.a(s_41), .b(gate502inter3), .O(gate502inter10));
  nor2  gate838(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate839(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate840(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1303(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1304(.a(gate503inter0), .b(s_108), .O(gate503inter1));
  and2  gate1305(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1306(.a(s_108), .O(gate503inter3));
  inv1  gate1307(.a(s_109), .O(gate503inter4));
  nand2 gate1308(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1309(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1310(.a(G1268), .O(gate503inter7));
  inv1  gate1311(.a(G1269), .O(gate503inter8));
  nand2 gate1312(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1313(.a(s_109), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1314(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1315(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1316(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1415(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1416(.a(gate507inter0), .b(s_124), .O(gate507inter1));
  and2  gate1417(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1418(.a(s_124), .O(gate507inter3));
  inv1  gate1419(.a(s_125), .O(gate507inter4));
  nand2 gate1420(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1421(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1422(.a(G1276), .O(gate507inter7));
  inv1  gate1423(.a(G1277), .O(gate507inter8));
  nand2 gate1424(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1425(.a(s_125), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1426(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1427(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1428(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate659(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate660(.a(gate508inter0), .b(s_16), .O(gate508inter1));
  and2  gate661(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate662(.a(s_16), .O(gate508inter3));
  inv1  gate663(.a(s_17), .O(gate508inter4));
  nand2 gate664(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate665(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate666(.a(G1278), .O(gate508inter7));
  inv1  gate667(.a(G1279), .O(gate508inter8));
  nand2 gate668(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate669(.a(s_17), .b(gate508inter3), .O(gate508inter10));
  nor2  gate670(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate671(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate672(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate701(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate702(.a(gate509inter0), .b(s_22), .O(gate509inter1));
  and2  gate703(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate704(.a(s_22), .O(gate509inter3));
  inv1  gate705(.a(s_23), .O(gate509inter4));
  nand2 gate706(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate707(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate708(.a(G1280), .O(gate509inter7));
  inv1  gate709(.a(G1281), .O(gate509inter8));
  nand2 gate710(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate711(.a(s_23), .b(gate509inter3), .O(gate509inter10));
  nor2  gate712(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate713(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate714(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule