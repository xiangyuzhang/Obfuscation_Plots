module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );

  xor2  gate371(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate372(.a(gate20inter0), .b(s_30), .O(gate20inter1));
  and2  gate373(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate374(.a(s_30), .O(gate20inter3));
  inv1  gate375(.a(s_31), .O(gate20inter4));
  nand2 gate376(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate377(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate378(.a(N8), .O(gate20inter7));
  inv1  gate379(.a(N119), .O(gate20inter8));
  nand2 gate380(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate381(.a(s_31), .b(gate20inter3), .O(gate20inter10));
  nor2  gate382(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate383(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate384(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate231(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate232(.a(gate24inter0), .b(s_10), .O(gate24inter1));
  and2  gate233(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate234(.a(s_10), .O(gate24inter3));
  inv1  gate235(.a(s_11), .O(gate24inter4));
  nand2 gate236(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate237(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate238(.a(N130), .O(gate24inter7));
  inv1  gate239(.a(N43), .O(gate24inter8));
  nand2 gate240(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate241(.a(s_11), .b(gate24inter3), .O(gate24inter10));
  nor2  gate242(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate243(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate244(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate175(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate176(.a(gate27inter0), .b(s_2), .O(gate27inter1));
  and2  gate177(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate178(.a(s_2), .O(gate27inter3));
  inv1  gate179(.a(s_3), .O(gate27inter4));
  nand2 gate180(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate181(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate182(.a(N142), .O(gate27inter7));
  inv1  gate183(.a(N82), .O(gate27inter8));
  nand2 gate184(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate185(.a(s_3), .b(gate27inter3), .O(gate27inter10));
  nor2  gate186(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate187(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate188(.a(gate27inter12), .b(gate27inter1), .O(N174));

  xor2  gate273(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate274(.a(gate28inter0), .b(s_16), .O(gate28inter1));
  and2  gate275(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate276(.a(s_16), .O(gate28inter3));
  inv1  gate277(.a(s_17), .O(gate28inter4));
  nand2 gate278(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate279(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate280(.a(N146), .O(gate28inter7));
  inv1  gate281(.a(N95), .O(gate28inter8));
  nand2 gate282(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate283(.a(s_17), .b(gate28inter3), .O(gate28inter10));
  nor2  gate284(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate285(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate286(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );

  xor2  gate259(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate260(.a(gate35inter0), .b(s_14), .O(gate35inter1));
  and2  gate261(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate262(.a(s_14), .O(gate35inter3));
  inv1  gate263(.a(s_15), .O(gate35inter4));
  nand2 gate264(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate265(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate266(.a(N53), .O(gate35inter7));
  inv1  gate267(.a(N131), .O(gate35inter8));
  nand2 gate268(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate269(.a(s_15), .b(gate35inter3), .O(gate35inter10));
  nor2  gate270(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate271(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate272(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate203(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate204(.a(gate38inter0), .b(s_6), .O(gate38inter1));
  and2  gate205(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate206(.a(s_6), .O(gate38inter3));
  inv1  gate207(.a(s_7), .O(gate38inter4));
  nand2 gate208(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate209(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate210(.a(N73), .O(gate38inter7));
  inv1  gate211(.a(N139), .O(gate38inter8));
  nand2 gate212(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate213(.a(s_7), .b(gate38inter3), .O(gate38inter10));
  nor2  gate214(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate215(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate216(.a(gate38inter12), .b(gate38inter1), .O(N191));
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );

  xor2  gate315(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate316(.a(gate44inter0), .b(s_22), .O(gate44inter1));
  and2  gate317(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate318(.a(s_22), .O(gate44inter3));
  inv1  gate319(.a(s_23), .O(gate44inter4));
  nand2 gate320(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate321(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate322(.a(N112), .O(gate44inter7));
  inv1  gate323(.a(N151), .O(gate44inter8));
  nand2 gate324(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate325(.a(s_23), .b(gate44inter3), .O(gate44inter10));
  nor2  gate326(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate327(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate328(.a(gate44inter12), .b(gate44inter1), .O(N197));
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate161(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate162(.a(gate60inter0), .b(s_0), .O(gate60inter1));
  and2  gate163(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate164(.a(s_0), .O(gate60inter3));
  inv1  gate165(.a(s_1), .O(gate60inter4));
  nand2 gate166(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate167(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate168(.a(N213), .O(gate60inter7));
  inv1  gate169(.a(N24), .O(gate60inter8));
  nand2 gate170(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate171(.a(s_1), .b(gate60inter3), .O(gate60inter10));
  nor2  gate172(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate173(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate174(.a(gate60inter12), .b(gate60inter1), .O(N250));
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate301(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate302(.a(gate71inter0), .b(s_20), .O(gate71inter1));
  and2  gate303(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate304(.a(s_20), .O(gate71inter3));
  inv1  gate305(.a(s_21), .O(gate71inter4));
  nand2 gate306(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate307(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate308(.a(N230), .O(gate71inter7));
  inv1  gate309(.a(N185), .O(gate71inter8));
  nand2 gate310(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate311(.a(s_21), .b(gate71inter3), .O(gate71inter10));
  nor2  gate312(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate313(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate314(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );

  xor2  gate343(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate344(.a(gate84inter0), .b(s_26), .O(gate84inter1));
  and2  gate345(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate346(.a(s_26), .O(gate84inter3));
  inv1  gate347(.a(s_27), .O(gate84inter4));
  nand2 gate348(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate349(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate350(.a(N247), .O(gate84inter7));
  inv1  gate351(.a(N196), .O(gate84inter8));
  nand2 gate352(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate353(.a(s_27), .b(gate84inter3), .O(gate84inter10));
  nor2  gate354(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate355(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate356(.a(gate84inter12), .b(gate84inter1), .O(N294));
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate357(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate358(.a(gate105inter0), .b(s_28), .O(gate105inter1));
  and2  gate359(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate360(.a(s_28), .O(gate105inter3));
  inv1  gate361(.a(s_29), .O(gate105inter4));
  nand2 gate362(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate363(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate364(.a(N319), .O(gate105inter7));
  inv1  gate365(.a(N21), .O(gate105inter8));
  nand2 gate366(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate367(.a(s_29), .b(gate105inter3), .O(gate105inter10));
  nor2  gate368(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate369(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate370(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate287(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate288(.a(gate113inter0), .b(s_18), .O(gate113inter1));
  and2  gate289(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate290(.a(s_18), .O(gate113inter3));
  inv1  gate291(.a(s_19), .O(gate113inter4));
  nand2 gate292(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate293(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate294(.a(N319), .O(gate113inter7));
  inv1  gate295(.a(N73), .O(gate113inter8));
  nand2 gate296(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate297(.a(s_19), .b(gate113inter3), .O(gate113inter10));
  nor2  gate298(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate299(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate300(.a(gate113inter12), .b(gate113inter1), .O(N344));

  xor2  gate217(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate218(.a(gate114inter0), .b(s_8), .O(gate114inter1));
  and2  gate219(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate220(.a(s_8), .O(gate114inter3));
  inv1  gate221(.a(s_9), .O(gate114inter4));
  nand2 gate222(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate223(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate224(.a(N319), .O(gate114inter7));
  inv1  gate225(.a(N86), .O(gate114inter8));
  nand2 gate226(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate227(.a(s_9), .b(gate114inter3), .O(gate114inter10));
  nor2  gate228(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate229(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate230(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate245(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate246(.a(gate118inter0), .b(s_12), .O(gate118inter1));
  and2  gate247(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate248(.a(s_12), .O(gate118inter3));
  inv1  gate249(.a(s_13), .O(gate118inter4));
  nand2 gate250(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate251(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate252(.a(N331), .O(gate118inter7));
  inv1  gate253(.a(N301), .O(gate118inter8));
  nand2 gate254(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate255(.a(s_13), .b(gate118inter3), .O(gate118inter10));
  nor2  gate256(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate257(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate258(.a(gate118inter12), .b(gate118inter1), .O(N349));
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );

  xor2  gate329(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate330(.a(gate134inter0), .b(s_24), .O(gate134inter1));
  and2  gate331(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate332(.a(s_24), .O(gate134inter3));
  inv1  gate333(.a(s_25), .O(gate134inter4));
  nand2 gate334(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate335(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate336(.a(N360), .O(gate134inter7));
  inv1  gate337(.a(N79), .O(gate134inter8));
  nand2 gate338(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate339(.a(s_25), .b(gate134inter3), .O(gate134inter10));
  nor2  gate340(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate341(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate342(.a(gate134inter12), .b(gate134inter1), .O(N376));
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );

  xor2  gate189(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate190(.a(gate137inter0), .b(s_4), .O(gate137inter1));
  and2  gate191(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate192(.a(s_4), .O(gate137inter3));
  inv1  gate193(.a(s_5), .O(gate137inter4));
  nand2 gate194(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate195(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate196(.a(N360), .O(gate137inter7));
  inv1  gate197(.a(N115), .O(gate137inter8));
  nand2 gate198(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate199(.a(s_5), .b(gate137inter3), .O(gate137inter10));
  nor2  gate200(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate201(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate202(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule