module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate617(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate618(.a(gate9inter0), .b(s_10), .O(gate9inter1));
  and2  gate619(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate620(.a(s_10), .O(gate9inter3));
  inv1  gate621(.a(s_11), .O(gate9inter4));
  nand2 gate622(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate623(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate624(.a(G1), .O(gate9inter7));
  inv1  gate625(.a(G2), .O(gate9inter8));
  nand2 gate626(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate627(.a(s_11), .b(gate9inter3), .O(gate9inter10));
  nor2  gate628(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate629(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate630(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate561(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate562(.a(gate12inter0), .b(s_2), .O(gate12inter1));
  and2  gate563(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate564(.a(s_2), .O(gate12inter3));
  inv1  gate565(.a(s_3), .O(gate12inter4));
  nand2 gate566(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate567(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate568(.a(G7), .O(gate12inter7));
  inv1  gate569(.a(G8), .O(gate12inter8));
  nand2 gate570(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate571(.a(s_3), .b(gate12inter3), .O(gate12inter10));
  nor2  gate572(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate573(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate574(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1331(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1332(.a(gate15inter0), .b(s_112), .O(gate15inter1));
  and2  gate1333(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1334(.a(s_112), .O(gate15inter3));
  inv1  gate1335(.a(s_113), .O(gate15inter4));
  nand2 gate1336(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1337(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1338(.a(G13), .O(gate15inter7));
  inv1  gate1339(.a(G14), .O(gate15inter8));
  nand2 gate1340(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1341(.a(s_113), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1342(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1343(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1344(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate575(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate576(.a(gate22inter0), .b(s_4), .O(gate22inter1));
  and2  gate577(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate578(.a(s_4), .O(gate22inter3));
  inv1  gate579(.a(s_5), .O(gate22inter4));
  nand2 gate580(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate581(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate582(.a(G27), .O(gate22inter7));
  inv1  gate583(.a(G28), .O(gate22inter8));
  nand2 gate584(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate585(.a(s_5), .b(gate22inter3), .O(gate22inter10));
  nor2  gate586(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate587(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate588(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1023(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1024(.a(gate26inter0), .b(s_68), .O(gate26inter1));
  and2  gate1025(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1026(.a(s_68), .O(gate26inter3));
  inv1  gate1027(.a(s_69), .O(gate26inter4));
  nand2 gate1028(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1029(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1030(.a(G9), .O(gate26inter7));
  inv1  gate1031(.a(G13), .O(gate26inter8));
  nand2 gate1032(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1033(.a(s_69), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1034(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1035(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1036(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate1359(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1360(.a(gate27inter0), .b(s_116), .O(gate27inter1));
  and2  gate1361(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1362(.a(s_116), .O(gate27inter3));
  inv1  gate1363(.a(s_117), .O(gate27inter4));
  nand2 gate1364(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1365(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1366(.a(G2), .O(gate27inter7));
  inv1  gate1367(.a(G6), .O(gate27inter8));
  nand2 gate1368(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1369(.a(s_117), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1370(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1371(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1372(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1275(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1276(.a(gate36inter0), .b(s_104), .O(gate36inter1));
  and2  gate1277(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1278(.a(s_104), .O(gate36inter3));
  inv1  gate1279(.a(s_105), .O(gate36inter4));
  nand2 gate1280(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1281(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1282(.a(G26), .O(gate36inter7));
  inv1  gate1283(.a(G30), .O(gate36inter8));
  nand2 gate1284(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1285(.a(s_105), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1286(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1287(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1288(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate897(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate898(.a(gate46inter0), .b(s_50), .O(gate46inter1));
  and2  gate899(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate900(.a(s_50), .O(gate46inter3));
  inv1  gate901(.a(s_51), .O(gate46inter4));
  nand2 gate902(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate903(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate904(.a(G6), .O(gate46inter7));
  inv1  gate905(.a(G272), .O(gate46inter8));
  nand2 gate906(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate907(.a(s_51), .b(gate46inter3), .O(gate46inter10));
  nor2  gate908(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate909(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate910(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate743(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate744(.a(gate52inter0), .b(s_28), .O(gate52inter1));
  and2  gate745(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate746(.a(s_28), .O(gate52inter3));
  inv1  gate747(.a(s_29), .O(gate52inter4));
  nand2 gate748(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate749(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate750(.a(G12), .O(gate52inter7));
  inv1  gate751(.a(G281), .O(gate52inter8));
  nand2 gate752(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate753(.a(s_29), .b(gate52inter3), .O(gate52inter10));
  nor2  gate754(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate755(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate756(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate771(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate772(.a(gate53inter0), .b(s_32), .O(gate53inter1));
  and2  gate773(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate774(.a(s_32), .O(gate53inter3));
  inv1  gate775(.a(s_33), .O(gate53inter4));
  nand2 gate776(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate777(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate778(.a(G13), .O(gate53inter7));
  inv1  gate779(.a(G284), .O(gate53inter8));
  nand2 gate780(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate781(.a(s_33), .b(gate53inter3), .O(gate53inter10));
  nor2  gate782(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate783(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate784(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1163(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1164(.a(gate62inter0), .b(s_88), .O(gate62inter1));
  and2  gate1165(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1166(.a(s_88), .O(gate62inter3));
  inv1  gate1167(.a(s_89), .O(gate62inter4));
  nand2 gate1168(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1169(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1170(.a(G22), .O(gate62inter7));
  inv1  gate1171(.a(G296), .O(gate62inter8));
  nand2 gate1172(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1173(.a(s_89), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1174(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1175(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1176(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate785(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate786(.a(gate67inter0), .b(s_34), .O(gate67inter1));
  and2  gate787(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate788(.a(s_34), .O(gate67inter3));
  inv1  gate789(.a(s_35), .O(gate67inter4));
  nand2 gate790(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate791(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate792(.a(G27), .O(gate67inter7));
  inv1  gate793(.a(G305), .O(gate67inter8));
  nand2 gate794(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate795(.a(s_35), .b(gate67inter3), .O(gate67inter10));
  nor2  gate796(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate797(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate798(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate841(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate842(.a(gate75inter0), .b(s_42), .O(gate75inter1));
  and2  gate843(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate844(.a(s_42), .O(gate75inter3));
  inv1  gate845(.a(s_43), .O(gate75inter4));
  nand2 gate846(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate847(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate848(.a(G9), .O(gate75inter7));
  inv1  gate849(.a(G317), .O(gate75inter8));
  nand2 gate850(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate851(.a(s_43), .b(gate75inter3), .O(gate75inter10));
  nor2  gate852(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate853(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate854(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate855(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate856(.a(gate78inter0), .b(s_44), .O(gate78inter1));
  and2  gate857(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate858(.a(s_44), .O(gate78inter3));
  inv1  gate859(.a(s_45), .O(gate78inter4));
  nand2 gate860(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate861(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate862(.a(G6), .O(gate78inter7));
  inv1  gate863(.a(G320), .O(gate78inter8));
  nand2 gate864(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate865(.a(s_45), .b(gate78inter3), .O(gate78inter10));
  nor2  gate866(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate867(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate868(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate659(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate660(.a(gate80inter0), .b(s_16), .O(gate80inter1));
  and2  gate661(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate662(.a(s_16), .O(gate80inter3));
  inv1  gate663(.a(s_17), .O(gate80inter4));
  nand2 gate664(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate665(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate666(.a(G14), .O(gate80inter7));
  inv1  gate667(.a(G323), .O(gate80inter8));
  nand2 gate668(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate669(.a(s_17), .b(gate80inter3), .O(gate80inter10));
  nor2  gate670(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate671(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate672(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1149(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1150(.a(gate85inter0), .b(s_86), .O(gate85inter1));
  and2  gate1151(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1152(.a(s_86), .O(gate85inter3));
  inv1  gate1153(.a(s_87), .O(gate85inter4));
  nand2 gate1154(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1155(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1156(.a(G4), .O(gate85inter7));
  inv1  gate1157(.a(G332), .O(gate85inter8));
  nand2 gate1158(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1159(.a(s_87), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1160(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1161(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1162(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate701(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate702(.a(gate91inter0), .b(s_22), .O(gate91inter1));
  and2  gate703(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate704(.a(s_22), .O(gate91inter3));
  inv1  gate705(.a(s_23), .O(gate91inter4));
  nand2 gate706(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate707(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate708(.a(G25), .O(gate91inter7));
  inv1  gate709(.a(G341), .O(gate91inter8));
  nand2 gate710(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate711(.a(s_23), .b(gate91inter3), .O(gate91inter10));
  nor2  gate712(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate713(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate714(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1135(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1136(.a(gate111inter0), .b(s_84), .O(gate111inter1));
  and2  gate1137(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1138(.a(s_84), .O(gate111inter3));
  inv1  gate1139(.a(s_85), .O(gate111inter4));
  nand2 gate1140(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1141(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1142(.a(G374), .O(gate111inter7));
  inv1  gate1143(.a(G375), .O(gate111inter8));
  nand2 gate1144(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1145(.a(s_85), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1146(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1147(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1148(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1289(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1290(.a(gate114inter0), .b(s_106), .O(gate114inter1));
  and2  gate1291(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1292(.a(s_106), .O(gate114inter3));
  inv1  gate1293(.a(s_107), .O(gate114inter4));
  nand2 gate1294(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1295(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1296(.a(G380), .O(gate114inter7));
  inv1  gate1297(.a(G381), .O(gate114inter8));
  nand2 gate1298(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1299(.a(s_107), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1300(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1301(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1302(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1261(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1262(.a(gate117inter0), .b(s_102), .O(gate117inter1));
  and2  gate1263(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1264(.a(s_102), .O(gate117inter3));
  inv1  gate1265(.a(s_103), .O(gate117inter4));
  nand2 gate1266(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1267(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1268(.a(G386), .O(gate117inter7));
  inv1  gate1269(.a(G387), .O(gate117inter8));
  nand2 gate1270(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1271(.a(s_103), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1272(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1273(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1274(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate939(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate940(.a(gate126inter0), .b(s_56), .O(gate126inter1));
  and2  gate941(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate942(.a(s_56), .O(gate126inter3));
  inv1  gate943(.a(s_57), .O(gate126inter4));
  nand2 gate944(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate945(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate946(.a(G404), .O(gate126inter7));
  inv1  gate947(.a(G405), .O(gate126inter8));
  nand2 gate948(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate949(.a(s_57), .b(gate126inter3), .O(gate126inter10));
  nor2  gate950(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate951(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate952(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1093(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1094(.a(gate140inter0), .b(s_78), .O(gate140inter1));
  and2  gate1095(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1096(.a(s_78), .O(gate140inter3));
  inv1  gate1097(.a(s_79), .O(gate140inter4));
  nand2 gate1098(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1099(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1100(.a(G444), .O(gate140inter7));
  inv1  gate1101(.a(G447), .O(gate140inter8));
  nand2 gate1102(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1103(.a(s_79), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1104(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1105(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1106(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate827(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate828(.a(gate141inter0), .b(s_40), .O(gate141inter1));
  and2  gate829(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate830(.a(s_40), .O(gate141inter3));
  inv1  gate831(.a(s_41), .O(gate141inter4));
  nand2 gate832(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate833(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate834(.a(G450), .O(gate141inter7));
  inv1  gate835(.a(G453), .O(gate141inter8));
  nand2 gate836(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate837(.a(s_41), .b(gate141inter3), .O(gate141inter10));
  nor2  gate838(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate839(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate840(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1345(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1346(.a(gate157inter0), .b(s_114), .O(gate157inter1));
  and2  gate1347(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1348(.a(s_114), .O(gate157inter3));
  inv1  gate1349(.a(s_115), .O(gate157inter4));
  nand2 gate1350(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1351(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1352(.a(G438), .O(gate157inter7));
  inv1  gate1353(.a(G528), .O(gate157inter8));
  nand2 gate1354(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1355(.a(s_115), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1356(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1357(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1358(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate925(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate926(.a(gate204inter0), .b(s_54), .O(gate204inter1));
  and2  gate927(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate928(.a(s_54), .O(gate204inter3));
  inv1  gate929(.a(s_55), .O(gate204inter4));
  nand2 gate930(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate931(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate932(.a(G607), .O(gate204inter7));
  inv1  gate933(.a(G617), .O(gate204inter8));
  nand2 gate934(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate935(.a(s_55), .b(gate204inter3), .O(gate204inter10));
  nor2  gate936(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate937(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate938(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1107(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1108(.a(gate207inter0), .b(s_80), .O(gate207inter1));
  and2  gate1109(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1110(.a(s_80), .O(gate207inter3));
  inv1  gate1111(.a(s_81), .O(gate207inter4));
  nand2 gate1112(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1113(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1114(.a(G622), .O(gate207inter7));
  inv1  gate1115(.a(G632), .O(gate207inter8));
  nand2 gate1116(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1117(.a(s_81), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1118(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1119(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1120(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate631(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate632(.a(gate214inter0), .b(s_12), .O(gate214inter1));
  and2  gate633(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate634(.a(s_12), .O(gate214inter3));
  inv1  gate635(.a(s_13), .O(gate214inter4));
  nand2 gate636(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate637(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate638(.a(G612), .O(gate214inter7));
  inv1  gate639(.a(G672), .O(gate214inter8));
  nand2 gate640(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate641(.a(s_13), .b(gate214inter3), .O(gate214inter10));
  nor2  gate642(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate643(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate644(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1219(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1220(.a(gate225inter0), .b(s_96), .O(gate225inter1));
  and2  gate1221(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1222(.a(s_96), .O(gate225inter3));
  inv1  gate1223(.a(s_97), .O(gate225inter4));
  nand2 gate1224(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1225(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1226(.a(G690), .O(gate225inter7));
  inv1  gate1227(.a(G691), .O(gate225inter8));
  nand2 gate1228(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1229(.a(s_97), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1230(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1231(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1232(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1247(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1248(.a(gate229inter0), .b(s_100), .O(gate229inter1));
  and2  gate1249(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1250(.a(s_100), .O(gate229inter3));
  inv1  gate1251(.a(s_101), .O(gate229inter4));
  nand2 gate1252(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1253(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1254(.a(G698), .O(gate229inter7));
  inv1  gate1255(.a(G699), .O(gate229inter8));
  nand2 gate1256(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1257(.a(s_101), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1258(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1259(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1260(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate981(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate982(.a(gate235inter0), .b(s_62), .O(gate235inter1));
  and2  gate983(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate984(.a(s_62), .O(gate235inter3));
  inv1  gate985(.a(s_63), .O(gate235inter4));
  nand2 gate986(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate987(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate988(.a(G248), .O(gate235inter7));
  inv1  gate989(.a(G724), .O(gate235inter8));
  nand2 gate990(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate991(.a(s_63), .b(gate235inter3), .O(gate235inter10));
  nor2  gate992(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate993(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate994(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate967(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate968(.a(gate247inter0), .b(s_60), .O(gate247inter1));
  and2  gate969(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate970(.a(s_60), .O(gate247inter3));
  inv1  gate971(.a(s_61), .O(gate247inter4));
  nand2 gate972(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate973(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate974(.a(G251), .O(gate247inter7));
  inv1  gate975(.a(G739), .O(gate247inter8));
  nand2 gate976(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate977(.a(s_61), .b(gate247inter3), .O(gate247inter10));
  nor2  gate978(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate979(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate980(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate995(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate996(.a(gate248inter0), .b(s_64), .O(gate248inter1));
  and2  gate997(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate998(.a(s_64), .O(gate248inter3));
  inv1  gate999(.a(s_65), .O(gate248inter4));
  nand2 gate1000(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1001(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1002(.a(G727), .O(gate248inter7));
  inv1  gate1003(.a(G739), .O(gate248inter8));
  nand2 gate1004(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1005(.a(s_65), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1006(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1007(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1008(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1051(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1052(.a(gate253inter0), .b(s_72), .O(gate253inter1));
  and2  gate1053(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1054(.a(s_72), .O(gate253inter3));
  inv1  gate1055(.a(s_73), .O(gate253inter4));
  nand2 gate1056(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1057(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1058(.a(G260), .O(gate253inter7));
  inv1  gate1059(.a(G748), .O(gate253inter8));
  nand2 gate1060(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1061(.a(s_73), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1062(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1063(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1064(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate589(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate590(.a(gate260inter0), .b(s_6), .O(gate260inter1));
  and2  gate591(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate592(.a(s_6), .O(gate260inter3));
  inv1  gate593(.a(s_7), .O(gate260inter4));
  nand2 gate594(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate595(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate596(.a(G760), .O(gate260inter7));
  inv1  gate597(.a(G761), .O(gate260inter8));
  nand2 gate598(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate599(.a(s_7), .b(gate260inter3), .O(gate260inter10));
  nor2  gate600(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate601(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate602(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1233(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1234(.a(gate269inter0), .b(s_98), .O(gate269inter1));
  and2  gate1235(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1236(.a(s_98), .O(gate269inter3));
  inv1  gate1237(.a(s_99), .O(gate269inter4));
  nand2 gate1238(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1239(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1240(.a(G654), .O(gate269inter7));
  inv1  gate1241(.a(G782), .O(gate269inter8));
  nand2 gate1242(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1243(.a(s_99), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1244(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1245(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1246(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate715(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate716(.a(gate283inter0), .b(s_24), .O(gate283inter1));
  and2  gate717(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate718(.a(s_24), .O(gate283inter3));
  inv1  gate719(.a(s_25), .O(gate283inter4));
  nand2 gate720(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate721(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate722(.a(G657), .O(gate283inter7));
  inv1  gate723(.a(G809), .O(gate283inter8));
  nand2 gate724(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate725(.a(s_25), .b(gate283inter3), .O(gate283inter10));
  nor2  gate726(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate727(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate728(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1079(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1080(.a(gate284inter0), .b(s_76), .O(gate284inter1));
  and2  gate1081(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1082(.a(s_76), .O(gate284inter3));
  inv1  gate1083(.a(s_77), .O(gate284inter4));
  nand2 gate1084(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1085(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1086(.a(G785), .O(gate284inter7));
  inv1  gate1087(.a(G809), .O(gate284inter8));
  nand2 gate1088(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1089(.a(s_77), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1090(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1091(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1092(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1387(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1388(.a(gate288inter0), .b(s_120), .O(gate288inter1));
  and2  gate1389(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1390(.a(s_120), .O(gate288inter3));
  inv1  gate1391(.a(s_121), .O(gate288inter4));
  nand2 gate1392(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1393(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1394(.a(G791), .O(gate288inter7));
  inv1  gate1395(.a(G815), .O(gate288inter8));
  nand2 gate1396(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1397(.a(s_121), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1398(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1399(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1400(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1303(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1304(.a(gate291inter0), .b(s_108), .O(gate291inter1));
  and2  gate1305(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1306(.a(s_108), .O(gate291inter3));
  inv1  gate1307(.a(s_109), .O(gate291inter4));
  nand2 gate1308(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1309(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1310(.a(G822), .O(gate291inter7));
  inv1  gate1311(.a(G823), .O(gate291inter8));
  nand2 gate1312(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1313(.a(s_109), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1314(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1315(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1316(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate757(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate758(.a(gate293inter0), .b(s_30), .O(gate293inter1));
  and2  gate759(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate760(.a(s_30), .O(gate293inter3));
  inv1  gate761(.a(s_31), .O(gate293inter4));
  nand2 gate762(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate763(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate764(.a(G828), .O(gate293inter7));
  inv1  gate765(.a(G829), .O(gate293inter8));
  nand2 gate766(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate767(.a(s_31), .b(gate293inter3), .O(gate293inter10));
  nor2  gate768(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate769(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate770(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate813(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate814(.a(gate387inter0), .b(s_38), .O(gate387inter1));
  and2  gate815(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate816(.a(s_38), .O(gate387inter3));
  inv1  gate817(.a(s_39), .O(gate387inter4));
  nand2 gate818(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate819(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate820(.a(G1), .O(gate387inter7));
  inv1  gate821(.a(G1036), .O(gate387inter8));
  nand2 gate822(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate823(.a(s_39), .b(gate387inter3), .O(gate387inter10));
  nor2  gate824(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate825(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate826(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1121(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1122(.a(gate390inter0), .b(s_82), .O(gate390inter1));
  and2  gate1123(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1124(.a(s_82), .O(gate390inter3));
  inv1  gate1125(.a(s_83), .O(gate390inter4));
  nand2 gate1126(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1127(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1128(.a(G4), .O(gate390inter7));
  inv1  gate1129(.a(G1045), .O(gate390inter8));
  nand2 gate1130(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1131(.a(s_83), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1132(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1133(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1134(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1191(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1192(.a(gate395inter0), .b(s_92), .O(gate395inter1));
  and2  gate1193(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1194(.a(s_92), .O(gate395inter3));
  inv1  gate1195(.a(s_93), .O(gate395inter4));
  nand2 gate1196(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1197(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1198(.a(G9), .O(gate395inter7));
  inv1  gate1199(.a(G1060), .O(gate395inter8));
  nand2 gate1200(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1201(.a(s_93), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1202(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1203(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1204(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate883(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate884(.a(gate402inter0), .b(s_48), .O(gate402inter1));
  and2  gate885(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate886(.a(s_48), .O(gate402inter3));
  inv1  gate887(.a(s_49), .O(gate402inter4));
  nand2 gate888(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate889(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate890(.a(G16), .O(gate402inter7));
  inv1  gate891(.a(G1081), .O(gate402inter8));
  nand2 gate892(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate893(.a(s_49), .b(gate402inter3), .O(gate402inter10));
  nor2  gate894(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate895(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate896(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1065(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1066(.a(gate416inter0), .b(s_74), .O(gate416inter1));
  and2  gate1067(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1068(.a(s_74), .O(gate416inter3));
  inv1  gate1069(.a(s_75), .O(gate416inter4));
  nand2 gate1070(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1071(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1072(.a(G30), .O(gate416inter7));
  inv1  gate1073(.a(G1123), .O(gate416inter8));
  nand2 gate1074(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1075(.a(s_75), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1076(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1077(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1078(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1205(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1206(.a(gate418inter0), .b(s_94), .O(gate418inter1));
  and2  gate1207(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1208(.a(s_94), .O(gate418inter3));
  inv1  gate1209(.a(s_95), .O(gate418inter4));
  nand2 gate1210(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1211(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1212(.a(G32), .O(gate418inter7));
  inv1  gate1213(.a(G1129), .O(gate418inter8));
  nand2 gate1214(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1215(.a(s_95), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1216(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1217(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1218(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1009(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1010(.a(gate446inter0), .b(s_66), .O(gate446inter1));
  and2  gate1011(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1012(.a(s_66), .O(gate446inter3));
  inv1  gate1013(.a(s_67), .O(gate446inter4));
  nand2 gate1014(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1015(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1016(.a(G1075), .O(gate446inter7));
  inv1  gate1017(.a(G1171), .O(gate446inter8));
  nand2 gate1018(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1019(.a(s_67), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1020(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1021(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1022(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1037(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1038(.a(gate460inter0), .b(s_70), .O(gate460inter1));
  and2  gate1039(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1040(.a(s_70), .O(gate460inter3));
  inv1  gate1041(.a(s_71), .O(gate460inter4));
  nand2 gate1042(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1043(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1044(.a(G1096), .O(gate460inter7));
  inv1  gate1045(.a(G1192), .O(gate460inter8));
  nand2 gate1046(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1047(.a(s_71), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1048(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1049(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1050(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate603(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate604(.a(gate475inter0), .b(s_8), .O(gate475inter1));
  and2  gate605(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate606(.a(s_8), .O(gate475inter3));
  inv1  gate607(.a(s_9), .O(gate475inter4));
  nand2 gate608(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate609(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate610(.a(G29), .O(gate475inter7));
  inv1  gate611(.a(G1216), .O(gate475inter8));
  nand2 gate612(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate613(.a(s_9), .b(gate475inter3), .O(gate475inter10));
  nor2  gate614(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate615(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate616(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate645(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate646(.a(gate476inter0), .b(s_14), .O(gate476inter1));
  and2  gate647(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate648(.a(s_14), .O(gate476inter3));
  inv1  gate649(.a(s_15), .O(gate476inter4));
  nand2 gate650(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate651(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate652(.a(G1120), .O(gate476inter7));
  inv1  gate653(.a(G1216), .O(gate476inter8));
  nand2 gate654(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate655(.a(s_15), .b(gate476inter3), .O(gate476inter10));
  nor2  gate656(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate657(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate658(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1373(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1374(.a(gate477inter0), .b(s_118), .O(gate477inter1));
  and2  gate1375(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1376(.a(s_118), .O(gate477inter3));
  inv1  gate1377(.a(s_119), .O(gate477inter4));
  nand2 gate1378(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1379(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1380(.a(G30), .O(gate477inter7));
  inv1  gate1381(.a(G1219), .O(gate477inter8));
  nand2 gate1382(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1383(.a(s_119), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1384(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1385(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1386(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate869(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate870(.a(gate478inter0), .b(s_46), .O(gate478inter1));
  and2  gate871(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate872(.a(s_46), .O(gate478inter3));
  inv1  gate873(.a(s_47), .O(gate478inter4));
  nand2 gate874(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate875(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate876(.a(G1123), .O(gate478inter7));
  inv1  gate877(.a(G1219), .O(gate478inter8));
  nand2 gate878(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate879(.a(s_47), .b(gate478inter3), .O(gate478inter10));
  nor2  gate880(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate881(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate882(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate799(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate800(.a(gate479inter0), .b(s_36), .O(gate479inter1));
  and2  gate801(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate802(.a(s_36), .O(gate479inter3));
  inv1  gate803(.a(s_37), .O(gate479inter4));
  nand2 gate804(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate805(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate806(.a(G31), .O(gate479inter7));
  inv1  gate807(.a(G1222), .O(gate479inter8));
  nand2 gate808(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate809(.a(s_37), .b(gate479inter3), .O(gate479inter10));
  nor2  gate810(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate811(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate812(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate953(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate954(.a(gate482inter0), .b(s_58), .O(gate482inter1));
  and2  gate955(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate956(.a(s_58), .O(gate482inter3));
  inv1  gate957(.a(s_59), .O(gate482inter4));
  nand2 gate958(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate959(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate960(.a(G1129), .O(gate482inter7));
  inv1  gate961(.a(G1225), .O(gate482inter8));
  nand2 gate962(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate963(.a(s_59), .b(gate482inter3), .O(gate482inter10));
  nor2  gate964(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate965(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate966(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1177(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1178(.a(gate488inter0), .b(s_90), .O(gate488inter1));
  and2  gate1179(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1180(.a(s_90), .O(gate488inter3));
  inv1  gate1181(.a(s_91), .O(gate488inter4));
  nand2 gate1182(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1183(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1184(.a(G1238), .O(gate488inter7));
  inv1  gate1185(.a(G1239), .O(gate488inter8));
  nand2 gate1186(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1187(.a(s_91), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1188(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1189(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1190(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1317(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1318(.a(gate493inter0), .b(s_110), .O(gate493inter1));
  and2  gate1319(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1320(.a(s_110), .O(gate493inter3));
  inv1  gate1321(.a(s_111), .O(gate493inter4));
  nand2 gate1322(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1323(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1324(.a(G1248), .O(gate493inter7));
  inv1  gate1325(.a(G1249), .O(gate493inter8));
  nand2 gate1326(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1327(.a(s_111), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1328(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1329(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1330(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate687(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate688(.a(gate495inter0), .b(s_20), .O(gate495inter1));
  and2  gate689(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate690(.a(s_20), .O(gate495inter3));
  inv1  gate691(.a(s_21), .O(gate495inter4));
  nand2 gate692(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate693(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate694(.a(G1252), .O(gate495inter7));
  inv1  gate695(.a(G1253), .O(gate495inter8));
  nand2 gate696(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate697(.a(s_21), .b(gate495inter3), .O(gate495inter10));
  nor2  gate698(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate699(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate700(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate911(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate912(.a(gate496inter0), .b(s_52), .O(gate496inter1));
  and2  gate913(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate914(.a(s_52), .O(gate496inter3));
  inv1  gate915(.a(s_53), .O(gate496inter4));
  nand2 gate916(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate917(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate918(.a(G1254), .O(gate496inter7));
  inv1  gate919(.a(G1255), .O(gate496inter8));
  nand2 gate920(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate921(.a(s_53), .b(gate496inter3), .O(gate496inter10));
  nor2  gate922(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate923(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate924(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate673(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate674(.a(gate507inter0), .b(s_18), .O(gate507inter1));
  and2  gate675(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate676(.a(s_18), .O(gate507inter3));
  inv1  gate677(.a(s_19), .O(gate507inter4));
  nand2 gate678(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate679(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate680(.a(G1276), .O(gate507inter7));
  inv1  gate681(.a(G1277), .O(gate507inter8));
  nand2 gate682(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate683(.a(s_19), .b(gate507inter3), .O(gate507inter10));
  nor2  gate684(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate685(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate686(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate547(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate548(.a(gate511inter0), .b(s_0), .O(gate511inter1));
  and2  gate549(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate550(.a(s_0), .O(gate511inter3));
  inv1  gate551(.a(s_1), .O(gate511inter4));
  nand2 gate552(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate553(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate554(.a(G1284), .O(gate511inter7));
  inv1  gate555(.a(G1285), .O(gate511inter8));
  nand2 gate556(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate557(.a(s_1), .b(gate511inter3), .O(gate511inter10));
  nor2  gate558(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate559(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate560(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate729(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate730(.a(gate514inter0), .b(s_26), .O(gate514inter1));
  and2  gate731(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate732(.a(s_26), .O(gate514inter3));
  inv1  gate733(.a(s_27), .O(gate514inter4));
  nand2 gate734(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate735(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate736(.a(G1290), .O(gate514inter7));
  inv1  gate737(.a(G1291), .O(gate514inter8));
  nand2 gate738(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate739(.a(s_27), .b(gate514inter3), .O(gate514inter10));
  nor2  gate740(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate741(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate742(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule