module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate967(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate968(.a(gate10inter0), .b(s_60), .O(gate10inter1));
  and2  gate969(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate970(.a(s_60), .O(gate10inter3));
  inv1  gate971(.a(s_61), .O(gate10inter4));
  nand2 gate972(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate973(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate974(.a(G3), .O(gate10inter7));
  inv1  gate975(.a(G4), .O(gate10inter8));
  nand2 gate976(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate977(.a(s_61), .b(gate10inter3), .O(gate10inter10));
  nor2  gate978(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate979(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate980(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate995(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate996(.a(gate19inter0), .b(s_64), .O(gate19inter1));
  and2  gate997(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate998(.a(s_64), .O(gate19inter3));
  inv1  gate999(.a(s_65), .O(gate19inter4));
  nand2 gate1000(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1001(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1002(.a(G21), .O(gate19inter7));
  inv1  gate1003(.a(G22), .O(gate19inter8));
  nand2 gate1004(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1005(.a(s_65), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1006(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1007(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1008(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1443(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1444(.a(gate22inter0), .b(s_128), .O(gate22inter1));
  and2  gate1445(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1446(.a(s_128), .O(gate22inter3));
  inv1  gate1447(.a(s_129), .O(gate22inter4));
  nand2 gate1448(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1449(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1450(.a(G27), .O(gate22inter7));
  inv1  gate1451(.a(G28), .O(gate22inter8));
  nand2 gate1452(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1453(.a(s_129), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1454(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1455(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1456(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1415(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1416(.a(gate30inter0), .b(s_124), .O(gate30inter1));
  and2  gate1417(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1418(.a(s_124), .O(gate30inter3));
  inv1  gate1419(.a(s_125), .O(gate30inter4));
  nand2 gate1420(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1421(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1422(.a(G11), .O(gate30inter7));
  inv1  gate1423(.a(G15), .O(gate30inter8));
  nand2 gate1424(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1425(.a(s_125), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1426(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1427(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1428(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate841(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate842(.a(gate33inter0), .b(s_42), .O(gate33inter1));
  and2  gate843(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate844(.a(s_42), .O(gate33inter3));
  inv1  gate845(.a(s_43), .O(gate33inter4));
  nand2 gate846(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate847(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate848(.a(G17), .O(gate33inter7));
  inv1  gate849(.a(G21), .O(gate33inter8));
  nand2 gate850(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate851(.a(s_43), .b(gate33inter3), .O(gate33inter10));
  nor2  gate852(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate853(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate854(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1527(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1528(.a(gate34inter0), .b(s_140), .O(gate34inter1));
  and2  gate1529(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1530(.a(s_140), .O(gate34inter3));
  inv1  gate1531(.a(s_141), .O(gate34inter4));
  nand2 gate1532(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1533(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1534(.a(G25), .O(gate34inter7));
  inv1  gate1535(.a(G29), .O(gate34inter8));
  nand2 gate1536(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1537(.a(s_141), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1538(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1539(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1540(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate981(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate982(.a(gate39inter0), .b(s_62), .O(gate39inter1));
  and2  gate983(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate984(.a(s_62), .O(gate39inter3));
  inv1  gate985(.a(s_63), .O(gate39inter4));
  nand2 gate986(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate987(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate988(.a(G20), .O(gate39inter7));
  inv1  gate989(.a(G24), .O(gate39inter8));
  nand2 gate990(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate991(.a(s_63), .b(gate39inter3), .O(gate39inter10));
  nor2  gate992(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate993(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate994(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1639(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1640(.a(gate40inter0), .b(s_156), .O(gate40inter1));
  and2  gate1641(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1642(.a(s_156), .O(gate40inter3));
  inv1  gate1643(.a(s_157), .O(gate40inter4));
  nand2 gate1644(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1645(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1646(.a(G28), .O(gate40inter7));
  inv1  gate1647(.a(G32), .O(gate40inter8));
  nand2 gate1648(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1649(.a(s_157), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1650(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1651(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1652(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate827(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate828(.a(gate42inter0), .b(s_40), .O(gate42inter1));
  and2  gate829(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate830(.a(s_40), .O(gate42inter3));
  inv1  gate831(.a(s_41), .O(gate42inter4));
  nand2 gate832(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate833(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate834(.a(G2), .O(gate42inter7));
  inv1  gate835(.a(G266), .O(gate42inter8));
  nand2 gate836(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate837(.a(s_41), .b(gate42inter3), .O(gate42inter10));
  nor2  gate838(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate839(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate840(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1023(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1024(.a(gate43inter0), .b(s_68), .O(gate43inter1));
  and2  gate1025(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1026(.a(s_68), .O(gate43inter3));
  inv1  gate1027(.a(s_69), .O(gate43inter4));
  nand2 gate1028(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1029(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1030(.a(G3), .O(gate43inter7));
  inv1  gate1031(.a(G269), .O(gate43inter8));
  nand2 gate1032(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1033(.a(s_69), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1034(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1035(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1036(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1177(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1178(.a(gate52inter0), .b(s_90), .O(gate52inter1));
  and2  gate1179(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1180(.a(s_90), .O(gate52inter3));
  inv1  gate1181(.a(s_91), .O(gate52inter4));
  nand2 gate1182(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1183(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1184(.a(G12), .O(gate52inter7));
  inv1  gate1185(.a(G281), .O(gate52inter8));
  nand2 gate1186(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1187(.a(s_91), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1188(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1189(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1190(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1219(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1220(.a(gate53inter0), .b(s_96), .O(gate53inter1));
  and2  gate1221(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1222(.a(s_96), .O(gate53inter3));
  inv1  gate1223(.a(s_97), .O(gate53inter4));
  nand2 gate1224(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1225(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1226(.a(G13), .O(gate53inter7));
  inv1  gate1227(.a(G284), .O(gate53inter8));
  nand2 gate1228(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1229(.a(s_97), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1230(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1231(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1232(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1765(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1766(.a(gate59inter0), .b(s_174), .O(gate59inter1));
  and2  gate1767(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1768(.a(s_174), .O(gate59inter3));
  inv1  gate1769(.a(s_175), .O(gate59inter4));
  nand2 gate1770(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1771(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1772(.a(G19), .O(gate59inter7));
  inv1  gate1773(.a(G293), .O(gate59inter8));
  nand2 gate1774(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1775(.a(s_175), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1776(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1777(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1778(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate673(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate674(.a(gate60inter0), .b(s_18), .O(gate60inter1));
  and2  gate675(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate676(.a(s_18), .O(gate60inter3));
  inv1  gate677(.a(s_19), .O(gate60inter4));
  nand2 gate678(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate679(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate680(.a(G20), .O(gate60inter7));
  inv1  gate681(.a(G293), .O(gate60inter8));
  nand2 gate682(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate683(.a(s_19), .b(gate60inter3), .O(gate60inter10));
  nor2  gate684(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate685(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate686(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1331(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1332(.a(gate62inter0), .b(s_112), .O(gate62inter1));
  and2  gate1333(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1334(.a(s_112), .O(gate62inter3));
  inv1  gate1335(.a(s_113), .O(gate62inter4));
  nand2 gate1336(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1337(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1338(.a(G22), .O(gate62inter7));
  inv1  gate1339(.a(G296), .O(gate62inter8));
  nand2 gate1340(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1341(.a(s_113), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1342(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1343(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1344(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate869(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate870(.a(gate64inter0), .b(s_46), .O(gate64inter1));
  and2  gate871(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate872(.a(s_46), .O(gate64inter3));
  inv1  gate873(.a(s_47), .O(gate64inter4));
  nand2 gate874(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate875(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate876(.a(G24), .O(gate64inter7));
  inv1  gate877(.a(G299), .O(gate64inter8));
  nand2 gate878(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate879(.a(s_47), .b(gate64inter3), .O(gate64inter10));
  nor2  gate880(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate881(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate882(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate855(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate856(.a(gate67inter0), .b(s_44), .O(gate67inter1));
  and2  gate857(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate858(.a(s_44), .O(gate67inter3));
  inv1  gate859(.a(s_45), .O(gate67inter4));
  nand2 gate860(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate861(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate862(.a(G27), .O(gate67inter7));
  inv1  gate863(.a(G305), .O(gate67inter8));
  nand2 gate864(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate865(.a(s_45), .b(gate67inter3), .O(gate67inter10));
  nor2  gate866(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate867(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate868(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1695(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1696(.a(gate71inter0), .b(s_164), .O(gate71inter1));
  and2  gate1697(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1698(.a(s_164), .O(gate71inter3));
  inv1  gate1699(.a(s_165), .O(gate71inter4));
  nand2 gate1700(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1701(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1702(.a(G31), .O(gate71inter7));
  inv1  gate1703(.a(G311), .O(gate71inter8));
  nand2 gate1704(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1705(.a(s_165), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1706(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1707(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1708(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1863(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1864(.a(gate72inter0), .b(s_188), .O(gate72inter1));
  and2  gate1865(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1866(.a(s_188), .O(gate72inter3));
  inv1  gate1867(.a(s_189), .O(gate72inter4));
  nand2 gate1868(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1869(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1870(.a(G32), .O(gate72inter7));
  inv1  gate1871(.a(G311), .O(gate72inter8));
  nand2 gate1872(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1873(.a(s_189), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1874(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1875(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1876(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate799(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate800(.a(gate75inter0), .b(s_36), .O(gate75inter1));
  and2  gate801(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate802(.a(s_36), .O(gate75inter3));
  inv1  gate803(.a(s_37), .O(gate75inter4));
  nand2 gate804(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate805(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate806(.a(G9), .O(gate75inter7));
  inv1  gate807(.a(G317), .O(gate75inter8));
  nand2 gate808(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate809(.a(s_37), .b(gate75inter3), .O(gate75inter10));
  nor2  gate810(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate811(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate812(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1345(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1346(.a(gate78inter0), .b(s_114), .O(gate78inter1));
  and2  gate1347(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1348(.a(s_114), .O(gate78inter3));
  inv1  gate1349(.a(s_115), .O(gate78inter4));
  nand2 gate1350(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1351(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1352(.a(G6), .O(gate78inter7));
  inv1  gate1353(.a(G320), .O(gate78inter8));
  nand2 gate1354(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1355(.a(s_115), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1356(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1357(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1358(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate575(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate576(.a(gate82inter0), .b(s_4), .O(gate82inter1));
  and2  gate577(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate578(.a(s_4), .O(gate82inter3));
  inv1  gate579(.a(s_5), .O(gate82inter4));
  nand2 gate580(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate581(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate582(.a(G7), .O(gate82inter7));
  inv1  gate583(.a(G326), .O(gate82inter8));
  nand2 gate584(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate585(.a(s_5), .b(gate82inter3), .O(gate82inter10));
  nor2  gate586(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate587(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate588(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate785(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate786(.a(gate91inter0), .b(s_34), .O(gate91inter1));
  and2  gate787(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate788(.a(s_34), .O(gate91inter3));
  inv1  gate789(.a(s_35), .O(gate91inter4));
  nand2 gate790(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate791(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate792(.a(G25), .O(gate91inter7));
  inv1  gate793(.a(G341), .O(gate91inter8));
  nand2 gate794(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate795(.a(s_35), .b(gate91inter3), .O(gate91inter10));
  nor2  gate796(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate797(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate798(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1583(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1584(.a(gate95inter0), .b(s_148), .O(gate95inter1));
  and2  gate1585(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1586(.a(s_148), .O(gate95inter3));
  inv1  gate1587(.a(s_149), .O(gate95inter4));
  nand2 gate1588(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1589(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1590(.a(G26), .O(gate95inter7));
  inv1  gate1591(.a(G347), .O(gate95inter8));
  nand2 gate1592(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1593(.a(s_149), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1594(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1595(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1596(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1359(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1360(.a(gate97inter0), .b(s_116), .O(gate97inter1));
  and2  gate1361(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1362(.a(s_116), .O(gate97inter3));
  inv1  gate1363(.a(s_117), .O(gate97inter4));
  nand2 gate1364(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1365(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1366(.a(G19), .O(gate97inter7));
  inv1  gate1367(.a(G350), .O(gate97inter8));
  nand2 gate1368(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1369(.a(s_117), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1370(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1371(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1372(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1401(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1402(.a(gate103inter0), .b(s_122), .O(gate103inter1));
  and2  gate1403(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1404(.a(s_122), .O(gate103inter3));
  inv1  gate1405(.a(s_123), .O(gate103inter4));
  nand2 gate1406(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1407(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1408(.a(G28), .O(gate103inter7));
  inv1  gate1409(.a(G359), .O(gate103inter8));
  nand2 gate1410(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1411(.a(s_123), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1412(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1413(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1414(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1919(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1920(.a(gate104inter0), .b(s_196), .O(gate104inter1));
  and2  gate1921(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1922(.a(s_196), .O(gate104inter3));
  inv1  gate1923(.a(s_197), .O(gate104inter4));
  nand2 gate1924(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1925(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1926(.a(G32), .O(gate104inter7));
  inv1  gate1927(.a(G359), .O(gate104inter8));
  nand2 gate1928(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1929(.a(s_197), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1930(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1931(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1932(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1093(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1094(.a(gate116inter0), .b(s_78), .O(gate116inter1));
  and2  gate1095(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1096(.a(s_78), .O(gate116inter3));
  inv1  gate1097(.a(s_79), .O(gate116inter4));
  nand2 gate1098(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1099(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1100(.a(G384), .O(gate116inter7));
  inv1  gate1101(.a(G385), .O(gate116inter8));
  nand2 gate1102(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1103(.a(s_79), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1104(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1105(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1106(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1877(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1878(.a(gate118inter0), .b(s_190), .O(gate118inter1));
  and2  gate1879(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1880(.a(s_190), .O(gate118inter3));
  inv1  gate1881(.a(s_191), .O(gate118inter4));
  nand2 gate1882(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1883(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1884(.a(G388), .O(gate118inter7));
  inv1  gate1885(.a(G389), .O(gate118inter8));
  nand2 gate1886(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1887(.a(s_191), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1888(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1889(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1890(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1541(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1542(.a(gate124inter0), .b(s_142), .O(gate124inter1));
  and2  gate1543(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1544(.a(s_142), .O(gate124inter3));
  inv1  gate1545(.a(s_143), .O(gate124inter4));
  nand2 gate1546(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1547(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1548(.a(G400), .O(gate124inter7));
  inv1  gate1549(.a(G401), .O(gate124inter8));
  nand2 gate1550(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1551(.a(s_143), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1552(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1553(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1554(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1807(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1808(.a(gate128inter0), .b(s_180), .O(gate128inter1));
  and2  gate1809(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1810(.a(s_180), .O(gate128inter3));
  inv1  gate1811(.a(s_181), .O(gate128inter4));
  nand2 gate1812(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1813(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1814(.a(G408), .O(gate128inter7));
  inv1  gate1815(.a(G409), .O(gate128inter8));
  nand2 gate1816(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1817(.a(s_181), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1818(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1819(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1820(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1611(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1612(.a(gate130inter0), .b(s_152), .O(gate130inter1));
  and2  gate1613(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1614(.a(s_152), .O(gate130inter3));
  inv1  gate1615(.a(s_153), .O(gate130inter4));
  nand2 gate1616(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1617(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1618(.a(G412), .O(gate130inter7));
  inv1  gate1619(.a(G413), .O(gate130inter8));
  nand2 gate1620(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1621(.a(s_153), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1622(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1623(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1624(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1499(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1500(.a(gate135inter0), .b(s_136), .O(gate135inter1));
  and2  gate1501(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1502(.a(s_136), .O(gate135inter3));
  inv1  gate1503(.a(s_137), .O(gate135inter4));
  nand2 gate1504(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1505(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1506(.a(G422), .O(gate135inter7));
  inv1  gate1507(.a(G423), .O(gate135inter8));
  nand2 gate1508(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1509(.a(s_137), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1510(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1511(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1512(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1261(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1262(.a(gate142inter0), .b(s_102), .O(gate142inter1));
  and2  gate1263(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1264(.a(s_102), .O(gate142inter3));
  inv1  gate1265(.a(s_103), .O(gate142inter4));
  nand2 gate1266(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1267(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1268(.a(G456), .O(gate142inter7));
  inv1  gate1269(.a(G459), .O(gate142inter8));
  nand2 gate1270(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1271(.a(s_103), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1272(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1273(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1274(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate813(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate814(.a(gate144inter0), .b(s_38), .O(gate144inter1));
  and2  gate815(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate816(.a(s_38), .O(gate144inter3));
  inv1  gate817(.a(s_39), .O(gate144inter4));
  nand2 gate818(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate819(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate820(.a(G468), .O(gate144inter7));
  inv1  gate821(.a(G471), .O(gate144inter8));
  nand2 gate822(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate823(.a(s_39), .b(gate144inter3), .O(gate144inter10));
  nor2  gate824(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate825(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate826(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1709(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1710(.a(gate148inter0), .b(s_166), .O(gate148inter1));
  and2  gate1711(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1712(.a(s_166), .O(gate148inter3));
  inv1  gate1713(.a(s_167), .O(gate148inter4));
  nand2 gate1714(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1715(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1716(.a(G492), .O(gate148inter7));
  inv1  gate1717(.a(G495), .O(gate148inter8));
  nand2 gate1718(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1719(.a(s_167), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1720(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1721(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1722(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1205(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1206(.a(gate155inter0), .b(s_94), .O(gate155inter1));
  and2  gate1207(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1208(.a(s_94), .O(gate155inter3));
  inv1  gate1209(.a(s_95), .O(gate155inter4));
  nand2 gate1210(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1211(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1212(.a(G432), .O(gate155inter7));
  inv1  gate1213(.a(G525), .O(gate155inter8));
  nand2 gate1214(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1215(.a(s_95), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1216(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1217(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1218(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1247(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1248(.a(gate158inter0), .b(s_100), .O(gate158inter1));
  and2  gate1249(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1250(.a(s_100), .O(gate158inter3));
  inv1  gate1251(.a(s_101), .O(gate158inter4));
  nand2 gate1252(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1253(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1254(.a(G441), .O(gate158inter7));
  inv1  gate1255(.a(G528), .O(gate158inter8));
  nand2 gate1256(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1257(.a(s_101), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1258(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1259(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1260(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate743(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate744(.a(gate159inter0), .b(s_28), .O(gate159inter1));
  and2  gate745(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate746(.a(s_28), .O(gate159inter3));
  inv1  gate747(.a(s_29), .O(gate159inter4));
  nand2 gate748(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate749(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate750(.a(G444), .O(gate159inter7));
  inv1  gate751(.a(G531), .O(gate159inter8));
  nand2 gate752(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate753(.a(s_29), .b(gate159inter3), .O(gate159inter10));
  nor2  gate754(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate755(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate756(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate631(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate632(.a(gate162inter0), .b(s_12), .O(gate162inter1));
  and2  gate633(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate634(.a(s_12), .O(gate162inter3));
  inv1  gate635(.a(s_13), .O(gate162inter4));
  nand2 gate636(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate637(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate638(.a(G453), .O(gate162inter7));
  inv1  gate639(.a(G534), .O(gate162inter8));
  nand2 gate640(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate641(.a(s_13), .b(gate162inter3), .O(gate162inter10));
  nor2  gate642(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate643(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate644(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate939(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate940(.a(gate164inter0), .b(s_56), .O(gate164inter1));
  and2  gate941(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate942(.a(s_56), .O(gate164inter3));
  inv1  gate943(.a(s_57), .O(gate164inter4));
  nand2 gate944(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate945(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate946(.a(G459), .O(gate164inter7));
  inv1  gate947(.a(G537), .O(gate164inter8));
  nand2 gate948(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate949(.a(s_57), .b(gate164inter3), .O(gate164inter10));
  nor2  gate950(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate951(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate952(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate1429(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1430(.a(gate165inter0), .b(s_126), .O(gate165inter1));
  and2  gate1431(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1432(.a(s_126), .O(gate165inter3));
  inv1  gate1433(.a(s_127), .O(gate165inter4));
  nand2 gate1434(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1435(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1436(.a(G462), .O(gate165inter7));
  inv1  gate1437(.a(G540), .O(gate165inter8));
  nand2 gate1438(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1439(.a(s_127), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1440(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1441(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1442(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1009(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1010(.a(gate168inter0), .b(s_66), .O(gate168inter1));
  and2  gate1011(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1012(.a(s_66), .O(gate168inter3));
  inv1  gate1013(.a(s_67), .O(gate168inter4));
  nand2 gate1014(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1015(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1016(.a(G471), .O(gate168inter7));
  inv1  gate1017(.a(G543), .O(gate168inter8));
  nand2 gate1018(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1019(.a(s_67), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1020(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1021(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1022(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1317(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1318(.a(gate170inter0), .b(s_110), .O(gate170inter1));
  and2  gate1319(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1320(.a(s_110), .O(gate170inter3));
  inv1  gate1321(.a(s_111), .O(gate170inter4));
  nand2 gate1322(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1323(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1324(.a(G477), .O(gate170inter7));
  inv1  gate1325(.a(G546), .O(gate170inter8));
  nand2 gate1326(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1327(.a(s_111), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1328(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1329(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1330(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate589(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate590(.a(gate171inter0), .b(s_6), .O(gate171inter1));
  and2  gate591(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate592(.a(s_6), .O(gate171inter3));
  inv1  gate593(.a(s_7), .O(gate171inter4));
  nand2 gate594(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate595(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate596(.a(G480), .O(gate171inter7));
  inv1  gate597(.a(G549), .O(gate171inter8));
  nand2 gate598(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate599(.a(s_7), .b(gate171inter3), .O(gate171inter10));
  nor2  gate600(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate601(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate602(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1191(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1192(.a(gate173inter0), .b(s_92), .O(gate173inter1));
  and2  gate1193(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1194(.a(s_92), .O(gate173inter3));
  inv1  gate1195(.a(s_93), .O(gate173inter4));
  nand2 gate1196(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1197(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1198(.a(G486), .O(gate173inter7));
  inv1  gate1199(.a(G552), .O(gate173inter8));
  nand2 gate1200(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1201(.a(s_93), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1202(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1203(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1204(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate603(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate604(.a(gate175inter0), .b(s_8), .O(gate175inter1));
  and2  gate605(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate606(.a(s_8), .O(gate175inter3));
  inv1  gate607(.a(s_9), .O(gate175inter4));
  nand2 gate608(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate609(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate610(.a(G492), .O(gate175inter7));
  inv1  gate611(.a(G555), .O(gate175inter8));
  nand2 gate612(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate613(.a(s_9), .b(gate175inter3), .O(gate175inter10));
  nor2  gate614(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate615(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate616(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate561(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate562(.a(gate187inter0), .b(s_2), .O(gate187inter1));
  and2  gate563(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate564(.a(s_2), .O(gate187inter3));
  inv1  gate565(.a(s_3), .O(gate187inter4));
  nand2 gate566(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate567(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate568(.a(G574), .O(gate187inter7));
  inv1  gate569(.a(G575), .O(gate187inter8));
  nand2 gate570(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate571(.a(s_3), .b(gate187inter3), .O(gate187inter10));
  nor2  gate572(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate573(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate574(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate715(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate716(.a(gate189inter0), .b(s_24), .O(gate189inter1));
  and2  gate717(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate718(.a(s_24), .O(gate189inter3));
  inv1  gate719(.a(s_25), .O(gate189inter4));
  nand2 gate720(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate721(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate722(.a(G578), .O(gate189inter7));
  inv1  gate723(.a(G579), .O(gate189inter8));
  nand2 gate724(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate725(.a(s_25), .b(gate189inter3), .O(gate189inter10));
  nor2  gate726(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate727(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate728(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1079(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1080(.a(gate190inter0), .b(s_76), .O(gate190inter1));
  and2  gate1081(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1082(.a(s_76), .O(gate190inter3));
  inv1  gate1083(.a(s_77), .O(gate190inter4));
  nand2 gate1084(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1085(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1086(.a(G580), .O(gate190inter7));
  inv1  gate1087(.a(G581), .O(gate190inter8));
  nand2 gate1088(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1089(.a(s_77), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1090(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1091(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1092(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate757(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate758(.a(gate191inter0), .b(s_30), .O(gate191inter1));
  and2  gate759(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate760(.a(s_30), .O(gate191inter3));
  inv1  gate761(.a(s_31), .O(gate191inter4));
  nand2 gate762(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate763(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate764(.a(G582), .O(gate191inter7));
  inv1  gate765(.a(G583), .O(gate191inter8));
  nand2 gate766(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate767(.a(s_31), .b(gate191inter3), .O(gate191inter10));
  nor2  gate768(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate769(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate770(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate687(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate688(.a(gate193inter0), .b(s_20), .O(gate193inter1));
  and2  gate689(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate690(.a(s_20), .O(gate193inter3));
  inv1  gate691(.a(s_21), .O(gate193inter4));
  nand2 gate692(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate693(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate694(.a(G586), .O(gate193inter7));
  inv1  gate695(.a(G587), .O(gate193inter8));
  nand2 gate696(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate697(.a(s_21), .b(gate193inter3), .O(gate193inter10));
  nor2  gate698(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate699(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate700(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1569(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1570(.a(gate196inter0), .b(s_146), .O(gate196inter1));
  and2  gate1571(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1572(.a(s_146), .O(gate196inter3));
  inv1  gate1573(.a(s_147), .O(gate196inter4));
  nand2 gate1574(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1575(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1576(.a(G592), .O(gate196inter7));
  inv1  gate1577(.a(G593), .O(gate196inter8));
  nand2 gate1578(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1579(.a(s_147), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1580(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1581(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1582(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1723(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1724(.a(gate199inter0), .b(s_168), .O(gate199inter1));
  and2  gate1725(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1726(.a(s_168), .O(gate199inter3));
  inv1  gate1727(.a(s_169), .O(gate199inter4));
  nand2 gate1728(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1729(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1730(.a(G598), .O(gate199inter7));
  inv1  gate1731(.a(G599), .O(gate199inter8));
  nand2 gate1732(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1733(.a(s_169), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1734(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1735(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1736(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1233(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1234(.a(gate201inter0), .b(s_98), .O(gate201inter1));
  and2  gate1235(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1236(.a(s_98), .O(gate201inter3));
  inv1  gate1237(.a(s_99), .O(gate201inter4));
  nand2 gate1238(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1239(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1240(.a(G602), .O(gate201inter7));
  inv1  gate1241(.a(G607), .O(gate201inter8));
  nand2 gate1242(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1243(.a(s_99), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1244(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1245(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1246(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1065(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1066(.a(gate202inter0), .b(s_74), .O(gate202inter1));
  and2  gate1067(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1068(.a(s_74), .O(gate202inter3));
  inv1  gate1069(.a(s_75), .O(gate202inter4));
  nand2 gate1070(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1071(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1072(.a(G612), .O(gate202inter7));
  inv1  gate1073(.a(G617), .O(gate202inter8));
  nand2 gate1074(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1075(.a(s_75), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1076(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1077(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1078(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1793(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1794(.a(gate216inter0), .b(s_178), .O(gate216inter1));
  and2  gate1795(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1796(.a(s_178), .O(gate216inter3));
  inv1  gate1797(.a(s_179), .O(gate216inter4));
  nand2 gate1798(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1799(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1800(.a(G617), .O(gate216inter7));
  inv1  gate1801(.a(G675), .O(gate216inter8));
  nand2 gate1802(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1803(.a(s_179), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1804(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1805(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1806(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate925(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate926(.a(gate217inter0), .b(s_54), .O(gate217inter1));
  and2  gate927(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate928(.a(s_54), .O(gate217inter3));
  inv1  gate929(.a(s_55), .O(gate217inter4));
  nand2 gate930(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate931(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate932(.a(G622), .O(gate217inter7));
  inv1  gate933(.a(G678), .O(gate217inter8));
  nand2 gate934(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate935(.a(s_55), .b(gate217inter3), .O(gate217inter10));
  nor2  gate936(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate937(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate938(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1373(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1374(.a(gate218inter0), .b(s_118), .O(gate218inter1));
  and2  gate1375(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1376(.a(s_118), .O(gate218inter3));
  inv1  gate1377(.a(s_119), .O(gate218inter4));
  nand2 gate1378(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1379(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1380(.a(G627), .O(gate218inter7));
  inv1  gate1381(.a(G678), .O(gate218inter8));
  nand2 gate1382(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1383(.a(s_119), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1384(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1385(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1386(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate911(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate912(.a(gate229inter0), .b(s_52), .O(gate229inter1));
  and2  gate913(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate914(.a(s_52), .O(gate229inter3));
  inv1  gate915(.a(s_53), .O(gate229inter4));
  nand2 gate916(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate917(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate918(.a(G698), .O(gate229inter7));
  inv1  gate919(.a(G699), .O(gate229inter8));
  nand2 gate920(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate921(.a(s_53), .b(gate229inter3), .O(gate229inter10));
  nor2  gate922(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate923(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate924(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate729(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate730(.a(gate236inter0), .b(s_26), .O(gate236inter1));
  and2  gate731(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate732(.a(s_26), .O(gate236inter3));
  inv1  gate733(.a(s_27), .O(gate236inter4));
  nand2 gate734(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate735(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate736(.a(G251), .O(gate236inter7));
  inv1  gate737(.a(G727), .O(gate236inter8));
  nand2 gate738(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate739(.a(s_27), .b(gate236inter3), .O(gate236inter10));
  nor2  gate740(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate741(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate742(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1555(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1556(.a(gate246inter0), .b(s_144), .O(gate246inter1));
  and2  gate1557(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1558(.a(s_144), .O(gate246inter3));
  inv1  gate1559(.a(s_145), .O(gate246inter4));
  nand2 gate1560(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1561(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1562(.a(G724), .O(gate246inter7));
  inv1  gate1563(.a(G736), .O(gate246inter8));
  nand2 gate1564(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1565(.a(s_145), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1566(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1567(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1568(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate953(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate954(.a(gate248inter0), .b(s_58), .O(gate248inter1));
  and2  gate955(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate956(.a(s_58), .O(gate248inter3));
  inv1  gate957(.a(s_59), .O(gate248inter4));
  nand2 gate958(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate959(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate960(.a(G727), .O(gate248inter7));
  inv1  gate961(.a(G739), .O(gate248inter8));
  nand2 gate962(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate963(.a(s_59), .b(gate248inter3), .O(gate248inter10));
  nor2  gate964(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate965(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate966(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1947(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1948(.a(gate255inter0), .b(s_200), .O(gate255inter1));
  and2  gate1949(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1950(.a(s_200), .O(gate255inter3));
  inv1  gate1951(.a(s_201), .O(gate255inter4));
  nand2 gate1952(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1953(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1954(.a(G263), .O(gate255inter7));
  inv1  gate1955(.a(G751), .O(gate255inter8));
  nand2 gate1956(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1957(.a(s_201), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1958(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1959(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1960(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1779(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1780(.a(gate256inter0), .b(s_176), .O(gate256inter1));
  and2  gate1781(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1782(.a(s_176), .O(gate256inter3));
  inv1  gate1783(.a(s_177), .O(gate256inter4));
  nand2 gate1784(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1785(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1786(.a(G715), .O(gate256inter7));
  inv1  gate1787(.a(G751), .O(gate256inter8));
  nand2 gate1788(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1789(.a(s_177), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1790(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1791(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1792(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1275(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1276(.a(gate260inter0), .b(s_104), .O(gate260inter1));
  and2  gate1277(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1278(.a(s_104), .O(gate260inter3));
  inv1  gate1279(.a(s_105), .O(gate260inter4));
  nand2 gate1280(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1281(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1282(.a(G760), .O(gate260inter7));
  inv1  gate1283(.a(G761), .O(gate260inter8));
  nand2 gate1284(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1285(.a(s_105), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1286(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1287(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1288(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate701(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate702(.a(gate262inter0), .b(s_22), .O(gate262inter1));
  and2  gate703(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate704(.a(s_22), .O(gate262inter3));
  inv1  gate705(.a(s_23), .O(gate262inter4));
  nand2 gate706(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate707(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate708(.a(G764), .O(gate262inter7));
  inv1  gate709(.a(G765), .O(gate262inter8));
  nand2 gate710(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate711(.a(s_23), .b(gate262inter3), .O(gate262inter10));
  nor2  gate712(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate713(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate714(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1597(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1598(.a(gate264inter0), .b(s_150), .O(gate264inter1));
  and2  gate1599(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1600(.a(s_150), .O(gate264inter3));
  inv1  gate1601(.a(s_151), .O(gate264inter4));
  nand2 gate1602(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1603(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1604(.a(G768), .O(gate264inter7));
  inv1  gate1605(.a(G769), .O(gate264inter8));
  nand2 gate1606(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1607(.a(s_151), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1608(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1609(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1610(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate659(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate660(.a(gate269inter0), .b(s_16), .O(gate269inter1));
  and2  gate661(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate662(.a(s_16), .O(gate269inter3));
  inv1  gate663(.a(s_17), .O(gate269inter4));
  nand2 gate664(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate665(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate666(.a(G654), .O(gate269inter7));
  inv1  gate667(.a(G782), .O(gate269inter8));
  nand2 gate668(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate669(.a(s_17), .b(gate269inter3), .O(gate269inter10));
  nor2  gate670(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate671(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate672(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate1835(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1836(.a(gate270inter0), .b(s_184), .O(gate270inter1));
  and2  gate1837(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1838(.a(s_184), .O(gate270inter3));
  inv1  gate1839(.a(s_185), .O(gate270inter4));
  nand2 gate1840(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1841(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1842(.a(G657), .O(gate270inter7));
  inv1  gate1843(.a(G785), .O(gate270inter8));
  nand2 gate1844(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1845(.a(s_185), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1846(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1847(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1848(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1121(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1122(.a(gate274inter0), .b(s_82), .O(gate274inter1));
  and2  gate1123(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1124(.a(s_82), .O(gate274inter3));
  inv1  gate1125(.a(s_83), .O(gate274inter4));
  nand2 gate1126(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1127(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1128(.a(G770), .O(gate274inter7));
  inv1  gate1129(.a(G794), .O(gate274inter8));
  nand2 gate1130(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1131(.a(s_83), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1132(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1133(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1134(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1653(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1654(.a(gate282inter0), .b(s_158), .O(gate282inter1));
  and2  gate1655(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1656(.a(s_158), .O(gate282inter3));
  inv1  gate1657(.a(s_159), .O(gate282inter4));
  nand2 gate1658(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1659(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1660(.a(G782), .O(gate282inter7));
  inv1  gate1661(.a(G806), .O(gate282inter8));
  nand2 gate1662(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1663(.a(s_159), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1664(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1665(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1666(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1667(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1668(.a(gate289inter0), .b(s_160), .O(gate289inter1));
  and2  gate1669(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1670(.a(s_160), .O(gate289inter3));
  inv1  gate1671(.a(s_161), .O(gate289inter4));
  nand2 gate1672(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1673(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1674(.a(G818), .O(gate289inter7));
  inv1  gate1675(.a(G819), .O(gate289inter8));
  nand2 gate1676(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1677(.a(s_161), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1678(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1679(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1680(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1751(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1752(.a(gate388inter0), .b(s_172), .O(gate388inter1));
  and2  gate1753(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1754(.a(s_172), .O(gate388inter3));
  inv1  gate1755(.a(s_173), .O(gate388inter4));
  nand2 gate1756(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1757(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1758(.a(G2), .O(gate388inter7));
  inv1  gate1759(.a(G1039), .O(gate388inter8));
  nand2 gate1760(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1761(.a(s_173), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1762(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1763(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1764(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate645(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate646(.a(gate397inter0), .b(s_14), .O(gate397inter1));
  and2  gate647(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate648(.a(s_14), .O(gate397inter3));
  inv1  gate649(.a(s_15), .O(gate397inter4));
  nand2 gate650(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate651(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate652(.a(G11), .O(gate397inter7));
  inv1  gate653(.a(G1066), .O(gate397inter8));
  nand2 gate654(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate655(.a(s_15), .b(gate397inter3), .O(gate397inter10));
  nor2  gate656(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate657(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate658(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1051(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1052(.a(gate405inter0), .b(s_72), .O(gate405inter1));
  and2  gate1053(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1054(.a(s_72), .O(gate405inter3));
  inv1  gate1055(.a(s_73), .O(gate405inter4));
  nand2 gate1056(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1057(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1058(.a(G19), .O(gate405inter7));
  inv1  gate1059(.a(G1090), .O(gate405inter8));
  nand2 gate1060(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1061(.a(s_73), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1062(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1063(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1064(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1891(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1892(.a(gate407inter0), .b(s_192), .O(gate407inter1));
  and2  gate1893(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1894(.a(s_192), .O(gate407inter3));
  inv1  gate1895(.a(s_193), .O(gate407inter4));
  nand2 gate1896(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1897(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1898(.a(G21), .O(gate407inter7));
  inv1  gate1899(.a(G1096), .O(gate407inter8));
  nand2 gate1900(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1901(.a(s_193), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1902(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1903(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1904(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1625(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1626(.a(gate410inter0), .b(s_154), .O(gate410inter1));
  and2  gate1627(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1628(.a(s_154), .O(gate410inter3));
  inv1  gate1629(.a(s_155), .O(gate410inter4));
  nand2 gate1630(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1631(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1632(.a(G24), .O(gate410inter7));
  inv1  gate1633(.a(G1105), .O(gate410inter8));
  nand2 gate1634(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1635(.a(s_155), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1636(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1637(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1638(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1457(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1458(.a(gate411inter0), .b(s_130), .O(gate411inter1));
  and2  gate1459(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1460(.a(s_130), .O(gate411inter3));
  inv1  gate1461(.a(s_131), .O(gate411inter4));
  nand2 gate1462(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1463(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1464(.a(G25), .O(gate411inter7));
  inv1  gate1465(.a(G1108), .O(gate411inter8));
  nand2 gate1466(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1467(.a(s_131), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1468(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1469(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1470(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1933(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1934(.a(gate416inter0), .b(s_198), .O(gate416inter1));
  and2  gate1935(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1936(.a(s_198), .O(gate416inter3));
  inv1  gate1937(.a(s_199), .O(gate416inter4));
  nand2 gate1938(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1939(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1940(.a(G30), .O(gate416inter7));
  inv1  gate1941(.a(G1123), .O(gate416inter8));
  nand2 gate1942(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1943(.a(s_199), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1944(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1945(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1946(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1513(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1514(.a(gate418inter0), .b(s_138), .O(gate418inter1));
  and2  gate1515(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1516(.a(s_138), .O(gate418inter3));
  inv1  gate1517(.a(s_139), .O(gate418inter4));
  nand2 gate1518(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1519(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1520(.a(G32), .O(gate418inter7));
  inv1  gate1521(.a(G1129), .O(gate418inter8));
  nand2 gate1522(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1523(.a(s_139), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1524(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1525(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1526(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1737(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1738(.a(gate422inter0), .b(s_170), .O(gate422inter1));
  and2  gate1739(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1740(.a(s_170), .O(gate422inter3));
  inv1  gate1741(.a(s_171), .O(gate422inter4));
  nand2 gate1742(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1743(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1744(.a(G1039), .O(gate422inter7));
  inv1  gate1745(.a(G1135), .O(gate422inter8));
  nand2 gate1746(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1747(.a(s_171), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1748(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1749(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1750(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1303(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1304(.a(gate423inter0), .b(s_108), .O(gate423inter1));
  and2  gate1305(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1306(.a(s_108), .O(gate423inter3));
  inv1  gate1307(.a(s_109), .O(gate423inter4));
  nand2 gate1308(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1309(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1310(.a(G3), .O(gate423inter7));
  inv1  gate1311(.a(G1138), .O(gate423inter8));
  nand2 gate1312(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1313(.a(s_109), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1314(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1315(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1316(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate547(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate548(.a(gate424inter0), .b(s_0), .O(gate424inter1));
  and2  gate549(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate550(.a(s_0), .O(gate424inter3));
  inv1  gate551(.a(s_1), .O(gate424inter4));
  nand2 gate552(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate553(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate554(.a(G1042), .O(gate424inter7));
  inv1  gate555(.a(G1138), .O(gate424inter8));
  nand2 gate556(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate557(.a(s_1), .b(gate424inter3), .O(gate424inter10));
  nor2  gate558(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate559(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate560(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1037(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1038(.a(gate436inter0), .b(s_70), .O(gate436inter1));
  and2  gate1039(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1040(.a(s_70), .O(gate436inter3));
  inv1  gate1041(.a(s_71), .O(gate436inter4));
  nand2 gate1042(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1043(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1044(.a(G1060), .O(gate436inter7));
  inv1  gate1045(.a(G1156), .O(gate436inter8));
  nand2 gate1046(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1047(.a(s_71), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1048(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1049(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1050(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1289(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1290(.a(gate437inter0), .b(s_106), .O(gate437inter1));
  and2  gate1291(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1292(.a(s_106), .O(gate437inter3));
  inv1  gate1293(.a(s_107), .O(gate437inter4));
  nand2 gate1294(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1295(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1296(.a(G10), .O(gate437inter7));
  inv1  gate1297(.a(G1159), .O(gate437inter8));
  nand2 gate1298(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1299(.a(s_107), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1300(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1301(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1302(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1849(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1850(.a(gate439inter0), .b(s_186), .O(gate439inter1));
  and2  gate1851(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1852(.a(s_186), .O(gate439inter3));
  inv1  gate1853(.a(s_187), .O(gate439inter4));
  nand2 gate1854(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1855(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1856(.a(G11), .O(gate439inter7));
  inv1  gate1857(.a(G1162), .O(gate439inter8));
  nand2 gate1858(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1859(.a(s_187), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1860(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1861(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1862(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1135(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1136(.a(gate443inter0), .b(s_84), .O(gate443inter1));
  and2  gate1137(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1138(.a(s_84), .O(gate443inter3));
  inv1  gate1139(.a(s_85), .O(gate443inter4));
  nand2 gate1140(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1141(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1142(.a(G13), .O(gate443inter7));
  inv1  gate1143(.a(G1168), .O(gate443inter8));
  nand2 gate1144(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1145(.a(s_85), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1146(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1147(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1148(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1821(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1822(.a(gate447inter0), .b(s_182), .O(gate447inter1));
  and2  gate1823(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1824(.a(s_182), .O(gate447inter3));
  inv1  gate1825(.a(s_183), .O(gate447inter4));
  nand2 gate1826(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1827(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1828(.a(G15), .O(gate447inter7));
  inv1  gate1829(.a(G1174), .O(gate447inter8));
  nand2 gate1830(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1831(.a(s_183), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1832(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1833(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1834(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate771(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate772(.a(gate452inter0), .b(s_32), .O(gate452inter1));
  and2  gate773(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate774(.a(s_32), .O(gate452inter3));
  inv1  gate775(.a(s_33), .O(gate452inter4));
  nand2 gate776(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate777(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate778(.a(G1084), .O(gate452inter7));
  inv1  gate779(.a(G1180), .O(gate452inter8));
  nand2 gate780(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate781(.a(s_33), .b(gate452inter3), .O(gate452inter10));
  nor2  gate782(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate783(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate784(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1681(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1682(.a(gate459inter0), .b(s_162), .O(gate459inter1));
  and2  gate1683(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1684(.a(s_162), .O(gate459inter3));
  inv1  gate1685(.a(s_163), .O(gate459inter4));
  nand2 gate1686(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1687(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1688(.a(G21), .O(gate459inter7));
  inv1  gate1689(.a(G1192), .O(gate459inter8));
  nand2 gate1690(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1691(.a(s_163), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1692(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1693(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1694(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1149(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1150(.a(gate465inter0), .b(s_86), .O(gate465inter1));
  and2  gate1151(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1152(.a(s_86), .O(gate465inter3));
  inv1  gate1153(.a(s_87), .O(gate465inter4));
  nand2 gate1154(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1155(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1156(.a(G24), .O(gate465inter7));
  inv1  gate1157(.a(G1201), .O(gate465inter8));
  nand2 gate1158(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1159(.a(s_87), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1160(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1161(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1162(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate883(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate884(.a(gate471inter0), .b(s_48), .O(gate471inter1));
  and2  gate885(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate886(.a(s_48), .O(gate471inter3));
  inv1  gate887(.a(s_49), .O(gate471inter4));
  nand2 gate888(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate889(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate890(.a(G27), .O(gate471inter7));
  inv1  gate891(.a(G1210), .O(gate471inter8));
  nand2 gate892(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate893(.a(s_49), .b(gate471inter3), .O(gate471inter10));
  nor2  gate894(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate895(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate896(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate897(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate898(.a(gate480inter0), .b(s_50), .O(gate480inter1));
  and2  gate899(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate900(.a(s_50), .O(gate480inter3));
  inv1  gate901(.a(s_51), .O(gate480inter4));
  nand2 gate902(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate903(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate904(.a(G1126), .O(gate480inter7));
  inv1  gate905(.a(G1222), .O(gate480inter8));
  nand2 gate906(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate907(.a(s_51), .b(gate480inter3), .O(gate480inter10));
  nor2  gate908(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate909(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate910(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1905(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1906(.a(gate487inter0), .b(s_194), .O(gate487inter1));
  and2  gate1907(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1908(.a(s_194), .O(gate487inter3));
  inv1  gate1909(.a(s_195), .O(gate487inter4));
  nand2 gate1910(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1911(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1912(.a(G1236), .O(gate487inter7));
  inv1  gate1913(.a(G1237), .O(gate487inter8));
  nand2 gate1914(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1915(.a(s_195), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1916(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1917(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1918(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1107(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1108(.a(gate490inter0), .b(s_80), .O(gate490inter1));
  and2  gate1109(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1110(.a(s_80), .O(gate490inter3));
  inv1  gate1111(.a(s_81), .O(gate490inter4));
  nand2 gate1112(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1113(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1114(.a(G1242), .O(gate490inter7));
  inv1  gate1115(.a(G1243), .O(gate490inter8));
  nand2 gate1116(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1117(.a(s_81), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1118(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1119(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1120(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate617(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate618(.a(gate493inter0), .b(s_10), .O(gate493inter1));
  and2  gate619(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate620(.a(s_10), .O(gate493inter3));
  inv1  gate621(.a(s_11), .O(gate493inter4));
  nand2 gate622(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate623(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate624(.a(G1248), .O(gate493inter7));
  inv1  gate625(.a(G1249), .O(gate493inter8));
  nand2 gate626(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate627(.a(s_11), .b(gate493inter3), .O(gate493inter10));
  nor2  gate628(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate629(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate630(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1471(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1472(.a(gate494inter0), .b(s_132), .O(gate494inter1));
  and2  gate1473(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1474(.a(s_132), .O(gate494inter3));
  inv1  gate1475(.a(s_133), .O(gate494inter4));
  nand2 gate1476(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1477(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1478(.a(G1250), .O(gate494inter7));
  inv1  gate1479(.a(G1251), .O(gate494inter8));
  nand2 gate1480(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1481(.a(s_133), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1482(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1483(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1484(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1485(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1486(.a(gate506inter0), .b(s_134), .O(gate506inter1));
  and2  gate1487(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1488(.a(s_134), .O(gate506inter3));
  inv1  gate1489(.a(s_135), .O(gate506inter4));
  nand2 gate1490(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1491(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1492(.a(G1274), .O(gate506inter7));
  inv1  gate1493(.a(G1275), .O(gate506inter8));
  nand2 gate1494(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1495(.a(s_135), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1496(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1497(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1498(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1387(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1388(.a(gate507inter0), .b(s_120), .O(gate507inter1));
  and2  gate1389(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1390(.a(s_120), .O(gate507inter3));
  inv1  gate1391(.a(s_121), .O(gate507inter4));
  nand2 gate1392(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1393(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1394(.a(G1276), .O(gate507inter7));
  inv1  gate1395(.a(G1277), .O(gate507inter8));
  nand2 gate1396(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1397(.a(s_121), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1398(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1399(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1400(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1163(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1164(.a(gate509inter0), .b(s_88), .O(gate509inter1));
  and2  gate1165(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1166(.a(s_88), .O(gate509inter3));
  inv1  gate1167(.a(s_89), .O(gate509inter4));
  nand2 gate1168(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1169(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1170(.a(G1280), .O(gate509inter7));
  inv1  gate1171(.a(G1281), .O(gate509inter8));
  nand2 gate1172(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1173(.a(s_89), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1174(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1175(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1176(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule