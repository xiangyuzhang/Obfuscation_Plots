module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381, s_382, s_383, s_384, s_385, s_386, s_387, s_388, s_389, s_390, s_391;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate939(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate940(.a(gate12inter0), .b(s_56), .O(gate12inter1));
  and2  gate941(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate942(.a(s_56), .O(gate12inter3));
  inv1  gate943(.a(s_57), .O(gate12inter4));
  nand2 gate944(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate945(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate946(.a(G7), .O(gate12inter7));
  inv1  gate947(.a(G8), .O(gate12inter8));
  nand2 gate948(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate949(.a(s_57), .b(gate12inter3), .O(gate12inter10));
  nor2  gate950(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate951(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate952(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2787(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2788(.a(gate13inter0), .b(s_320), .O(gate13inter1));
  and2  gate2789(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2790(.a(s_320), .O(gate13inter3));
  inv1  gate2791(.a(s_321), .O(gate13inter4));
  nand2 gate2792(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2793(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2794(.a(G9), .O(gate13inter7));
  inv1  gate2795(.a(G10), .O(gate13inter8));
  nand2 gate2796(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2797(.a(s_321), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2798(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2799(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2800(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1583(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1584(.a(gate14inter0), .b(s_148), .O(gate14inter1));
  and2  gate1585(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1586(.a(s_148), .O(gate14inter3));
  inv1  gate1587(.a(s_149), .O(gate14inter4));
  nand2 gate1588(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1589(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1590(.a(G11), .O(gate14inter7));
  inv1  gate1591(.a(G12), .O(gate14inter8));
  nand2 gate1592(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1593(.a(s_149), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1594(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1595(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1596(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2913(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2914(.a(gate16inter0), .b(s_338), .O(gate16inter1));
  and2  gate2915(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2916(.a(s_338), .O(gate16inter3));
  inv1  gate2917(.a(s_339), .O(gate16inter4));
  nand2 gate2918(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2919(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2920(.a(G15), .O(gate16inter7));
  inv1  gate2921(.a(G16), .O(gate16inter8));
  nand2 gate2922(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2923(.a(s_339), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2924(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2925(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2926(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate701(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate702(.a(gate19inter0), .b(s_22), .O(gate19inter1));
  and2  gate703(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate704(.a(s_22), .O(gate19inter3));
  inv1  gate705(.a(s_23), .O(gate19inter4));
  nand2 gate706(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate707(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate708(.a(G21), .O(gate19inter7));
  inv1  gate709(.a(G22), .O(gate19inter8));
  nand2 gate710(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate711(.a(s_23), .b(gate19inter3), .O(gate19inter10));
  nor2  gate712(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate713(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate714(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate3249(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate3250(.a(gate23inter0), .b(s_386), .O(gate23inter1));
  and2  gate3251(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate3252(.a(s_386), .O(gate23inter3));
  inv1  gate3253(.a(s_387), .O(gate23inter4));
  nand2 gate3254(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate3255(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate3256(.a(G29), .O(gate23inter7));
  inv1  gate3257(.a(G30), .O(gate23inter8));
  nand2 gate3258(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate3259(.a(s_387), .b(gate23inter3), .O(gate23inter10));
  nor2  gate3260(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate3261(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate3262(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2087(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2088(.a(gate24inter0), .b(s_220), .O(gate24inter1));
  and2  gate2089(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2090(.a(s_220), .O(gate24inter3));
  inv1  gate2091(.a(s_221), .O(gate24inter4));
  nand2 gate2092(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2093(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2094(.a(G31), .O(gate24inter7));
  inv1  gate2095(.a(G32), .O(gate24inter8));
  nand2 gate2096(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2097(.a(s_221), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2098(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2099(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2100(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate659(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate660(.a(gate25inter0), .b(s_16), .O(gate25inter1));
  and2  gate661(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate662(.a(s_16), .O(gate25inter3));
  inv1  gate663(.a(s_17), .O(gate25inter4));
  nand2 gate664(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate665(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate666(.a(G1), .O(gate25inter7));
  inv1  gate667(.a(G5), .O(gate25inter8));
  nand2 gate668(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate669(.a(s_17), .b(gate25inter3), .O(gate25inter10));
  nor2  gate670(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate671(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate672(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate3053(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate3054(.a(gate35inter0), .b(s_358), .O(gate35inter1));
  and2  gate3055(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate3056(.a(s_358), .O(gate35inter3));
  inv1  gate3057(.a(s_359), .O(gate35inter4));
  nand2 gate3058(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate3059(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate3060(.a(G18), .O(gate35inter7));
  inv1  gate3061(.a(G22), .O(gate35inter8));
  nand2 gate3062(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate3063(.a(s_359), .b(gate35inter3), .O(gate35inter10));
  nor2  gate3064(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate3065(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate3066(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2325(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2326(.a(gate36inter0), .b(s_254), .O(gate36inter1));
  and2  gate2327(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2328(.a(s_254), .O(gate36inter3));
  inv1  gate2329(.a(s_255), .O(gate36inter4));
  nand2 gate2330(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2331(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2332(.a(G26), .O(gate36inter7));
  inv1  gate2333(.a(G30), .O(gate36inter8));
  nand2 gate2334(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2335(.a(s_255), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2336(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2337(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2338(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate3193(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate3194(.a(gate37inter0), .b(s_378), .O(gate37inter1));
  and2  gate3195(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate3196(.a(s_378), .O(gate37inter3));
  inv1  gate3197(.a(s_379), .O(gate37inter4));
  nand2 gate3198(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate3199(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate3200(.a(G19), .O(gate37inter7));
  inv1  gate3201(.a(G23), .O(gate37inter8));
  nand2 gate3202(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate3203(.a(s_379), .b(gate37inter3), .O(gate37inter10));
  nor2  gate3204(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate3205(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate3206(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate841(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate842(.a(gate39inter0), .b(s_42), .O(gate39inter1));
  and2  gate843(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate844(.a(s_42), .O(gate39inter3));
  inv1  gate845(.a(s_43), .O(gate39inter4));
  nand2 gate846(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate847(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate848(.a(G20), .O(gate39inter7));
  inv1  gate849(.a(G24), .O(gate39inter8));
  nand2 gate850(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate851(.a(s_43), .b(gate39inter3), .O(gate39inter10));
  nor2  gate852(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate853(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate854(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate2871(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2872(.a(gate40inter0), .b(s_332), .O(gate40inter1));
  and2  gate2873(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2874(.a(s_332), .O(gate40inter3));
  inv1  gate2875(.a(s_333), .O(gate40inter4));
  nand2 gate2876(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2877(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2878(.a(G28), .O(gate40inter7));
  inv1  gate2879(.a(G32), .O(gate40inter8));
  nand2 gate2880(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2881(.a(s_333), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2882(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2883(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2884(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2605(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2606(.a(gate42inter0), .b(s_294), .O(gate42inter1));
  and2  gate2607(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2608(.a(s_294), .O(gate42inter3));
  inv1  gate2609(.a(s_295), .O(gate42inter4));
  nand2 gate2610(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2611(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2612(.a(G2), .O(gate42inter7));
  inv1  gate2613(.a(G266), .O(gate42inter8));
  nand2 gate2614(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2615(.a(s_295), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2616(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2617(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2618(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate3235(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate3236(.a(gate45inter0), .b(s_384), .O(gate45inter1));
  and2  gate3237(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate3238(.a(s_384), .O(gate45inter3));
  inv1  gate3239(.a(s_385), .O(gate45inter4));
  nand2 gate3240(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate3241(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate3242(.a(G5), .O(gate45inter7));
  inv1  gate3243(.a(G272), .O(gate45inter8));
  nand2 gate3244(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate3245(.a(s_385), .b(gate45inter3), .O(gate45inter10));
  nor2  gate3246(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate3247(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate3248(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2969(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2970(.a(gate48inter0), .b(s_346), .O(gate48inter1));
  and2  gate2971(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2972(.a(s_346), .O(gate48inter3));
  inv1  gate2973(.a(s_347), .O(gate48inter4));
  nand2 gate2974(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2975(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2976(.a(G8), .O(gate48inter7));
  inv1  gate2977(.a(G275), .O(gate48inter8));
  nand2 gate2978(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2979(.a(s_347), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2980(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2981(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2982(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1065(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1066(.a(gate53inter0), .b(s_74), .O(gate53inter1));
  and2  gate1067(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1068(.a(s_74), .O(gate53inter3));
  inv1  gate1069(.a(s_75), .O(gate53inter4));
  nand2 gate1070(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1071(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1072(.a(G13), .O(gate53inter7));
  inv1  gate1073(.a(G284), .O(gate53inter8));
  nand2 gate1074(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1075(.a(s_75), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1076(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1077(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1078(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate2619(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2620(.a(gate54inter0), .b(s_296), .O(gate54inter1));
  and2  gate2621(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2622(.a(s_296), .O(gate54inter3));
  inv1  gate2623(.a(s_297), .O(gate54inter4));
  nand2 gate2624(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2625(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2626(.a(G14), .O(gate54inter7));
  inv1  gate2627(.a(G284), .O(gate54inter8));
  nand2 gate2628(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2629(.a(s_297), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2630(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2631(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2632(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1247(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1248(.a(gate55inter0), .b(s_100), .O(gate55inter1));
  and2  gate1249(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1250(.a(s_100), .O(gate55inter3));
  inv1  gate1251(.a(s_101), .O(gate55inter4));
  nand2 gate1252(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1253(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1254(.a(G15), .O(gate55inter7));
  inv1  gate1255(.a(G287), .O(gate55inter8));
  nand2 gate1256(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1257(.a(s_101), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1258(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1259(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1260(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1625(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1626(.a(gate57inter0), .b(s_154), .O(gate57inter1));
  and2  gate1627(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1628(.a(s_154), .O(gate57inter3));
  inv1  gate1629(.a(s_155), .O(gate57inter4));
  nand2 gate1630(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1631(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1632(.a(G17), .O(gate57inter7));
  inv1  gate1633(.a(G290), .O(gate57inter8));
  nand2 gate1634(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1635(.a(s_155), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1636(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1637(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1638(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate995(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate996(.a(gate59inter0), .b(s_64), .O(gate59inter1));
  and2  gate997(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate998(.a(s_64), .O(gate59inter3));
  inv1  gate999(.a(s_65), .O(gate59inter4));
  nand2 gate1000(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1001(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1002(.a(G19), .O(gate59inter7));
  inv1  gate1003(.a(G293), .O(gate59inter8));
  nand2 gate1004(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1005(.a(s_65), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1006(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1007(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1008(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate2955(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2956(.a(gate60inter0), .b(s_344), .O(gate60inter1));
  and2  gate2957(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2958(.a(s_344), .O(gate60inter3));
  inv1  gate2959(.a(s_345), .O(gate60inter4));
  nand2 gate2960(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2961(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2962(.a(G20), .O(gate60inter7));
  inv1  gate2963(.a(G293), .O(gate60inter8));
  nand2 gate2964(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2965(.a(s_345), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2966(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2967(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2968(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2157(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2158(.a(gate61inter0), .b(s_230), .O(gate61inter1));
  and2  gate2159(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2160(.a(s_230), .O(gate61inter3));
  inv1  gate2161(.a(s_231), .O(gate61inter4));
  nand2 gate2162(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2163(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2164(.a(G21), .O(gate61inter7));
  inv1  gate2165(.a(G296), .O(gate61inter8));
  nand2 gate2166(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2167(.a(s_231), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2168(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2169(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2170(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1723(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1724(.a(gate62inter0), .b(s_168), .O(gate62inter1));
  and2  gate1725(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1726(.a(s_168), .O(gate62inter3));
  inv1  gate1727(.a(s_169), .O(gate62inter4));
  nand2 gate1728(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1729(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1730(.a(G22), .O(gate62inter7));
  inv1  gate1731(.a(G296), .O(gate62inter8));
  nand2 gate1732(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1733(.a(s_169), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1734(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1735(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1736(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1919(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1920(.a(gate64inter0), .b(s_196), .O(gate64inter1));
  and2  gate1921(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1922(.a(s_196), .O(gate64inter3));
  inv1  gate1923(.a(s_197), .O(gate64inter4));
  nand2 gate1924(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1925(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1926(.a(G24), .O(gate64inter7));
  inv1  gate1927(.a(G299), .O(gate64inter8));
  nand2 gate1928(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1929(.a(s_197), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1930(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1931(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1932(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate2549(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2550(.a(gate65inter0), .b(s_286), .O(gate65inter1));
  and2  gate2551(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2552(.a(s_286), .O(gate65inter3));
  inv1  gate2553(.a(s_287), .O(gate65inter4));
  nand2 gate2554(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2555(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2556(.a(G25), .O(gate65inter7));
  inv1  gate2557(.a(G302), .O(gate65inter8));
  nand2 gate2558(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2559(.a(s_287), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2560(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2561(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2562(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate589(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate590(.a(gate67inter0), .b(s_6), .O(gate67inter1));
  and2  gate591(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate592(.a(s_6), .O(gate67inter3));
  inv1  gate593(.a(s_7), .O(gate67inter4));
  nand2 gate594(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate595(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate596(.a(G27), .O(gate67inter7));
  inv1  gate597(.a(G305), .O(gate67inter8));
  nand2 gate598(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate599(.a(s_7), .b(gate67inter3), .O(gate67inter10));
  nor2  gate600(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate601(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate602(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate3165(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate3166(.a(gate71inter0), .b(s_374), .O(gate71inter1));
  and2  gate3167(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate3168(.a(s_374), .O(gate71inter3));
  inv1  gate3169(.a(s_375), .O(gate71inter4));
  nand2 gate3170(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate3171(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate3172(.a(G31), .O(gate71inter7));
  inv1  gate3173(.a(G311), .O(gate71inter8));
  nand2 gate3174(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate3175(.a(s_375), .b(gate71inter3), .O(gate71inter10));
  nor2  gate3176(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate3177(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate3178(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate2675(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2676(.a(gate73inter0), .b(s_304), .O(gate73inter1));
  and2  gate2677(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2678(.a(s_304), .O(gate73inter3));
  inv1  gate2679(.a(s_305), .O(gate73inter4));
  nand2 gate2680(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2681(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2682(.a(G1), .O(gate73inter7));
  inv1  gate2683(.a(G314), .O(gate73inter8));
  nand2 gate2684(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2685(.a(s_305), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2686(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2687(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2688(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2591(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2592(.a(gate76inter0), .b(s_292), .O(gate76inter1));
  and2  gate2593(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2594(.a(s_292), .O(gate76inter3));
  inv1  gate2595(.a(s_293), .O(gate76inter4));
  nand2 gate2596(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2597(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2598(.a(G13), .O(gate76inter7));
  inv1  gate2599(.a(G317), .O(gate76inter8));
  nand2 gate2600(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2601(.a(s_293), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2602(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2603(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2604(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2773(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2774(.a(gate78inter0), .b(s_318), .O(gate78inter1));
  and2  gate2775(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2776(.a(s_318), .O(gate78inter3));
  inv1  gate2777(.a(s_319), .O(gate78inter4));
  nand2 gate2778(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2779(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2780(.a(G6), .O(gate78inter7));
  inv1  gate2781(.a(G320), .O(gate78inter8));
  nand2 gate2782(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2783(.a(s_319), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2784(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2785(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2786(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1821(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1822(.a(gate79inter0), .b(s_182), .O(gate79inter1));
  and2  gate1823(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1824(.a(s_182), .O(gate79inter3));
  inv1  gate1825(.a(s_183), .O(gate79inter4));
  nand2 gate1826(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1827(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1828(.a(G10), .O(gate79inter7));
  inv1  gate1829(.a(G323), .O(gate79inter8));
  nand2 gate1830(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1831(.a(s_183), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1832(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1833(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1834(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate897(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate898(.a(gate80inter0), .b(s_50), .O(gate80inter1));
  and2  gate899(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate900(.a(s_50), .O(gate80inter3));
  inv1  gate901(.a(s_51), .O(gate80inter4));
  nand2 gate902(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate903(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate904(.a(G14), .O(gate80inter7));
  inv1  gate905(.a(G323), .O(gate80inter8));
  nand2 gate906(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate907(.a(s_51), .b(gate80inter3), .O(gate80inter10));
  nor2  gate908(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate909(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate910(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate673(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate674(.a(gate82inter0), .b(s_18), .O(gate82inter1));
  and2  gate675(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate676(.a(s_18), .O(gate82inter3));
  inv1  gate677(.a(s_19), .O(gate82inter4));
  nand2 gate678(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate679(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate680(.a(G7), .O(gate82inter7));
  inv1  gate681(.a(G326), .O(gate82inter8));
  nand2 gate682(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate683(.a(s_19), .b(gate82inter3), .O(gate82inter10));
  nor2  gate684(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate685(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate686(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1555(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1556(.a(gate86inter0), .b(s_144), .O(gate86inter1));
  and2  gate1557(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1558(.a(s_144), .O(gate86inter3));
  inv1  gate1559(.a(s_145), .O(gate86inter4));
  nand2 gate1560(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1561(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1562(.a(G8), .O(gate86inter7));
  inv1  gate1563(.a(G332), .O(gate86inter8));
  nand2 gate1564(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1565(.a(s_145), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1566(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1567(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1568(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2731(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2732(.a(gate88inter0), .b(s_312), .O(gate88inter1));
  and2  gate2733(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2734(.a(s_312), .O(gate88inter3));
  inv1  gate2735(.a(s_313), .O(gate88inter4));
  nand2 gate2736(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2737(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2738(.a(G16), .O(gate88inter7));
  inv1  gate2739(.a(G335), .O(gate88inter8));
  nand2 gate2740(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2741(.a(s_313), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2742(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2743(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2744(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2577(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2578(.a(gate94inter0), .b(s_290), .O(gate94inter1));
  and2  gate2579(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2580(.a(s_290), .O(gate94inter3));
  inv1  gate2581(.a(s_291), .O(gate94inter4));
  nand2 gate2582(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2583(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2584(.a(G22), .O(gate94inter7));
  inv1  gate2585(.a(G344), .O(gate94inter8));
  nand2 gate2586(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2587(.a(s_291), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2588(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2589(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2590(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1765(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1766(.a(gate99inter0), .b(s_174), .O(gate99inter1));
  and2  gate1767(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1768(.a(s_174), .O(gate99inter3));
  inv1  gate1769(.a(s_175), .O(gate99inter4));
  nand2 gate1770(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1771(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1772(.a(G27), .O(gate99inter7));
  inv1  gate1773(.a(G353), .O(gate99inter8));
  nand2 gate1774(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1775(.a(s_175), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1776(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1777(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1778(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1387(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1388(.a(gate101inter0), .b(s_120), .O(gate101inter1));
  and2  gate1389(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1390(.a(s_120), .O(gate101inter3));
  inv1  gate1391(.a(s_121), .O(gate101inter4));
  nand2 gate1392(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1393(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1394(.a(G20), .O(gate101inter7));
  inv1  gate1395(.a(G356), .O(gate101inter8));
  nand2 gate1396(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1397(.a(s_121), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1398(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1399(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1400(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1877(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1878(.a(gate102inter0), .b(s_190), .O(gate102inter1));
  and2  gate1879(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1880(.a(s_190), .O(gate102inter3));
  inv1  gate1881(.a(s_191), .O(gate102inter4));
  nand2 gate1882(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1883(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1884(.a(G24), .O(gate102inter7));
  inv1  gate1885(.a(G356), .O(gate102inter8));
  nand2 gate1886(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1887(.a(s_191), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1888(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1889(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1890(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate2493(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2494(.a(gate103inter0), .b(s_278), .O(gate103inter1));
  and2  gate2495(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2496(.a(s_278), .O(gate103inter3));
  inv1  gate2497(.a(s_279), .O(gate103inter4));
  nand2 gate2498(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2499(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2500(.a(G28), .O(gate103inter7));
  inv1  gate2501(.a(G359), .O(gate103inter8));
  nand2 gate2502(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2503(.a(s_279), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2504(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2505(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2506(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate561(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate562(.a(gate104inter0), .b(s_2), .O(gate104inter1));
  and2  gate563(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate564(.a(s_2), .O(gate104inter3));
  inv1  gate565(.a(s_3), .O(gate104inter4));
  nand2 gate566(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate567(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate568(.a(G32), .O(gate104inter7));
  inv1  gate569(.a(G359), .O(gate104inter8));
  nand2 gate570(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate571(.a(s_3), .b(gate104inter3), .O(gate104inter10));
  nor2  gate572(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate573(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate574(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate3123(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate3124(.a(gate105inter0), .b(s_368), .O(gate105inter1));
  and2  gate3125(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate3126(.a(s_368), .O(gate105inter3));
  inv1  gate3127(.a(s_369), .O(gate105inter4));
  nand2 gate3128(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate3129(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate3130(.a(G362), .O(gate105inter7));
  inv1  gate3131(.a(G363), .O(gate105inter8));
  nand2 gate3132(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate3133(.a(s_369), .b(gate105inter3), .O(gate105inter10));
  nor2  gate3134(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate3135(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate3136(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate2241(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2242(.a(gate106inter0), .b(s_242), .O(gate106inter1));
  and2  gate2243(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2244(.a(s_242), .O(gate106inter3));
  inv1  gate2245(.a(s_243), .O(gate106inter4));
  nand2 gate2246(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2247(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2248(.a(G364), .O(gate106inter7));
  inv1  gate2249(.a(G365), .O(gate106inter8));
  nand2 gate2250(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2251(.a(s_243), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2252(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2253(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2254(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate2997(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2998(.a(gate109inter0), .b(s_350), .O(gate109inter1));
  and2  gate2999(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate3000(.a(s_350), .O(gate109inter3));
  inv1  gate3001(.a(s_351), .O(gate109inter4));
  nand2 gate3002(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate3003(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate3004(.a(G370), .O(gate109inter7));
  inv1  gate3005(.a(G371), .O(gate109inter8));
  nand2 gate3006(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate3007(.a(s_351), .b(gate109inter3), .O(gate109inter10));
  nor2  gate3008(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate3009(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate3010(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate799(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate800(.a(gate110inter0), .b(s_36), .O(gate110inter1));
  and2  gate801(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate802(.a(s_36), .O(gate110inter3));
  inv1  gate803(.a(s_37), .O(gate110inter4));
  nand2 gate804(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate805(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate806(.a(G372), .O(gate110inter7));
  inv1  gate807(.a(G373), .O(gate110inter8));
  nand2 gate808(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate809(.a(s_37), .b(gate110inter3), .O(gate110inter10));
  nor2  gate810(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate811(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate812(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate827(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate828(.a(gate112inter0), .b(s_40), .O(gate112inter1));
  and2  gate829(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate830(.a(s_40), .O(gate112inter3));
  inv1  gate831(.a(s_41), .O(gate112inter4));
  nand2 gate832(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate833(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate834(.a(G376), .O(gate112inter7));
  inv1  gate835(.a(G377), .O(gate112inter8));
  nand2 gate836(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate837(.a(s_41), .b(gate112inter3), .O(gate112inter10));
  nor2  gate838(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate839(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate840(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2983(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2984(.a(gate115inter0), .b(s_348), .O(gate115inter1));
  and2  gate2985(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2986(.a(s_348), .O(gate115inter3));
  inv1  gate2987(.a(s_349), .O(gate115inter4));
  nand2 gate2988(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2989(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2990(.a(G382), .O(gate115inter7));
  inv1  gate2991(.a(G383), .O(gate115inter8));
  nand2 gate2992(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2993(.a(s_349), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2994(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2995(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2996(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate631(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate632(.a(gate116inter0), .b(s_12), .O(gate116inter1));
  and2  gate633(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate634(.a(s_12), .O(gate116inter3));
  inv1  gate635(.a(s_13), .O(gate116inter4));
  nand2 gate636(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate637(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate638(.a(G384), .O(gate116inter7));
  inv1  gate639(.a(G385), .O(gate116inter8));
  nand2 gate640(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate641(.a(s_13), .b(gate116inter3), .O(gate116inter10));
  nor2  gate642(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate643(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate644(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1793(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1794(.a(gate118inter0), .b(s_178), .O(gate118inter1));
  and2  gate1795(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1796(.a(s_178), .O(gate118inter3));
  inv1  gate1797(.a(s_179), .O(gate118inter4));
  nand2 gate1798(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1799(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1800(.a(G388), .O(gate118inter7));
  inv1  gate1801(.a(G389), .O(gate118inter8));
  nand2 gate1802(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1803(.a(s_179), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1804(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1805(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1806(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1191(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1192(.a(gate121inter0), .b(s_92), .O(gate121inter1));
  and2  gate1193(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1194(.a(s_92), .O(gate121inter3));
  inv1  gate1195(.a(s_93), .O(gate121inter4));
  nand2 gate1196(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1197(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1198(.a(G394), .O(gate121inter7));
  inv1  gate1199(.a(G395), .O(gate121inter8));
  nand2 gate1200(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1201(.a(s_93), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1202(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1203(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1204(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1849(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1850(.a(gate125inter0), .b(s_186), .O(gate125inter1));
  and2  gate1851(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1852(.a(s_186), .O(gate125inter3));
  inv1  gate1853(.a(s_187), .O(gate125inter4));
  nand2 gate1854(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1855(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1856(.a(G402), .O(gate125inter7));
  inv1  gate1857(.a(G403), .O(gate125inter8));
  nand2 gate1858(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1859(.a(s_187), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1860(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1861(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1862(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2507(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2508(.a(gate127inter0), .b(s_280), .O(gate127inter1));
  and2  gate2509(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2510(.a(s_280), .O(gate127inter3));
  inv1  gate2511(.a(s_281), .O(gate127inter4));
  nand2 gate2512(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2513(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2514(.a(G406), .O(gate127inter7));
  inv1  gate2515(.a(G407), .O(gate127inter8));
  nand2 gate2516(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2517(.a(s_281), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2518(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2519(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2520(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1429(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1430(.a(gate129inter0), .b(s_126), .O(gate129inter1));
  and2  gate1431(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1432(.a(s_126), .O(gate129inter3));
  inv1  gate1433(.a(s_127), .O(gate129inter4));
  nand2 gate1434(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1435(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1436(.a(G410), .O(gate129inter7));
  inv1  gate1437(.a(G411), .O(gate129inter8));
  nand2 gate1438(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1439(.a(s_127), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1440(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1441(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1442(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2899(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2900(.a(gate130inter0), .b(s_336), .O(gate130inter1));
  and2  gate2901(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2902(.a(s_336), .O(gate130inter3));
  inv1  gate2903(.a(s_337), .O(gate130inter4));
  nand2 gate2904(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2905(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2906(.a(G412), .O(gate130inter7));
  inv1  gate2907(.a(G413), .O(gate130inter8));
  nand2 gate2908(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2909(.a(s_337), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2910(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2911(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2912(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate603(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate604(.a(gate131inter0), .b(s_8), .O(gate131inter1));
  and2  gate605(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate606(.a(s_8), .O(gate131inter3));
  inv1  gate607(.a(s_9), .O(gate131inter4));
  nand2 gate608(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate609(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate610(.a(G414), .O(gate131inter7));
  inv1  gate611(.a(G415), .O(gate131inter8));
  nand2 gate612(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate613(.a(s_9), .b(gate131inter3), .O(gate131inter10));
  nor2  gate614(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate615(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate616(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate2521(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2522(.a(gate132inter0), .b(s_282), .O(gate132inter1));
  and2  gate2523(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2524(.a(s_282), .O(gate132inter3));
  inv1  gate2525(.a(s_283), .O(gate132inter4));
  nand2 gate2526(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2527(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2528(.a(G416), .O(gate132inter7));
  inv1  gate2529(.a(G417), .O(gate132inter8));
  nand2 gate2530(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2531(.a(s_283), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2532(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2533(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2534(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1513(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1514(.a(gate133inter0), .b(s_138), .O(gate133inter1));
  and2  gate1515(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1516(.a(s_138), .O(gate133inter3));
  inv1  gate1517(.a(s_139), .O(gate133inter4));
  nand2 gate1518(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1519(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1520(.a(G418), .O(gate133inter7));
  inv1  gate1521(.a(G419), .O(gate133inter8));
  nand2 gate1522(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1523(.a(s_139), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1524(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1525(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1526(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1359(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1360(.a(gate134inter0), .b(s_116), .O(gate134inter1));
  and2  gate1361(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1362(.a(s_116), .O(gate134inter3));
  inv1  gate1363(.a(s_117), .O(gate134inter4));
  nand2 gate1364(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1365(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1366(.a(G420), .O(gate134inter7));
  inv1  gate1367(.a(G421), .O(gate134inter8));
  nand2 gate1368(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1369(.a(s_117), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1370(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1371(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1372(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1709(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1710(.a(gate136inter0), .b(s_166), .O(gate136inter1));
  and2  gate1711(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1712(.a(s_166), .O(gate136inter3));
  inv1  gate1713(.a(s_167), .O(gate136inter4));
  nand2 gate1714(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1715(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1716(.a(G424), .O(gate136inter7));
  inv1  gate1717(.a(G425), .O(gate136inter8));
  nand2 gate1718(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1719(.a(s_167), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1720(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1721(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1722(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1695(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1696(.a(gate137inter0), .b(s_164), .O(gate137inter1));
  and2  gate1697(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1698(.a(s_164), .O(gate137inter3));
  inv1  gate1699(.a(s_165), .O(gate137inter4));
  nand2 gate1700(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1701(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1702(.a(G426), .O(gate137inter7));
  inv1  gate1703(.a(G429), .O(gate137inter8));
  nand2 gate1704(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1705(.a(s_165), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1706(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1707(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1708(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1149(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1150(.a(gate139inter0), .b(s_86), .O(gate139inter1));
  and2  gate1151(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1152(.a(s_86), .O(gate139inter3));
  inv1  gate1153(.a(s_87), .O(gate139inter4));
  nand2 gate1154(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1155(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1156(.a(G438), .O(gate139inter7));
  inv1  gate1157(.a(G441), .O(gate139inter8));
  nand2 gate1158(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1159(.a(s_87), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1160(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1161(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1162(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate3151(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate3152(.a(gate141inter0), .b(s_372), .O(gate141inter1));
  and2  gate3153(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate3154(.a(s_372), .O(gate141inter3));
  inv1  gate3155(.a(s_373), .O(gate141inter4));
  nand2 gate3156(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate3157(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate3158(.a(G450), .O(gate141inter7));
  inv1  gate3159(.a(G453), .O(gate141inter8));
  nand2 gate3160(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate3161(.a(s_373), .b(gate141inter3), .O(gate141inter10));
  nor2  gate3162(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate3163(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate3164(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate687(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate688(.a(gate142inter0), .b(s_20), .O(gate142inter1));
  and2  gate689(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate690(.a(s_20), .O(gate142inter3));
  inv1  gate691(.a(s_21), .O(gate142inter4));
  nand2 gate692(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate693(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate694(.a(G456), .O(gate142inter7));
  inv1  gate695(.a(G459), .O(gate142inter8));
  nand2 gate696(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate697(.a(s_21), .b(gate142inter3), .O(gate142inter10));
  nor2  gate698(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate699(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate700(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2451(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2452(.a(gate144inter0), .b(s_272), .O(gate144inter1));
  and2  gate2453(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2454(.a(s_272), .O(gate144inter3));
  inv1  gate2455(.a(s_273), .O(gate144inter4));
  nand2 gate2456(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2457(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2458(.a(G468), .O(gate144inter7));
  inv1  gate2459(.a(G471), .O(gate144inter8));
  nand2 gate2460(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2461(.a(s_273), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2462(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2463(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2464(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2927(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2928(.a(gate145inter0), .b(s_340), .O(gate145inter1));
  and2  gate2929(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2930(.a(s_340), .O(gate145inter3));
  inv1  gate2931(.a(s_341), .O(gate145inter4));
  nand2 gate2932(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2933(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2934(.a(G474), .O(gate145inter7));
  inv1  gate2935(.a(G477), .O(gate145inter8));
  nand2 gate2936(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2937(.a(s_341), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2938(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2939(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2940(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate953(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate954(.a(gate147inter0), .b(s_58), .O(gate147inter1));
  and2  gate955(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate956(.a(s_58), .O(gate147inter3));
  inv1  gate957(.a(s_59), .O(gate147inter4));
  nand2 gate958(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate959(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate960(.a(G486), .O(gate147inter7));
  inv1  gate961(.a(G489), .O(gate147inter8));
  nand2 gate962(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate963(.a(s_59), .b(gate147inter3), .O(gate147inter10));
  nor2  gate964(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate965(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate966(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2031(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2032(.a(gate149inter0), .b(s_212), .O(gate149inter1));
  and2  gate2033(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2034(.a(s_212), .O(gate149inter3));
  inv1  gate2035(.a(s_213), .O(gate149inter4));
  nand2 gate2036(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2037(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2038(.a(G498), .O(gate149inter7));
  inv1  gate2039(.a(G501), .O(gate149inter8));
  nand2 gate2040(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2041(.a(s_213), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2042(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2043(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2044(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1499(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1500(.a(gate150inter0), .b(s_136), .O(gate150inter1));
  and2  gate1501(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1502(.a(s_136), .O(gate150inter3));
  inv1  gate1503(.a(s_137), .O(gate150inter4));
  nand2 gate1504(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1505(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1506(.a(G504), .O(gate150inter7));
  inv1  gate1507(.a(G507), .O(gate150inter8));
  nand2 gate1508(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1509(.a(s_137), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1510(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1511(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1512(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate3277(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate3278(.a(gate151inter0), .b(s_390), .O(gate151inter1));
  and2  gate3279(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate3280(.a(s_390), .O(gate151inter3));
  inv1  gate3281(.a(s_391), .O(gate151inter4));
  nand2 gate3282(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate3283(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate3284(.a(G510), .O(gate151inter7));
  inv1  gate3285(.a(G513), .O(gate151inter8));
  nand2 gate3286(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate3287(.a(s_391), .b(gate151inter3), .O(gate151inter10));
  nor2  gate3288(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate3289(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate3290(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1093(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1094(.a(gate155inter0), .b(s_78), .O(gate155inter1));
  and2  gate1095(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1096(.a(s_78), .O(gate155inter3));
  inv1  gate1097(.a(s_79), .O(gate155inter4));
  nand2 gate1098(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1099(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1100(.a(G432), .O(gate155inter7));
  inv1  gate1101(.a(G525), .O(gate155inter8));
  nand2 gate1102(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1103(.a(s_79), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1104(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1105(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1106(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2829(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2830(.a(gate159inter0), .b(s_326), .O(gate159inter1));
  and2  gate2831(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2832(.a(s_326), .O(gate159inter3));
  inv1  gate2833(.a(s_327), .O(gate159inter4));
  nand2 gate2834(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2835(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2836(.a(G444), .O(gate159inter7));
  inv1  gate2837(.a(G531), .O(gate159inter8));
  nand2 gate2838(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2839(.a(s_327), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2840(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2841(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2842(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1569(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1570(.a(gate163inter0), .b(s_146), .O(gate163inter1));
  and2  gate1571(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1572(.a(s_146), .O(gate163inter3));
  inv1  gate1573(.a(s_147), .O(gate163inter4));
  nand2 gate1574(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1575(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1576(.a(G456), .O(gate163inter7));
  inv1  gate1577(.a(G537), .O(gate163inter8));
  nand2 gate1578(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1579(.a(s_147), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1580(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1581(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1582(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1289(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1290(.a(gate166inter0), .b(s_106), .O(gate166inter1));
  and2  gate1291(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1292(.a(s_106), .O(gate166inter3));
  inv1  gate1293(.a(s_107), .O(gate166inter4));
  nand2 gate1294(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1295(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1296(.a(G465), .O(gate166inter7));
  inv1  gate1297(.a(G540), .O(gate166inter8));
  nand2 gate1298(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1299(.a(s_107), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1300(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1301(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1302(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2843(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2844(.a(gate167inter0), .b(s_328), .O(gate167inter1));
  and2  gate2845(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2846(.a(s_328), .O(gate167inter3));
  inv1  gate2847(.a(s_329), .O(gate167inter4));
  nand2 gate2848(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2849(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2850(.a(G468), .O(gate167inter7));
  inv1  gate2851(.a(G543), .O(gate167inter8));
  nand2 gate2852(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2853(.a(s_329), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2854(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2855(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2856(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2409(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2410(.a(gate170inter0), .b(s_266), .O(gate170inter1));
  and2  gate2411(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2412(.a(s_266), .O(gate170inter3));
  inv1  gate2413(.a(s_267), .O(gate170inter4));
  nand2 gate2414(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2415(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2416(.a(G477), .O(gate170inter7));
  inv1  gate2417(.a(G546), .O(gate170inter8));
  nand2 gate2418(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2419(.a(s_267), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2420(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2421(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2422(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate855(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate856(.a(gate173inter0), .b(s_44), .O(gate173inter1));
  and2  gate857(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate858(.a(s_44), .O(gate173inter3));
  inv1  gate859(.a(s_45), .O(gate173inter4));
  nand2 gate860(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate861(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate862(.a(G486), .O(gate173inter7));
  inv1  gate863(.a(G552), .O(gate173inter8));
  nand2 gate864(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate865(.a(s_45), .b(gate173inter3), .O(gate173inter10));
  nor2  gate866(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate867(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate868(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate2171(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2172(.a(gate174inter0), .b(s_232), .O(gate174inter1));
  and2  gate2173(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2174(.a(s_232), .O(gate174inter3));
  inv1  gate2175(.a(s_233), .O(gate174inter4));
  nand2 gate2176(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2177(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2178(.a(G489), .O(gate174inter7));
  inv1  gate2179(.a(G552), .O(gate174inter8));
  nand2 gate2180(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2181(.a(s_233), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2182(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2183(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2184(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate2017(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2018(.a(gate175inter0), .b(s_210), .O(gate175inter1));
  and2  gate2019(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2020(.a(s_210), .O(gate175inter3));
  inv1  gate2021(.a(s_211), .O(gate175inter4));
  nand2 gate2022(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2023(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2024(.a(G492), .O(gate175inter7));
  inv1  gate2025(.a(G555), .O(gate175inter8));
  nand2 gate2026(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2027(.a(s_211), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2028(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2029(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2030(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate3025(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate3026(.a(gate176inter0), .b(s_354), .O(gate176inter1));
  and2  gate3027(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate3028(.a(s_354), .O(gate176inter3));
  inv1  gate3029(.a(s_355), .O(gate176inter4));
  nand2 gate3030(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate3031(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate3032(.a(G495), .O(gate176inter7));
  inv1  gate3033(.a(G555), .O(gate176inter8));
  nand2 gate3034(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate3035(.a(s_355), .b(gate176inter3), .O(gate176inter10));
  nor2  gate3036(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate3037(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate3038(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate1905(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1906(.a(gate177inter0), .b(s_194), .O(gate177inter1));
  and2  gate1907(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1908(.a(s_194), .O(gate177inter3));
  inv1  gate1909(.a(s_195), .O(gate177inter4));
  nand2 gate1910(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1911(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1912(.a(G498), .O(gate177inter7));
  inv1  gate1913(.a(G558), .O(gate177inter8));
  nand2 gate1914(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1915(.a(s_195), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1916(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1917(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1918(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate2003(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2004(.a(gate178inter0), .b(s_208), .O(gate178inter1));
  and2  gate2005(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2006(.a(s_208), .O(gate178inter3));
  inv1  gate2007(.a(s_209), .O(gate178inter4));
  nand2 gate2008(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2009(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2010(.a(G501), .O(gate178inter7));
  inv1  gate2011(.a(G558), .O(gate178inter8));
  nand2 gate2012(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2013(.a(s_209), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2014(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2015(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2016(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate3263(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate3264(.a(gate180inter0), .b(s_388), .O(gate180inter1));
  and2  gate3265(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate3266(.a(s_388), .O(gate180inter3));
  inv1  gate3267(.a(s_389), .O(gate180inter4));
  nand2 gate3268(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate3269(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate3270(.a(G507), .O(gate180inter7));
  inv1  gate3271(.a(G561), .O(gate180inter8));
  nand2 gate3272(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate3273(.a(s_389), .b(gate180inter3), .O(gate180inter10));
  nor2  gate3274(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate3275(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate3276(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1541(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1542(.a(gate183inter0), .b(s_142), .O(gate183inter1));
  and2  gate1543(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1544(.a(s_142), .O(gate183inter3));
  inv1  gate1545(.a(s_143), .O(gate183inter4));
  nand2 gate1546(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1547(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1548(.a(G516), .O(gate183inter7));
  inv1  gate1549(.a(G567), .O(gate183inter8));
  nand2 gate1550(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1551(.a(s_143), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1552(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1553(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1554(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2269(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2270(.a(gate185inter0), .b(s_246), .O(gate185inter1));
  and2  gate2271(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2272(.a(s_246), .O(gate185inter3));
  inv1  gate2273(.a(s_247), .O(gate185inter4));
  nand2 gate2274(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2275(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2276(.a(G570), .O(gate185inter7));
  inv1  gate2277(.a(G571), .O(gate185inter8));
  nand2 gate2278(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2279(.a(s_247), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2280(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2281(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2282(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1527(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1528(.a(gate188inter0), .b(s_140), .O(gate188inter1));
  and2  gate1529(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1530(.a(s_140), .O(gate188inter3));
  inv1  gate1531(.a(s_141), .O(gate188inter4));
  nand2 gate1532(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1533(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1534(.a(G576), .O(gate188inter7));
  inv1  gate1535(.a(G577), .O(gate188inter8));
  nand2 gate1536(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1537(.a(s_141), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1538(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1539(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1540(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate3137(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate3138(.a(gate190inter0), .b(s_370), .O(gate190inter1));
  and2  gate3139(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate3140(.a(s_370), .O(gate190inter3));
  inv1  gate3141(.a(s_371), .O(gate190inter4));
  nand2 gate3142(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate3143(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate3144(.a(G580), .O(gate190inter7));
  inv1  gate3145(.a(G581), .O(gate190inter8));
  nand2 gate3146(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate3147(.a(s_371), .b(gate190inter3), .O(gate190inter10));
  nor2  gate3148(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate3149(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate3150(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1779(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1780(.a(gate194inter0), .b(s_176), .O(gate194inter1));
  and2  gate1781(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1782(.a(s_176), .O(gate194inter3));
  inv1  gate1783(.a(s_177), .O(gate194inter4));
  nand2 gate1784(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1785(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1786(.a(G588), .O(gate194inter7));
  inv1  gate1787(.a(G589), .O(gate194inter8));
  nand2 gate1788(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1789(.a(s_177), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1790(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1791(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1792(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate925(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate926(.a(gate198inter0), .b(s_54), .O(gate198inter1));
  and2  gate927(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate928(.a(s_54), .O(gate198inter3));
  inv1  gate929(.a(s_55), .O(gate198inter4));
  nand2 gate930(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate931(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate932(.a(G596), .O(gate198inter7));
  inv1  gate933(.a(G597), .O(gate198inter8));
  nand2 gate934(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate935(.a(s_55), .b(gate198inter3), .O(gate198inter10));
  nor2  gate936(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate937(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate938(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1863(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1864(.a(gate199inter0), .b(s_188), .O(gate199inter1));
  and2  gate1865(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1866(.a(s_188), .O(gate199inter3));
  inv1  gate1867(.a(s_189), .O(gate199inter4));
  nand2 gate1868(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1869(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1870(.a(G598), .O(gate199inter7));
  inv1  gate1871(.a(G599), .O(gate199inter8));
  nand2 gate1872(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1873(.a(s_189), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1874(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1875(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1876(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2101(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2102(.a(gate204inter0), .b(s_222), .O(gate204inter1));
  and2  gate2103(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2104(.a(s_222), .O(gate204inter3));
  inv1  gate2105(.a(s_223), .O(gate204inter4));
  nand2 gate2106(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2107(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2108(.a(G607), .O(gate204inter7));
  inv1  gate2109(.a(G617), .O(gate204inter8));
  nand2 gate2110(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2111(.a(s_223), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2112(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2113(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2114(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1163(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1164(.a(gate205inter0), .b(s_88), .O(gate205inter1));
  and2  gate1165(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1166(.a(s_88), .O(gate205inter3));
  inv1  gate1167(.a(s_89), .O(gate205inter4));
  nand2 gate1168(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1169(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1170(.a(G622), .O(gate205inter7));
  inv1  gate1171(.a(G627), .O(gate205inter8));
  nand2 gate1172(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1173(.a(s_89), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1174(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1175(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1176(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1681(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1682(.a(gate206inter0), .b(s_162), .O(gate206inter1));
  and2  gate1683(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1684(.a(s_162), .O(gate206inter3));
  inv1  gate1685(.a(s_163), .O(gate206inter4));
  nand2 gate1686(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1687(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1688(.a(G632), .O(gate206inter7));
  inv1  gate1689(.a(G637), .O(gate206inter8));
  nand2 gate1690(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1691(.a(s_163), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1692(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1693(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1694(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2115(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2116(.a(gate208inter0), .b(s_224), .O(gate208inter1));
  and2  gate2117(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2118(.a(s_224), .O(gate208inter3));
  inv1  gate2119(.a(s_225), .O(gate208inter4));
  nand2 gate2120(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2121(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2122(.a(G627), .O(gate208inter7));
  inv1  gate2123(.a(G637), .O(gate208inter8));
  nand2 gate2124(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2125(.a(s_225), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2126(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2127(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2128(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1835(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1836(.a(gate209inter0), .b(s_184), .O(gate209inter1));
  and2  gate1837(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1838(.a(s_184), .O(gate209inter3));
  inv1  gate1839(.a(s_185), .O(gate209inter4));
  nand2 gate1840(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1841(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1842(.a(G602), .O(gate209inter7));
  inv1  gate1843(.a(G666), .O(gate209inter8));
  nand2 gate1844(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1845(.a(s_185), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1846(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1847(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1848(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1373(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1374(.a(gate213inter0), .b(s_118), .O(gate213inter1));
  and2  gate1375(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1376(.a(s_118), .O(gate213inter3));
  inv1  gate1377(.a(s_119), .O(gate213inter4));
  nand2 gate1378(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1379(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1380(.a(G602), .O(gate213inter7));
  inv1  gate1381(.a(G672), .O(gate213inter8));
  nand2 gate1382(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1383(.a(s_119), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1384(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1385(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1386(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1891(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1892(.a(gate216inter0), .b(s_192), .O(gate216inter1));
  and2  gate1893(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1894(.a(s_192), .O(gate216inter3));
  inv1  gate1895(.a(s_193), .O(gate216inter4));
  nand2 gate1896(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1897(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1898(.a(G617), .O(gate216inter7));
  inv1  gate1899(.a(G675), .O(gate216inter8));
  nand2 gate1900(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1901(.a(s_193), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1902(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1903(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1904(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2381(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2382(.a(gate218inter0), .b(s_262), .O(gate218inter1));
  and2  gate2383(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2384(.a(s_262), .O(gate218inter3));
  inv1  gate2385(.a(s_263), .O(gate218inter4));
  nand2 gate2386(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2387(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2388(.a(G627), .O(gate218inter7));
  inv1  gate2389(.a(G678), .O(gate218inter8));
  nand2 gate2390(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2391(.a(s_263), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2392(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2393(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2394(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1471(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1472(.a(gate219inter0), .b(s_132), .O(gate219inter1));
  and2  gate1473(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1474(.a(s_132), .O(gate219inter3));
  inv1  gate1475(.a(s_133), .O(gate219inter4));
  nand2 gate1476(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1477(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1478(.a(G632), .O(gate219inter7));
  inv1  gate1479(.a(G681), .O(gate219inter8));
  nand2 gate1480(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1481(.a(s_133), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1482(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1483(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1484(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate2059(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2060(.a(gate221inter0), .b(s_216), .O(gate221inter1));
  and2  gate2061(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2062(.a(s_216), .O(gate221inter3));
  inv1  gate2063(.a(s_217), .O(gate221inter4));
  nand2 gate2064(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2065(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2066(.a(G622), .O(gate221inter7));
  inv1  gate2067(.a(G684), .O(gate221inter8));
  nand2 gate2068(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2069(.a(s_217), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2070(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2071(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2072(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2143(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2144(.a(gate223inter0), .b(s_228), .O(gate223inter1));
  and2  gate2145(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2146(.a(s_228), .O(gate223inter3));
  inv1  gate2147(.a(s_229), .O(gate223inter4));
  nand2 gate2148(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2149(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2150(.a(G627), .O(gate223inter7));
  inv1  gate2151(.a(G687), .O(gate223inter8));
  nand2 gate2152(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2153(.a(s_229), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2154(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2155(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2156(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1597(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1598(.a(gate228inter0), .b(s_150), .O(gate228inter1));
  and2  gate1599(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1600(.a(s_150), .O(gate228inter3));
  inv1  gate1601(.a(s_151), .O(gate228inter4));
  nand2 gate1602(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1603(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1604(.a(G696), .O(gate228inter7));
  inv1  gate1605(.a(G697), .O(gate228inter8));
  nand2 gate1606(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1607(.a(s_151), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1608(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1609(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1610(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1667(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1668(.a(gate230inter0), .b(s_160), .O(gate230inter1));
  and2  gate1669(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1670(.a(s_160), .O(gate230inter3));
  inv1  gate1671(.a(s_161), .O(gate230inter4));
  nand2 gate1672(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1673(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1674(.a(G700), .O(gate230inter7));
  inv1  gate1675(.a(G701), .O(gate230inter8));
  nand2 gate1676(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1677(.a(s_161), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1678(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1679(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1680(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2885(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2886(.a(gate231inter0), .b(s_334), .O(gate231inter1));
  and2  gate2887(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2888(.a(s_334), .O(gate231inter3));
  inv1  gate2889(.a(s_335), .O(gate231inter4));
  nand2 gate2890(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2891(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2892(.a(G702), .O(gate231inter7));
  inv1  gate2893(.a(G703), .O(gate231inter8));
  nand2 gate2894(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2895(.a(s_335), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2896(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2897(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2898(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate2801(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2802(.a(gate235inter0), .b(s_322), .O(gate235inter1));
  and2  gate2803(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2804(.a(s_322), .O(gate235inter3));
  inv1  gate2805(.a(s_323), .O(gate235inter4));
  nand2 gate2806(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2807(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2808(.a(G248), .O(gate235inter7));
  inv1  gate2809(.a(G724), .O(gate235inter8));
  nand2 gate2810(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2811(.a(s_323), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2812(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2813(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2814(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate1177(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1178(.a(gate236inter0), .b(s_90), .O(gate236inter1));
  and2  gate1179(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1180(.a(s_90), .O(gate236inter3));
  inv1  gate1181(.a(s_91), .O(gate236inter4));
  nand2 gate1182(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1183(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1184(.a(G251), .O(gate236inter7));
  inv1  gate1185(.a(G727), .O(gate236inter8));
  nand2 gate1186(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1187(.a(s_91), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1188(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1189(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1190(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate645(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate646(.a(gate239inter0), .b(s_14), .O(gate239inter1));
  and2  gate647(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate648(.a(s_14), .O(gate239inter3));
  inv1  gate649(.a(s_15), .O(gate239inter4));
  nand2 gate650(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate651(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate652(.a(G260), .O(gate239inter7));
  inv1  gate653(.a(G712), .O(gate239inter8));
  nand2 gate654(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate655(.a(s_15), .b(gate239inter3), .O(gate239inter10));
  nor2  gate656(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate657(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate658(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2479(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2480(.a(gate244inter0), .b(s_276), .O(gate244inter1));
  and2  gate2481(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2482(.a(s_276), .O(gate244inter3));
  inv1  gate2483(.a(s_277), .O(gate244inter4));
  nand2 gate2484(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2485(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2486(.a(G721), .O(gate244inter7));
  inv1  gate2487(.a(G733), .O(gate244inter8));
  nand2 gate2488(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2489(.a(s_277), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2490(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2491(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2492(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1401(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1402(.a(gate245inter0), .b(s_122), .O(gate245inter1));
  and2  gate1403(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1404(.a(s_122), .O(gate245inter3));
  inv1  gate1405(.a(s_123), .O(gate245inter4));
  nand2 gate1406(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1407(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1408(.a(G248), .O(gate245inter7));
  inv1  gate1409(.a(G736), .O(gate245inter8));
  nand2 gate1410(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1411(.a(s_123), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1412(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1413(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1414(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1233(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1234(.a(gate250inter0), .b(s_98), .O(gate250inter1));
  and2  gate1235(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1236(.a(s_98), .O(gate250inter3));
  inv1  gate1237(.a(s_99), .O(gate250inter4));
  nand2 gate1238(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1239(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1240(.a(G706), .O(gate250inter7));
  inv1  gate1241(.a(G742), .O(gate250inter8));
  nand2 gate1242(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1243(.a(s_99), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1244(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1245(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1246(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1611(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1612(.a(gate251inter0), .b(s_152), .O(gate251inter1));
  and2  gate1613(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1614(.a(s_152), .O(gate251inter3));
  inv1  gate1615(.a(s_153), .O(gate251inter4));
  nand2 gate1616(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1617(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1618(.a(G257), .O(gate251inter7));
  inv1  gate1619(.a(G745), .O(gate251inter8));
  nand2 gate1620(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1621(.a(s_153), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1622(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1623(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1624(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1205(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1206(.a(gate257inter0), .b(s_94), .O(gate257inter1));
  and2  gate1207(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1208(.a(s_94), .O(gate257inter3));
  inv1  gate1209(.a(s_95), .O(gate257inter4));
  nand2 gate1210(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1211(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1212(.a(G754), .O(gate257inter7));
  inv1  gate1213(.a(G755), .O(gate257inter8));
  nand2 gate1214(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1215(.a(s_95), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1216(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1217(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1218(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate813(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate814(.a(gate258inter0), .b(s_38), .O(gate258inter1));
  and2  gate815(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate816(.a(s_38), .O(gate258inter3));
  inv1  gate817(.a(s_39), .O(gate258inter4));
  nand2 gate818(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate819(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate820(.a(G756), .O(gate258inter7));
  inv1  gate821(.a(G757), .O(gate258inter8));
  nand2 gate822(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate823(.a(s_39), .b(gate258inter3), .O(gate258inter10));
  nor2  gate824(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate825(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate826(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2339(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2340(.a(gate262inter0), .b(s_256), .O(gate262inter1));
  and2  gate2341(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2342(.a(s_256), .O(gate262inter3));
  inv1  gate2343(.a(s_257), .O(gate262inter4));
  nand2 gate2344(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2345(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2346(.a(G764), .O(gate262inter7));
  inv1  gate2347(.a(G765), .O(gate262inter8));
  nand2 gate2348(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2349(.a(s_257), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2350(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2351(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2352(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate911(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate912(.a(gate264inter0), .b(s_52), .O(gate264inter1));
  and2  gate913(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate914(.a(s_52), .O(gate264inter3));
  inv1  gate915(.a(s_53), .O(gate264inter4));
  nand2 gate916(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate917(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate918(.a(G768), .O(gate264inter7));
  inv1  gate919(.a(G769), .O(gate264inter8));
  nand2 gate920(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate921(.a(s_53), .b(gate264inter3), .O(gate264inter10));
  nor2  gate922(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate923(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate924(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate2367(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2368(.a(gate266inter0), .b(s_260), .O(gate266inter1));
  and2  gate2369(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2370(.a(s_260), .O(gate266inter3));
  inv1  gate2371(.a(s_261), .O(gate266inter4));
  nand2 gate2372(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2373(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2374(.a(G645), .O(gate266inter7));
  inv1  gate2375(.a(G773), .O(gate266inter8));
  nand2 gate2376(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2377(.a(s_261), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2378(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2379(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2380(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2465(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2466(.a(gate270inter0), .b(s_274), .O(gate270inter1));
  and2  gate2467(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2468(.a(s_274), .O(gate270inter3));
  inv1  gate2469(.a(s_275), .O(gate270inter4));
  nand2 gate2470(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2471(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2472(.a(G657), .O(gate270inter7));
  inv1  gate2473(.a(G785), .O(gate270inter8));
  nand2 gate2474(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2475(.a(s_275), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2476(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2477(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2478(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1345(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1346(.a(gate271inter0), .b(s_114), .O(gate271inter1));
  and2  gate1347(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1348(.a(s_114), .O(gate271inter3));
  inv1  gate1349(.a(s_115), .O(gate271inter4));
  nand2 gate1350(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1351(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1352(.a(G660), .O(gate271inter7));
  inv1  gate1353(.a(G788), .O(gate271inter8));
  nand2 gate1354(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1355(.a(s_115), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1356(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1357(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1358(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2283(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2284(.a(gate272inter0), .b(s_248), .O(gate272inter1));
  and2  gate2285(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2286(.a(s_248), .O(gate272inter3));
  inv1  gate2287(.a(s_249), .O(gate272inter4));
  nand2 gate2288(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2289(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2290(.a(G663), .O(gate272inter7));
  inv1  gate2291(.a(G791), .O(gate272inter8));
  nand2 gate2292(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2293(.a(s_249), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2294(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2295(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2296(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1009(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1010(.a(gate276inter0), .b(s_66), .O(gate276inter1));
  and2  gate1011(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1012(.a(s_66), .O(gate276inter3));
  inv1  gate1013(.a(s_67), .O(gate276inter4));
  nand2 gate1014(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1015(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1016(.a(G773), .O(gate276inter7));
  inv1  gate1017(.a(G797), .O(gate276inter8));
  nand2 gate1018(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1019(.a(s_67), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1020(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1021(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1022(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate2535(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2536(.a(gate277inter0), .b(s_284), .O(gate277inter1));
  and2  gate2537(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2538(.a(s_284), .O(gate277inter3));
  inv1  gate2539(.a(s_285), .O(gate277inter4));
  nand2 gate2540(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2541(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2542(.a(G648), .O(gate277inter7));
  inv1  gate2543(.a(G800), .O(gate277inter8));
  nand2 gate2544(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2545(.a(s_285), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2546(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2547(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2548(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2717(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2718(.a(gate281inter0), .b(s_310), .O(gate281inter1));
  and2  gate2719(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2720(.a(s_310), .O(gate281inter3));
  inv1  gate2721(.a(s_311), .O(gate281inter4));
  nand2 gate2722(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2723(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2724(.a(G654), .O(gate281inter7));
  inv1  gate2725(.a(G806), .O(gate281inter8));
  nand2 gate2726(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2727(.a(s_311), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2728(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2729(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2730(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2185(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2186(.a(gate282inter0), .b(s_234), .O(gate282inter1));
  and2  gate2187(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2188(.a(s_234), .O(gate282inter3));
  inv1  gate2189(.a(s_235), .O(gate282inter4));
  nand2 gate2190(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2191(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2192(.a(G782), .O(gate282inter7));
  inv1  gate2193(.a(G806), .O(gate282inter8));
  nand2 gate2194(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2195(.a(s_235), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2196(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2197(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2198(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1975(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1976(.a(gate284inter0), .b(s_204), .O(gate284inter1));
  and2  gate1977(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1978(.a(s_204), .O(gate284inter3));
  inv1  gate1979(.a(s_205), .O(gate284inter4));
  nand2 gate1980(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1981(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1982(.a(G785), .O(gate284inter7));
  inv1  gate1983(.a(G809), .O(gate284inter8));
  nand2 gate1984(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1985(.a(s_205), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1986(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1987(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1988(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1485(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1486(.a(gate285inter0), .b(s_134), .O(gate285inter1));
  and2  gate1487(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1488(.a(s_134), .O(gate285inter3));
  inv1  gate1489(.a(s_135), .O(gate285inter4));
  nand2 gate1490(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1491(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1492(.a(G660), .O(gate285inter7));
  inv1  gate1493(.a(G812), .O(gate285inter8));
  nand2 gate1494(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1495(.a(s_135), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1496(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1497(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1498(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1751(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1752(.a(gate287inter0), .b(s_172), .O(gate287inter1));
  and2  gate1753(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1754(.a(s_172), .O(gate287inter3));
  inv1  gate1755(.a(s_173), .O(gate287inter4));
  nand2 gate1756(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1757(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1758(.a(G663), .O(gate287inter7));
  inv1  gate1759(.a(G815), .O(gate287inter8));
  nand2 gate1760(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1761(.a(s_173), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1762(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1763(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1764(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2227(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2228(.a(gate292inter0), .b(s_240), .O(gate292inter1));
  and2  gate2229(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2230(.a(s_240), .O(gate292inter3));
  inv1  gate2231(.a(s_241), .O(gate292inter4));
  nand2 gate2232(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2233(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2234(.a(G824), .O(gate292inter7));
  inv1  gate2235(.a(G825), .O(gate292inter8));
  nand2 gate2236(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2237(.a(s_241), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2238(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2239(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2240(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2703(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2704(.a(gate295inter0), .b(s_308), .O(gate295inter1));
  and2  gate2705(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2706(.a(s_308), .O(gate295inter3));
  inv1  gate2707(.a(s_309), .O(gate295inter4));
  nand2 gate2708(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2709(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2710(.a(G830), .O(gate295inter7));
  inv1  gate2711(.a(G831), .O(gate295inter8));
  nand2 gate2712(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2713(.a(s_309), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2714(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2715(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2716(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1317(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1318(.a(gate296inter0), .b(s_110), .O(gate296inter1));
  and2  gate1319(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1320(.a(s_110), .O(gate296inter3));
  inv1  gate1321(.a(s_111), .O(gate296inter4));
  nand2 gate1322(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1323(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1324(.a(G826), .O(gate296inter7));
  inv1  gate1325(.a(G827), .O(gate296inter8));
  nand2 gate1326(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1327(.a(s_111), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1328(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1329(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1330(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate3095(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate3096(.a(gate389inter0), .b(s_364), .O(gate389inter1));
  and2  gate3097(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate3098(.a(s_364), .O(gate389inter3));
  inv1  gate3099(.a(s_365), .O(gate389inter4));
  nand2 gate3100(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate3101(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate3102(.a(G3), .O(gate389inter7));
  inv1  gate3103(.a(G1042), .O(gate389inter8));
  nand2 gate3104(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate3105(.a(s_365), .b(gate389inter3), .O(gate389inter10));
  nor2  gate3106(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate3107(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate3108(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1415(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1416(.a(gate391inter0), .b(s_124), .O(gate391inter1));
  and2  gate1417(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1418(.a(s_124), .O(gate391inter3));
  inv1  gate1419(.a(s_125), .O(gate391inter4));
  nand2 gate1420(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1421(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1422(.a(G5), .O(gate391inter7));
  inv1  gate1423(.a(G1048), .O(gate391inter8));
  nand2 gate1424(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1425(.a(s_125), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1426(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1427(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1428(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate2633(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2634(.a(gate392inter0), .b(s_298), .O(gate392inter1));
  and2  gate2635(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2636(.a(s_298), .O(gate392inter3));
  inv1  gate2637(.a(s_299), .O(gate392inter4));
  nand2 gate2638(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2639(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2640(.a(G6), .O(gate392inter7));
  inv1  gate2641(.a(G1051), .O(gate392inter8));
  nand2 gate2642(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2643(.a(s_299), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2644(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2645(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2646(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate967(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate968(.a(gate395inter0), .b(s_60), .O(gate395inter1));
  and2  gate969(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate970(.a(s_60), .O(gate395inter3));
  inv1  gate971(.a(s_61), .O(gate395inter4));
  nand2 gate972(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate973(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate974(.a(G9), .O(gate395inter7));
  inv1  gate975(.a(G1060), .O(gate395inter8));
  nand2 gate976(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate977(.a(s_61), .b(gate395inter3), .O(gate395inter10));
  nor2  gate978(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate979(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate980(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate2073(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2074(.a(gate399inter0), .b(s_218), .O(gate399inter1));
  and2  gate2075(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2076(.a(s_218), .O(gate399inter3));
  inv1  gate2077(.a(s_219), .O(gate399inter4));
  nand2 gate2078(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2079(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2080(.a(G13), .O(gate399inter7));
  inv1  gate2081(.a(G1072), .O(gate399inter8));
  nand2 gate2082(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2083(.a(s_219), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2084(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2085(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2086(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2759(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2760(.a(gate400inter0), .b(s_316), .O(gate400inter1));
  and2  gate2761(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2762(.a(s_316), .O(gate400inter3));
  inv1  gate2763(.a(s_317), .O(gate400inter4));
  nand2 gate2764(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2765(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2766(.a(G14), .O(gate400inter7));
  inv1  gate2767(.a(G1075), .O(gate400inter8));
  nand2 gate2768(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2769(.a(s_317), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2770(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2771(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2772(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate869(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate870(.a(gate403inter0), .b(s_46), .O(gate403inter1));
  and2  gate871(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate872(.a(s_46), .O(gate403inter3));
  inv1  gate873(.a(s_47), .O(gate403inter4));
  nand2 gate874(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate875(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate876(.a(G17), .O(gate403inter7));
  inv1  gate877(.a(G1084), .O(gate403inter8));
  nand2 gate878(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate879(.a(s_47), .b(gate403inter3), .O(gate403inter10));
  nor2  gate880(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate881(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate882(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1639(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1640(.a(gate404inter0), .b(s_156), .O(gate404inter1));
  and2  gate1641(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1642(.a(s_156), .O(gate404inter3));
  inv1  gate1643(.a(s_157), .O(gate404inter4));
  nand2 gate1644(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1645(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1646(.a(G18), .O(gate404inter7));
  inv1  gate1647(.a(G1087), .O(gate404inter8));
  nand2 gate1648(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1649(.a(s_157), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1650(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1651(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1652(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate617(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate618(.a(gate407inter0), .b(s_10), .O(gate407inter1));
  and2  gate619(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate620(.a(s_10), .O(gate407inter3));
  inv1  gate621(.a(s_11), .O(gate407inter4));
  nand2 gate622(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate623(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate624(.a(G21), .O(gate407inter7));
  inv1  gate625(.a(G1096), .O(gate407inter8));
  nand2 gate626(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate627(.a(s_11), .b(gate407inter3), .O(gate407inter10));
  nor2  gate628(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate629(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate630(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2941(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2942(.a(gate409inter0), .b(s_342), .O(gate409inter1));
  and2  gate2943(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2944(.a(s_342), .O(gate409inter3));
  inv1  gate2945(.a(s_343), .O(gate409inter4));
  nand2 gate2946(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2947(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2948(.a(G23), .O(gate409inter7));
  inv1  gate2949(.a(G1102), .O(gate409inter8));
  nand2 gate2950(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2951(.a(s_343), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2952(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2953(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2954(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2395(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2396(.a(gate410inter0), .b(s_264), .O(gate410inter1));
  and2  gate2397(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2398(.a(s_264), .O(gate410inter3));
  inv1  gate2399(.a(s_265), .O(gate410inter4));
  nand2 gate2400(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2401(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2402(.a(G24), .O(gate410inter7));
  inv1  gate2403(.a(G1105), .O(gate410inter8));
  nand2 gate2404(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2405(.a(s_265), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2406(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2407(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2408(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate3011(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate3012(.a(gate412inter0), .b(s_352), .O(gate412inter1));
  and2  gate3013(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate3014(.a(s_352), .O(gate412inter3));
  inv1  gate3015(.a(s_353), .O(gate412inter4));
  nand2 gate3016(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate3017(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate3018(.a(G26), .O(gate412inter7));
  inv1  gate3019(.a(G1111), .O(gate412inter8));
  nand2 gate3020(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate3021(.a(s_353), .b(gate412inter3), .O(gate412inter10));
  nor2  gate3022(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate3023(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate3024(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1653(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1654(.a(gate413inter0), .b(s_158), .O(gate413inter1));
  and2  gate1655(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1656(.a(s_158), .O(gate413inter3));
  inv1  gate1657(.a(s_159), .O(gate413inter4));
  nand2 gate1658(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1659(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1660(.a(G27), .O(gate413inter7));
  inv1  gate1661(.a(G1114), .O(gate413inter8));
  nand2 gate1662(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1663(.a(s_159), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1664(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1665(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1666(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2199(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2200(.a(gate414inter0), .b(s_236), .O(gate414inter1));
  and2  gate2201(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2202(.a(s_236), .O(gate414inter3));
  inv1  gate2203(.a(s_237), .O(gate414inter4));
  nand2 gate2204(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2205(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2206(.a(G28), .O(gate414inter7));
  inv1  gate2207(.a(G1117), .O(gate414inter8));
  nand2 gate2208(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2209(.a(s_237), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2210(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2211(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2212(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate2857(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2858(.a(gate415inter0), .b(s_330), .O(gate415inter1));
  and2  gate2859(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2860(.a(s_330), .O(gate415inter3));
  inv1  gate2861(.a(s_331), .O(gate415inter4));
  nand2 gate2862(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2863(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2864(.a(G29), .O(gate415inter7));
  inv1  gate2865(.a(G1120), .O(gate415inter8));
  nand2 gate2866(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2867(.a(s_331), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2868(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2869(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2870(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1331(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1332(.a(gate416inter0), .b(s_112), .O(gate416inter1));
  and2  gate1333(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1334(.a(s_112), .O(gate416inter3));
  inv1  gate1335(.a(s_113), .O(gate416inter4));
  nand2 gate1336(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1337(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1338(.a(G30), .O(gate416inter7));
  inv1  gate1339(.a(G1123), .O(gate416inter8));
  nand2 gate1340(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1341(.a(s_113), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1342(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1343(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1344(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate883(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate884(.a(gate417inter0), .b(s_48), .O(gate417inter1));
  and2  gate885(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate886(.a(s_48), .O(gate417inter3));
  inv1  gate887(.a(s_49), .O(gate417inter4));
  nand2 gate888(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate889(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate890(.a(G31), .O(gate417inter7));
  inv1  gate891(.a(G1126), .O(gate417inter8));
  nand2 gate892(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate893(.a(s_49), .b(gate417inter3), .O(gate417inter10));
  nor2  gate894(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate895(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate896(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2255(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2256(.a(gate418inter0), .b(s_244), .O(gate418inter1));
  and2  gate2257(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2258(.a(s_244), .O(gate418inter3));
  inv1  gate2259(.a(s_245), .O(gate418inter4));
  nand2 gate2260(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2261(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2262(.a(G32), .O(gate418inter7));
  inv1  gate2263(.a(G1129), .O(gate418inter8));
  nand2 gate2264(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2265(.a(s_245), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2266(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2267(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2268(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2353(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2354(.a(gate419inter0), .b(s_258), .O(gate419inter1));
  and2  gate2355(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2356(.a(s_258), .O(gate419inter3));
  inv1  gate2357(.a(s_259), .O(gate419inter4));
  nand2 gate2358(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2359(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2360(.a(G1), .O(gate419inter7));
  inv1  gate2361(.a(G1132), .O(gate419inter8));
  nand2 gate2362(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2363(.a(s_259), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2364(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2365(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2366(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1807(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1808(.a(gate420inter0), .b(s_180), .O(gate420inter1));
  and2  gate1809(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1810(.a(s_180), .O(gate420inter3));
  inv1  gate1811(.a(s_181), .O(gate420inter4));
  nand2 gate1812(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1813(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1814(.a(G1036), .O(gate420inter7));
  inv1  gate1815(.a(G1132), .O(gate420inter8));
  nand2 gate1816(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1817(.a(s_181), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1818(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1819(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1820(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1079(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1080(.a(gate423inter0), .b(s_76), .O(gate423inter1));
  and2  gate1081(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1082(.a(s_76), .O(gate423inter3));
  inv1  gate1083(.a(s_77), .O(gate423inter4));
  nand2 gate1084(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1085(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1086(.a(G3), .O(gate423inter7));
  inv1  gate1087(.a(G1138), .O(gate423inter8));
  nand2 gate1088(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1089(.a(s_77), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1090(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1091(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1092(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate715(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate716(.a(gate425inter0), .b(s_24), .O(gate425inter1));
  and2  gate717(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate718(.a(s_24), .O(gate425inter3));
  inv1  gate719(.a(s_25), .O(gate425inter4));
  nand2 gate720(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate721(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate722(.a(G4), .O(gate425inter7));
  inv1  gate723(.a(G1141), .O(gate425inter8));
  nand2 gate724(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate725(.a(s_25), .b(gate425inter3), .O(gate425inter10));
  nor2  gate726(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate727(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate728(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1219(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1220(.a(gate426inter0), .b(s_96), .O(gate426inter1));
  and2  gate1221(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1222(.a(s_96), .O(gate426inter3));
  inv1  gate1223(.a(s_97), .O(gate426inter4));
  nand2 gate1224(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1225(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1226(.a(G1045), .O(gate426inter7));
  inv1  gate1227(.a(G1141), .O(gate426inter8));
  nand2 gate1228(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1229(.a(s_97), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1230(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1231(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1232(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate3109(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate3110(.a(gate428inter0), .b(s_366), .O(gate428inter1));
  and2  gate3111(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate3112(.a(s_366), .O(gate428inter3));
  inv1  gate3113(.a(s_367), .O(gate428inter4));
  nand2 gate3114(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate3115(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate3116(.a(G1048), .O(gate428inter7));
  inv1  gate3117(.a(G1144), .O(gate428inter8));
  nand2 gate3118(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate3119(.a(s_367), .b(gate428inter3), .O(gate428inter10));
  nor2  gate3120(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate3121(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate3122(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1261(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1262(.a(gate429inter0), .b(s_102), .O(gate429inter1));
  and2  gate1263(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1264(.a(s_102), .O(gate429inter3));
  inv1  gate1265(.a(s_103), .O(gate429inter4));
  nand2 gate1266(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1267(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1268(.a(G6), .O(gate429inter7));
  inv1  gate1269(.a(G1147), .O(gate429inter8));
  nand2 gate1270(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1271(.a(s_103), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1272(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1273(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1274(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate3039(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate3040(.a(gate432inter0), .b(s_356), .O(gate432inter1));
  and2  gate3041(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate3042(.a(s_356), .O(gate432inter3));
  inv1  gate3043(.a(s_357), .O(gate432inter4));
  nand2 gate3044(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate3045(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate3046(.a(G1054), .O(gate432inter7));
  inv1  gate3047(.a(G1150), .O(gate432inter8));
  nand2 gate3048(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate3049(.a(s_357), .b(gate432inter3), .O(gate432inter10));
  nor2  gate3050(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate3051(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate3052(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1443(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1444(.a(gate433inter0), .b(s_128), .O(gate433inter1));
  and2  gate1445(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1446(.a(s_128), .O(gate433inter3));
  inv1  gate1447(.a(s_129), .O(gate433inter4));
  nand2 gate1448(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1449(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1450(.a(G8), .O(gate433inter7));
  inv1  gate1451(.a(G1153), .O(gate433inter8));
  nand2 gate1452(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1453(.a(s_129), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1454(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1455(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1456(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate743(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate744(.a(gate434inter0), .b(s_28), .O(gate434inter1));
  and2  gate745(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate746(.a(s_28), .O(gate434inter3));
  inv1  gate747(.a(s_29), .O(gate434inter4));
  nand2 gate748(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate749(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate750(.a(G1057), .O(gate434inter7));
  inv1  gate751(.a(G1153), .O(gate434inter8));
  nand2 gate752(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate753(.a(s_29), .b(gate434inter3), .O(gate434inter10));
  nor2  gate754(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate755(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate756(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2045(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2046(.a(gate435inter0), .b(s_214), .O(gate435inter1));
  and2  gate2047(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2048(.a(s_214), .O(gate435inter3));
  inv1  gate2049(.a(s_215), .O(gate435inter4));
  nand2 gate2050(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2051(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2052(.a(G9), .O(gate435inter7));
  inv1  gate2053(.a(G1156), .O(gate435inter8));
  nand2 gate2054(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2055(.a(s_215), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2056(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2057(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2058(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate3221(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate3222(.a(gate437inter0), .b(s_382), .O(gate437inter1));
  and2  gate3223(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate3224(.a(s_382), .O(gate437inter3));
  inv1  gate3225(.a(s_383), .O(gate437inter4));
  nand2 gate3226(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate3227(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate3228(.a(G10), .O(gate437inter7));
  inv1  gate3229(.a(G1159), .O(gate437inter8));
  nand2 gate3230(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate3231(.a(s_383), .b(gate437inter3), .O(gate437inter10));
  nor2  gate3232(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate3233(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate3234(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1303(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1304(.a(gate438inter0), .b(s_108), .O(gate438inter1));
  and2  gate1305(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1306(.a(s_108), .O(gate438inter3));
  inv1  gate1307(.a(s_109), .O(gate438inter4));
  nand2 gate1308(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1309(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1310(.a(G1063), .O(gate438inter7));
  inv1  gate1311(.a(G1159), .O(gate438inter8));
  nand2 gate1312(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1313(.a(s_109), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1314(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1315(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1316(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate3067(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate3068(.a(gate439inter0), .b(s_360), .O(gate439inter1));
  and2  gate3069(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate3070(.a(s_360), .O(gate439inter3));
  inv1  gate3071(.a(s_361), .O(gate439inter4));
  nand2 gate3072(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate3073(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate3074(.a(G11), .O(gate439inter7));
  inv1  gate3075(.a(G1162), .O(gate439inter8));
  nand2 gate3076(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate3077(.a(s_361), .b(gate439inter3), .O(gate439inter10));
  nor2  gate3078(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate3079(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate3080(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1947(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1948(.a(gate441inter0), .b(s_200), .O(gate441inter1));
  and2  gate1949(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1950(.a(s_200), .O(gate441inter3));
  inv1  gate1951(.a(s_201), .O(gate441inter4));
  nand2 gate1952(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1953(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1954(.a(G12), .O(gate441inter7));
  inv1  gate1955(.a(G1165), .O(gate441inter8));
  nand2 gate1956(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1957(.a(s_201), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1958(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1959(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1960(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1933(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1934(.a(gate442inter0), .b(s_198), .O(gate442inter1));
  and2  gate1935(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1936(.a(s_198), .O(gate442inter3));
  inv1  gate1937(.a(s_199), .O(gate442inter4));
  nand2 gate1938(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1939(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1940(.a(G1069), .O(gate442inter7));
  inv1  gate1941(.a(G1165), .O(gate442inter8));
  nand2 gate1942(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1943(.a(s_199), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1944(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1945(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1946(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2297(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2298(.a(gate444inter0), .b(s_250), .O(gate444inter1));
  and2  gate2299(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2300(.a(s_250), .O(gate444inter3));
  inv1  gate2301(.a(s_251), .O(gate444inter4));
  nand2 gate2302(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2303(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2304(.a(G1072), .O(gate444inter7));
  inv1  gate2305(.a(G1168), .O(gate444inter8));
  nand2 gate2306(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2307(.a(s_251), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2308(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2309(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2310(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1275(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1276(.a(gate446inter0), .b(s_104), .O(gate446inter1));
  and2  gate1277(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1278(.a(s_104), .O(gate446inter3));
  inv1  gate1279(.a(s_105), .O(gate446inter4));
  nand2 gate1280(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1281(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1282(.a(G1075), .O(gate446inter7));
  inv1  gate1283(.a(G1171), .O(gate446inter8));
  nand2 gate1284(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1285(.a(s_105), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1286(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1287(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1288(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1457(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1458(.a(gate451inter0), .b(s_130), .O(gate451inter1));
  and2  gate1459(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1460(.a(s_130), .O(gate451inter3));
  inv1  gate1461(.a(s_131), .O(gate451inter4));
  nand2 gate1462(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1463(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1464(.a(G17), .O(gate451inter7));
  inv1  gate1465(.a(G1180), .O(gate451inter8));
  nand2 gate1466(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1467(.a(s_131), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1468(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1469(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1470(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate575(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate576(.a(gate452inter0), .b(s_4), .O(gate452inter1));
  and2  gate577(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate578(.a(s_4), .O(gate452inter3));
  inv1  gate579(.a(s_5), .O(gate452inter4));
  nand2 gate580(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate581(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate582(.a(G1084), .O(gate452inter7));
  inv1  gate583(.a(G1180), .O(gate452inter8));
  nand2 gate584(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate585(.a(s_5), .b(gate452inter3), .O(gate452inter10));
  nor2  gate586(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate587(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate588(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate547(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate548(.a(gate453inter0), .b(s_0), .O(gate453inter1));
  and2  gate549(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate550(.a(s_0), .O(gate453inter3));
  inv1  gate551(.a(s_1), .O(gate453inter4));
  nand2 gate552(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate553(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate554(.a(G18), .O(gate453inter7));
  inv1  gate555(.a(G1183), .O(gate453inter8));
  nand2 gate556(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate557(.a(s_1), .b(gate453inter3), .O(gate453inter10));
  nor2  gate558(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate559(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate560(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2815(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2816(.a(gate456inter0), .b(s_324), .O(gate456inter1));
  and2  gate2817(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2818(.a(s_324), .O(gate456inter3));
  inv1  gate2819(.a(s_325), .O(gate456inter4));
  nand2 gate2820(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2821(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2822(.a(G1090), .O(gate456inter7));
  inv1  gate2823(.a(G1186), .O(gate456inter8));
  nand2 gate2824(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2825(.a(s_325), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2826(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2827(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2828(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate785(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate786(.a(gate457inter0), .b(s_34), .O(gate457inter1));
  and2  gate787(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate788(.a(s_34), .O(gate457inter3));
  inv1  gate789(.a(s_35), .O(gate457inter4));
  nand2 gate790(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate791(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate792(.a(G20), .O(gate457inter7));
  inv1  gate793(.a(G1189), .O(gate457inter8));
  nand2 gate794(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate795(.a(s_35), .b(gate457inter3), .O(gate457inter10));
  nor2  gate796(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate797(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate798(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1989(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1990(.a(gate459inter0), .b(s_206), .O(gate459inter1));
  and2  gate1991(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1992(.a(s_206), .O(gate459inter3));
  inv1  gate1993(.a(s_207), .O(gate459inter4));
  nand2 gate1994(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1995(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1996(.a(G21), .O(gate459inter7));
  inv1  gate1997(.a(G1192), .O(gate459inter8));
  nand2 gate1998(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1999(.a(s_207), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2000(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2001(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2002(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate2311(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2312(.a(gate460inter0), .b(s_252), .O(gate460inter1));
  and2  gate2313(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2314(.a(s_252), .O(gate460inter3));
  inv1  gate2315(.a(s_253), .O(gate460inter4));
  nand2 gate2316(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2317(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2318(.a(G1096), .O(gate460inter7));
  inv1  gate2319(.a(G1192), .O(gate460inter8));
  nand2 gate2320(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2321(.a(s_253), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2322(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2323(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2324(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate1737(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1738(.a(gate461inter0), .b(s_170), .O(gate461inter1));
  and2  gate1739(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1740(.a(s_170), .O(gate461inter3));
  inv1  gate1741(.a(s_171), .O(gate461inter4));
  nand2 gate1742(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1743(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1744(.a(G22), .O(gate461inter7));
  inv1  gate1745(.a(G1195), .O(gate461inter8));
  nand2 gate1746(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1747(.a(s_171), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1748(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1749(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1750(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate729(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate730(.a(gate463inter0), .b(s_26), .O(gate463inter1));
  and2  gate731(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate732(.a(s_26), .O(gate463inter3));
  inv1  gate733(.a(s_27), .O(gate463inter4));
  nand2 gate734(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate735(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate736(.a(G23), .O(gate463inter7));
  inv1  gate737(.a(G1198), .O(gate463inter8));
  nand2 gate738(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate739(.a(s_27), .b(gate463inter3), .O(gate463inter10));
  nor2  gate740(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate741(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate742(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2437(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2438(.a(gate467inter0), .b(s_270), .O(gate467inter1));
  and2  gate2439(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2440(.a(s_270), .O(gate467inter3));
  inv1  gate2441(.a(s_271), .O(gate467inter4));
  nand2 gate2442(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2443(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2444(.a(G25), .O(gate467inter7));
  inv1  gate2445(.a(G1204), .O(gate467inter8));
  nand2 gate2446(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2447(.a(s_271), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2448(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2449(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2450(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2563(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2564(.a(gate469inter0), .b(s_288), .O(gate469inter1));
  and2  gate2565(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2566(.a(s_288), .O(gate469inter3));
  inv1  gate2567(.a(s_289), .O(gate469inter4));
  nand2 gate2568(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2569(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2570(.a(G26), .O(gate469inter7));
  inv1  gate2571(.a(G1207), .O(gate469inter8));
  nand2 gate2572(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2573(.a(s_289), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2574(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2575(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2576(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate981(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate982(.a(gate471inter0), .b(s_62), .O(gate471inter1));
  and2  gate983(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate984(.a(s_62), .O(gate471inter3));
  inv1  gate985(.a(s_63), .O(gate471inter4));
  nand2 gate986(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate987(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate988(.a(G27), .O(gate471inter7));
  inv1  gate989(.a(G1210), .O(gate471inter8));
  nand2 gate990(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate991(.a(s_63), .b(gate471inter3), .O(gate471inter10));
  nor2  gate992(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate993(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate994(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1135(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1136(.a(gate473inter0), .b(s_84), .O(gate473inter1));
  and2  gate1137(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1138(.a(s_84), .O(gate473inter3));
  inv1  gate1139(.a(s_85), .O(gate473inter4));
  nand2 gate1140(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1141(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1142(.a(G28), .O(gate473inter7));
  inv1  gate1143(.a(G1213), .O(gate473inter8));
  nand2 gate1144(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1145(.a(s_85), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1146(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1147(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1148(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate1051(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1052(.a(gate474inter0), .b(s_72), .O(gate474inter1));
  and2  gate1053(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1054(.a(s_72), .O(gate474inter3));
  inv1  gate1055(.a(s_73), .O(gate474inter4));
  nand2 gate1056(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1057(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1058(.a(G1117), .O(gate474inter7));
  inv1  gate1059(.a(G1213), .O(gate474inter8));
  nand2 gate1060(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1061(.a(s_73), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1062(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1063(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1064(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1107(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1108(.a(gate476inter0), .b(s_80), .O(gate476inter1));
  and2  gate1109(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1110(.a(s_80), .O(gate476inter3));
  inv1  gate1111(.a(s_81), .O(gate476inter4));
  nand2 gate1112(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1113(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1114(.a(G1120), .O(gate476inter7));
  inv1  gate1115(.a(G1216), .O(gate476inter8));
  nand2 gate1116(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1117(.a(s_81), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1118(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1119(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1120(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate757(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate758(.a(gate478inter0), .b(s_30), .O(gate478inter1));
  and2  gate759(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate760(.a(s_30), .O(gate478inter3));
  inv1  gate761(.a(s_31), .O(gate478inter4));
  nand2 gate762(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate763(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate764(.a(G1123), .O(gate478inter7));
  inv1  gate765(.a(G1219), .O(gate478inter8));
  nand2 gate766(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate767(.a(s_31), .b(gate478inter3), .O(gate478inter10));
  nor2  gate768(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate769(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate770(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2745(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2746(.a(gate480inter0), .b(s_314), .O(gate480inter1));
  and2  gate2747(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2748(.a(s_314), .O(gate480inter3));
  inv1  gate2749(.a(s_315), .O(gate480inter4));
  nand2 gate2750(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2751(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2752(.a(G1126), .O(gate480inter7));
  inv1  gate2753(.a(G1222), .O(gate480inter8));
  nand2 gate2754(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2755(.a(s_315), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2756(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2757(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2758(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2129(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2130(.a(gate485inter0), .b(s_226), .O(gate485inter1));
  and2  gate2131(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2132(.a(s_226), .O(gate485inter3));
  inv1  gate2133(.a(s_227), .O(gate485inter4));
  nand2 gate2134(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2135(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2136(.a(G1232), .O(gate485inter7));
  inv1  gate2137(.a(G1233), .O(gate485inter8));
  nand2 gate2138(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2139(.a(s_227), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2140(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2141(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2142(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate771(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate772(.a(gate487inter0), .b(s_32), .O(gate487inter1));
  and2  gate773(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate774(.a(s_32), .O(gate487inter3));
  inv1  gate775(.a(s_33), .O(gate487inter4));
  nand2 gate776(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate777(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate778(.a(G1236), .O(gate487inter7));
  inv1  gate779(.a(G1237), .O(gate487inter8));
  nand2 gate780(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate781(.a(s_33), .b(gate487inter3), .O(gate487inter10));
  nor2  gate782(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate783(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate784(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate3081(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate3082(.a(gate489inter0), .b(s_362), .O(gate489inter1));
  and2  gate3083(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate3084(.a(s_362), .O(gate489inter3));
  inv1  gate3085(.a(s_363), .O(gate489inter4));
  nand2 gate3086(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate3087(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate3088(.a(G1240), .O(gate489inter7));
  inv1  gate3089(.a(G1241), .O(gate489inter8));
  nand2 gate3090(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate3091(.a(s_363), .b(gate489inter3), .O(gate489inter10));
  nor2  gate3092(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate3093(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate3094(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1121(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1122(.a(gate490inter0), .b(s_82), .O(gate490inter1));
  and2  gate1123(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1124(.a(s_82), .O(gate490inter3));
  inv1  gate1125(.a(s_83), .O(gate490inter4));
  nand2 gate1126(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1127(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1128(.a(G1242), .O(gate490inter7));
  inv1  gate1129(.a(G1243), .O(gate490inter8));
  nand2 gate1130(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1131(.a(s_83), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1132(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1133(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1134(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2213(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2214(.a(gate493inter0), .b(s_238), .O(gate493inter1));
  and2  gate2215(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2216(.a(s_238), .O(gate493inter3));
  inv1  gate2217(.a(s_239), .O(gate493inter4));
  nand2 gate2218(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2219(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2220(.a(G1248), .O(gate493inter7));
  inv1  gate2221(.a(G1249), .O(gate493inter8));
  nand2 gate2222(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2223(.a(s_239), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2224(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2225(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2226(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2689(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2690(.a(gate494inter0), .b(s_306), .O(gate494inter1));
  and2  gate2691(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2692(.a(s_306), .O(gate494inter3));
  inv1  gate2693(.a(s_307), .O(gate494inter4));
  nand2 gate2694(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2695(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2696(.a(G1250), .O(gate494inter7));
  inv1  gate2697(.a(G1251), .O(gate494inter8));
  nand2 gate2698(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2699(.a(s_307), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2700(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2701(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2702(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1037(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1038(.a(gate501inter0), .b(s_70), .O(gate501inter1));
  and2  gate1039(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1040(.a(s_70), .O(gate501inter3));
  inv1  gate1041(.a(s_71), .O(gate501inter4));
  nand2 gate1042(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1043(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1044(.a(G1264), .O(gate501inter7));
  inv1  gate1045(.a(G1265), .O(gate501inter8));
  nand2 gate1046(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1047(.a(s_71), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1048(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1049(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1050(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate3207(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate3208(.a(gate503inter0), .b(s_380), .O(gate503inter1));
  and2  gate3209(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate3210(.a(s_380), .O(gate503inter3));
  inv1  gate3211(.a(s_381), .O(gate503inter4));
  nand2 gate3212(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate3213(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate3214(.a(G1268), .O(gate503inter7));
  inv1  gate3215(.a(G1269), .O(gate503inter8));
  nand2 gate3216(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate3217(.a(s_381), .b(gate503inter3), .O(gate503inter10));
  nor2  gate3218(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate3219(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate3220(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate3179(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate3180(.a(gate505inter0), .b(s_376), .O(gate505inter1));
  and2  gate3181(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate3182(.a(s_376), .O(gate505inter3));
  inv1  gate3183(.a(s_377), .O(gate505inter4));
  nand2 gate3184(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate3185(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate3186(.a(G1272), .O(gate505inter7));
  inv1  gate3187(.a(G1273), .O(gate505inter8));
  nand2 gate3188(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate3189(.a(s_377), .b(gate505inter3), .O(gate505inter10));
  nor2  gate3190(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate3191(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate3192(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1023(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1024(.a(gate507inter0), .b(s_68), .O(gate507inter1));
  and2  gate1025(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1026(.a(s_68), .O(gate507inter3));
  inv1  gate1027(.a(s_69), .O(gate507inter4));
  nand2 gate1028(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1029(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1030(.a(G1276), .O(gate507inter7));
  inv1  gate1031(.a(G1277), .O(gate507inter8));
  nand2 gate1032(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1033(.a(s_69), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1034(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1035(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1036(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2647(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2648(.a(gate508inter0), .b(s_300), .O(gate508inter1));
  and2  gate2649(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2650(.a(s_300), .O(gate508inter3));
  inv1  gate2651(.a(s_301), .O(gate508inter4));
  nand2 gate2652(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2653(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2654(.a(G1278), .O(gate508inter7));
  inv1  gate2655(.a(G1279), .O(gate508inter8));
  nand2 gate2656(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2657(.a(s_301), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2658(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2659(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2660(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2661(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2662(.a(gate510inter0), .b(s_302), .O(gate510inter1));
  and2  gate2663(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2664(.a(s_302), .O(gate510inter3));
  inv1  gate2665(.a(s_303), .O(gate510inter4));
  nand2 gate2666(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2667(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2668(.a(G1282), .O(gate510inter7));
  inv1  gate2669(.a(G1283), .O(gate510inter8));
  nand2 gate2670(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2671(.a(s_303), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2672(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2673(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2674(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1961(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1962(.a(gate512inter0), .b(s_202), .O(gate512inter1));
  and2  gate1963(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1964(.a(s_202), .O(gate512inter3));
  inv1  gate1965(.a(s_203), .O(gate512inter4));
  nand2 gate1966(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1967(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1968(.a(G1286), .O(gate512inter7));
  inv1  gate1969(.a(G1287), .O(gate512inter8));
  nand2 gate1970(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1971(.a(s_203), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1972(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1973(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1974(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate2423(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2424(.a(gate513inter0), .b(s_268), .O(gate513inter1));
  and2  gate2425(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2426(.a(s_268), .O(gate513inter3));
  inv1  gate2427(.a(s_269), .O(gate513inter4));
  nand2 gate2428(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2429(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2430(.a(G1288), .O(gate513inter7));
  inv1  gate2431(.a(G1289), .O(gate513inter8));
  nand2 gate2432(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2433(.a(s_269), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2434(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2435(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2436(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule