module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate771(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate772(.a(gate12inter0), .b(s_32), .O(gate12inter1));
  and2  gate773(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate774(.a(s_32), .O(gate12inter3));
  inv1  gate775(.a(s_33), .O(gate12inter4));
  nand2 gate776(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate777(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate778(.a(G7), .O(gate12inter7));
  inv1  gate779(.a(G8), .O(gate12inter8));
  nand2 gate780(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate781(.a(s_33), .b(gate12inter3), .O(gate12inter10));
  nor2  gate782(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate783(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate784(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1289(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1290(.a(gate13inter0), .b(s_106), .O(gate13inter1));
  and2  gate1291(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1292(.a(s_106), .O(gate13inter3));
  inv1  gate1293(.a(s_107), .O(gate13inter4));
  nand2 gate1294(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1295(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1296(.a(G9), .O(gate13inter7));
  inv1  gate1297(.a(G10), .O(gate13inter8));
  nand2 gate1298(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1299(.a(s_107), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1300(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1301(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1302(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1919(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1920(.a(gate15inter0), .b(s_196), .O(gate15inter1));
  and2  gate1921(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1922(.a(s_196), .O(gate15inter3));
  inv1  gate1923(.a(s_197), .O(gate15inter4));
  nand2 gate1924(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1925(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1926(.a(G13), .O(gate15inter7));
  inv1  gate1927(.a(G14), .O(gate15inter8));
  nand2 gate1928(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1929(.a(s_197), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1930(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1931(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1932(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2465(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2466(.a(gate16inter0), .b(s_274), .O(gate16inter1));
  and2  gate2467(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2468(.a(s_274), .O(gate16inter3));
  inv1  gate2469(.a(s_275), .O(gate16inter4));
  nand2 gate2470(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2471(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2472(.a(G15), .O(gate16inter7));
  inv1  gate2473(.a(G16), .O(gate16inter8));
  nand2 gate2474(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2475(.a(s_275), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2476(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2477(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2478(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2213(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2214(.a(gate17inter0), .b(s_238), .O(gate17inter1));
  and2  gate2215(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2216(.a(s_238), .O(gate17inter3));
  inv1  gate2217(.a(s_239), .O(gate17inter4));
  nand2 gate2218(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2219(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2220(.a(G17), .O(gate17inter7));
  inv1  gate2221(.a(G18), .O(gate17inter8));
  nand2 gate2222(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2223(.a(s_239), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2224(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2225(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2226(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1079(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1080(.a(gate18inter0), .b(s_76), .O(gate18inter1));
  and2  gate1081(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1082(.a(s_76), .O(gate18inter3));
  inv1  gate1083(.a(s_77), .O(gate18inter4));
  nand2 gate1084(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1085(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1086(.a(G19), .O(gate18inter7));
  inv1  gate1087(.a(G20), .O(gate18inter8));
  nand2 gate1088(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1089(.a(s_77), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1090(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1091(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1092(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1933(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1934(.a(gate22inter0), .b(s_198), .O(gate22inter1));
  and2  gate1935(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1936(.a(s_198), .O(gate22inter3));
  inv1  gate1937(.a(s_199), .O(gate22inter4));
  nand2 gate1938(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1939(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1940(.a(G27), .O(gate22inter7));
  inv1  gate1941(.a(G28), .O(gate22inter8));
  nand2 gate1942(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1943(.a(s_199), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1944(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1945(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1946(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1261(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1262(.a(gate23inter0), .b(s_102), .O(gate23inter1));
  and2  gate1263(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1264(.a(s_102), .O(gate23inter3));
  inv1  gate1265(.a(s_103), .O(gate23inter4));
  nand2 gate1266(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1267(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1268(.a(G29), .O(gate23inter7));
  inv1  gate1269(.a(G30), .O(gate23inter8));
  nand2 gate1270(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1271(.a(s_103), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1272(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1273(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1274(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2185(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2186(.a(gate24inter0), .b(s_234), .O(gate24inter1));
  and2  gate2187(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2188(.a(s_234), .O(gate24inter3));
  inv1  gate2189(.a(s_235), .O(gate24inter4));
  nand2 gate2190(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2191(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2192(.a(G31), .O(gate24inter7));
  inv1  gate2193(.a(G32), .O(gate24inter8));
  nand2 gate2194(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2195(.a(s_235), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2196(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2197(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2198(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1597(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1598(.a(gate30inter0), .b(s_150), .O(gate30inter1));
  and2  gate1599(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1600(.a(s_150), .O(gate30inter3));
  inv1  gate1601(.a(s_151), .O(gate30inter4));
  nand2 gate1602(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1603(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1604(.a(G11), .O(gate30inter7));
  inv1  gate1605(.a(G15), .O(gate30inter8));
  nand2 gate1606(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1607(.a(s_151), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1608(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1609(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1610(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1191(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1192(.a(gate36inter0), .b(s_92), .O(gate36inter1));
  and2  gate1193(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1194(.a(s_92), .O(gate36inter3));
  inv1  gate1195(.a(s_93), .O(gate36inter4));
  nand2 gate1196(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1197(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1198(.a(G26), .O(gate36inter7));
  inv1  gate1199(.a(G30), .O(gate36inter8));
  nand2 gate1200(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1201(.a(s_93), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1202(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1203(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1204(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1625(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1626(.a(gate37inter0), .b(s_154), .O(gate37inter1));
  and2  gate1627(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1628(.a(s_154), .O(gate37inter3));
  inv1  gate1629(.a(s_155), .O(gate37inter4));
  nand2 gate1630(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1631(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1632(.a(G19), .O(gate37inter7));
  inv1  gate1633(.a(G23), .O(gate37inter8));
  nand2 gate1634(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1635(.a(s_155), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1636(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1637(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1638(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate701(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate702(.a(gate40inter0), .b(s_22), .O(gate40inter1));
  and2  gate703(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate704(.a(s_22), .O(gate40inter3));
  inv1  gate705(.a(s_23), .O(gate40inter4));
  nand2 gate706(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate707(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate708(.a(G28), .O(gate40inter7));
  inv1  gate709(.a(G32), .O(gate40inter8));
  nand2 gate710(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate711(.a(s_23), .b(gate40inter3), .O(gate40inter10));
  nor2  gate712(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate713(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate714(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1247(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1248(.a(gate41inter0), .b(s_100), .O(gate41inter1));
  and2  gate1249(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1250(.a(s_100), .O(gate41inter3));
  inv1  gate1251(.a(s_101), .O(gate41inter4));
  nand2 gate1252(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1253(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1254(.a(G1), .O(gate41inter7));
  inv1  gate1255(.a(G266), .O(gate41inter8));
  nand2 gate1256(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1257(.a(s_101), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1258(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1259(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1260(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1695(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1696(.a(gate42inter0), .b(s_164), .O(gate42inter1));
  and2  gate1697(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1698(.a(s_164), .O(gate42inter3));
  inv1  gate1699(.a(s_165), .O(gate42inter4));
  nand2 gate1700(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1701(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1702(.a(G2), .O(gate42inter7));
  inv1  gate1703(.a(G266), .O(gate42inter8));
  nand2 gate1704(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1705(.a(s_165), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1706(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1707(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1708(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1639(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1640(.a(gate43inter0), .b(s_156), .O(gate43inter1));
  and2  gate1641(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1642(.a(s_156), .O(gate43inter3));
  inv1  gate1643(.a(s_157), .O(gate43inter4));
  nand2 gate1644(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1645(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1646(.a(G3), .O(gate43inter7));
  inv1  gate1647(.a(G269), .O(gate43inter8));
  nand2 gate1648(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1649(.a(s_157), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1650(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1651(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1652(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1051(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1052(.a(gate47inter0), .b(s_72), .O(gate47inter1));
  and2  gate1053(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1054(.a(s_72), .O(gate47inter3));
  inv1  gate1055(.a(s_73), .O(gate47inter4));
  nand2 gate1056(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1057(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1058(.a(G7), .O(gate47inter7));
  inv1  gate1059(.a(G275), .O(gate47inter8));
  nand2 gate1060(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1061(.a(s_73), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1062(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1063(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1064(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1331(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1332(.a(gate50inter0), .b(s_112), .O(gate50inter1));
  and2  gate1333(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1334(.a(s_112), .O(gate50inter3));
  inv1  gate1335(.a(s_113), .O(gate50inter4));
  nand2 gate1336(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1337(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1338(.a(G10), .O(gate50inter7));
  inv1  gate1339(.a(G278), .O(gate50inter8));
  nand2 gate1340(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1341(.a(s_113), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1342(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1343(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1344(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1765(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1766(.a(gate53inter0), .b(s_174), .O(gate53inter1));
  and2  gate1767(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1768(.a(s_174), .O(gate53inter3));
  inv1  gate1769(.a(s_175), .O(gate53inter4));
  nand2 gate1770(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1771(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1772(.a(G13), .O(gate53inter7));
  inv1  gate1773(.a(G284), .O(gate53inter8));
  nand2 gate1774(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1775(.a(s_175), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1776(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1777(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1778(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate953(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate954(.a(gate55inter0), .b(s_58), .O(gate55inter1));
  and2  gate955(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate956(.a(s_58), .O(gate55inter3));
  inv1  gate957(.a(s_59), .O(gate55inter4));
  nand2 gate958(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate959(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate960(.a(G15), .O(gate55inter7));
  inv1  gate961(.a(G287), .O(gate55inter8));
  nand2 gate962(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate963(.a(s_59), .b(gate55inter3), .O(gate55inter10));
  nor2  gate964(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate965(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate966(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1989(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1990(.a(gate64inter0), .b(s_206), .O(gate64inter1));
  and2  gate1991(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1992(.a(s_206), .O(gate64inter3));
  inv1  gate1993(.a(s_207), .O(gate64inter4));
  nand2 gate1994(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1995(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1996(.a(G24), .O(gate64inter7));
  inv1  gate1997(.a(G299), .O(gate64inter8));
  nand2 gate1998(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1999(.a(s_207), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2000(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2001(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2002(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1163(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1164(.a(gate66inter0), .b(s_88), .O(gate66inter1));
  and2  gate1165(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1166(.a(s_88), .O(gate66inter3));
  inv1  gate1167(.a(s_89), .O(gate66inter4));
  nand2 gate1168(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1169(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1170(.a(G26), .O(gate66inter7));
  inv1  gate1171(.a(G302), .O(gate66inter8));
  nand2 gate1172(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1173(.a(s_89), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1174(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1175(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1176(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1443(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1444(.a(gate67inter0), .b(s_128), .O(gate67inter1));
  and2  gate1445(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1446(.a(s_128), .O(gate67inter3));
  inv1  gate1447(.a(s_129), .O(gate67inter4));
  nand2 gate1448(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1449(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1450(.a(G27), .O(gate67inter7));
  inv1  gate1451(.a(G305), .O(gate67inter8));
  nand2 gate1452(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1453(.a(s_129), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1454(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1455(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1456(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1121(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1122(.a(gate74inter0), .b(s_82), .O(gate74inter1));
  and2  gate1123(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1124(.a(s_82), .O(gate74inter3));
  inv1  gate1125(.a(s_83), .O(gate74inter4));
  nand2 gate1126(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1127(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1128(.a(G5), .O(gate74inter7));
  inv1  gate1129(.a(G314), .O(gate74inter8));
  nand2 gate1130(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1131(.a(s_83), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1132(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1133(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1134(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1527(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1528(.a(gate75inter0), .b(s_140), .O(gate75inter1));
  and2  gate1529(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1530(.a(s_140), .O(gate75inter3));
  inv1  gate1531(.a(s_141), .O(gate75inter4));
  nand2 gate1532(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1533(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1534(.a(G9), .O(gate75inter7));
  inv1  gate1535(.a(G317), .O(gate75inter8));
  nand2 gate1536(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1537(.a(s_141), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1538(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1539(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1540(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1751(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1752(.a(gate77inter0), .b(s_172), .O(gate77inter1));
  and2  gate1753(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1754(.a(s_172), .O(gate77inter3));
  inv1  gate1755(.a(s_173), .O(gate77inter4));
  nand2 gate1756(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1757(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1758(.a(G2), .O(gate77inter7));
  inv1  gate1759(.a(G320), .O(gate77inter8));
  nand2 gate1760(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1761(.a(s_173), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1762(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1763(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1764(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate2437(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2438(.a(gate78inter0), .b(s_270), .O(gate78inter1));
  and2  gate2439(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2440(.a(s_270), .O(gate78inter3));
  inv1  gate2441(.a(s_271), .O(gate78inter4));
  nand2 gate2442(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2443(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2444(.a(G6), .O(gate78inter7));
  inv1  gate2445(.a(G320), .O(gate78inter8));
  nand2 gate2446(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2447(.a(s_271), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2448(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2449(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2450(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2395(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2396(.a(gate81inter0), .b(s_264), .O(gate81inter1));
  and2  gate2397(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2398(.a(s_264), .O(gate81inter3));
  inv1  gate2399(.a(s_265), .O(gate81inter4));
  nand2 gate2400(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2401(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2402(.a(G3), .O(gate81inter7));
  inv1  gate2403(.a(G326), .O(gate81inter8));
  nand2 gate2404(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2405(.a(s_265), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2406(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2407(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2408(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate561(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate562(.a(gate82inter0), .b(s_2), .O(gate82inter1));
  and2  gate563(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate564(.a(s_2), .O(gate82inter3));
  inv1  gate565(.a(s_3), .O(gate82inter4));
  nand2 gate566(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate567(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate568(.a(G7), .O(gate82inter7));
  inv1  gate569(.a(G326), .O(gate82inter8));
  nand2 gate570(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate571(.a(s_3), .b(gate82inter3), .O(gate82inter10));
  nor2  gate572(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate573(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate574(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1793(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1794(.a(gate83inter0), .b(s_178), .O(gate83inter1));
  and2  gate1795(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1796(.a(s_178), .O(gate83inter3));
  inv1  gate1797(.a(s_179), .O(gate83inter4));
  nand2 gate1798(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1799(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1800(.a(G11), .O(gate83inter7));
  inv1  gate1801(.a(G329), .O(gate83inter8));
  nand2 gate1802(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1803(.a(s_179), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1804(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1805(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1806(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1093(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1094(.a(gate88inter0), .b(s_78), .O(gate88inter1));
  and2  gate1095(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1096(.a(s_78), .O(gate88inter3));
  inv1  gate1097(.a(s_79), .O(gate88inter4));
  nand2 gate1098(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1099(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1100(.a(G16), .O(gate88inter7));
  inv1  gate1101(.a(G335), .O(gate88inter8));
  nand2 gate1102(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1103(.a(s_79), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1104(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1105(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1106(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1485(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1486(.a(gate94inter0), .b(s_134), .O(gate94inter1));
  and2  gate1487(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1488(.a(s_134), .O(gate94inter3));
  inv1  gate1489(.a(s_135), .O(gate94inter4));
  nand2 gate1490(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1491(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1492(.a(G22), .O(gate94inter7));
  inv1  gate1493(.a(G344), .O(gate94inter8));
  nand2 gate1494(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1495(.a(s_135), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1496(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1497(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1498(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1275(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1276(.a(gate99inter0), .b(s_104), .O(gate99inter1));
  and2  gate1277(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1278(.a(s_104), .O(gate99inter3));
  inv1  gate1279(.a(s_105), .O(gate99inter4));
  nand2 gate1280(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1281(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1282(.a(G27), .O(gate99inter7));
  inv1  gate1283(.a(G353), .O(gate99inter8));
  nand2 gate1284(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1285(.a(s_105), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1286(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1287(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1288(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2157(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2158(.a(gate101inter0), .b(s_230), .O(gate101inter1));
  and2  gate2159(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2160(.a(s_230), .O(gate101inter3));
  inv1  gate2161(.a(s_231), .O(gate101inter4));
  nand2 gate2162(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2163(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2164(.a(G20), .O(gate101inter7));
  inv1  gate2165(.a(G356), .O(gate101inter8));
  nand2 gate2166(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2167(.a(s_231), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2168(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2169(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2170(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2101(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2102(.a(gate102inter0), .b(s_222), .O(gate102inter1));
  and2  gate2103(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2104(.a(s_222), .O(gate102inter3));
  inv1  gate2105(.a(s_223), .O(gate102inter4));
  nand2 gate2106(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2107(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2108(.a(G24), .O(gate102inter7));
  inv1  gate2109(.a(G356), .O(gate102inter8));
  nand2 gate2110(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2111(.a(s_223), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2112(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2113(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2114(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate631(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate632(.a(gate103inter0), .b(s_12), .O(gate103inter1));
  and2  gate633(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate634(.a(s_12), .O(gate103inter3));
  inv1  gate635(.a(s_13), .O(gate103inter4));
  nand2 gate636(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate637(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate638(.a(G28), .O(gate103inter7));
  inv1  gate639(.a(G359), .O(gate103inter8));
  nand2 gate640(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate641(.a(s_13), .b(gate103inter3), .O(gate103inter10));
  nor2  gate642(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate643(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate644(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1975(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1976(.a(gate104inter0), .b(s_204), .O(gate104inter1));
  and2  gate1977(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1978(.a(s_204), .O(gate104inter3));
  inv1  gate1979(.a(s_205), .O(gate104inter4));
  nand2 gate1980(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1981(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1982(.a(G32), .O(gate104inter7));
  inv1  gate1983(.a(G359), .O(gate104inter8));
  nand2 gate1984(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1985(.a(s_205), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1986(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1987(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1988(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate967(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate968(.a(gate108inter0), .b(s_60), .O(gate108inter1));
  and2  gate969(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate970(.a(s_60), .O(gate108inter3));
  inv1  gate971(.a(s_61), .O(gate108inter4));
  nand2 gate972(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate973(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate974(.a(G368), .O(gate108inter7));
  inv1  gate975(.a(G369), .O(gate108inter8));
  nand2 gate976(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate977(.a(s_61), .b(gate108inter3), .O(gate108inter10));
  nor2  gate978(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate979(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate980(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1709(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1710(.a(gate113inter0), .b(s_166), .O(gate113inter1));
  and2  gate1711(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1712(.a(s_166), .O(gate113inter3));
  inv1  gate1713(.a(s_167), .O(gate113inter4));
  nand2 gate1714(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1715(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1716(.a(G378), .O(gate113inter7));
  inv1  gate1717(.a(G379), .O(gate113inter8));
  nand2 gate1718(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1719(.a(s_167), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1720(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1721(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1722(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate2507(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2508(.a(gate116inter0), .b(s_280), .O(gate116inter1));
  and2  gate2509(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2510(.a(s_280), .O(gate116inter3));
  inv1  gate2511(.a(s_281), .O(gate116inter4));
  nand2 gate2512(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2513(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2514(.a(G384), .O(gate116inter7));
  inv1  gate2515(.a(G385), .O(gate116inter8));
  nand2 gate2516(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2517(.a(s_281), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2518(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2519(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2520(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate715(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate716(.a(gate118inter0), .b(s_24), .O(gate118inter1));
  and2  gate717(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate718(.a(s_24), .O(gate118inter3));
  inv1  gate719(.a(s_25), .O(gate118inter4));
  nand2 gate720(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate721(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate722(.a(G388), .O(gate118inter7));
  inv1  gate723(.a(G389), .O(gate118inter8));
  nand2 gate724(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate725(.a(s_25), .b(gate118inter3), .O(gate118inter10));
  nor2  gate726(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate727(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate728(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1863(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1864(.a(gate119inter0), .b(s_188), .O(gate119inter1));
  and2  gate1865(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1866(.a(s_188), .O(gate119inter3));
  inv1  gate1867(.a(s_189), .O(gate119inter4));
  nand2 gate1868(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1869(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1870(.a(G390), .O(gate119inter7));
  inv1  gate1871(.a(G391), .O(gate119inter8));
  nand2 gate1872(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1873(.a(s_189), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1874(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1875(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1876(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate785(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate786(.a(gate120inter0), .b(s_34), .O(gate120inter1));
  and2  gate787(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate788(.a(s_34), .O(gate120inter3));
  inv1  gate789(.a(s_35), .O(gate120inter4));
  nand2 gate790(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate791(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate792(.a(G392), .O(gate120inter7));
  inv1  gate793(.a(G393), .O(gate120inter8));
  nand2 gate794(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate795(.a(s_35), .b(gate120inter3), .O(gate120inter10));
  nor2  gate796(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate797(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate798(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1205(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1206(.a(gate124inter0), .b(s_94), .O(gate124inter1));
  and2  gate1207(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1208(.a(s_94), .O(gate124inter3));
  inv1  gate1209(.a(s_95), .O(gate124inter4));
  nand2 gate1210(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1211(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1212(.a(G400), .O(gate124inter7));
  inv1  gate1213(.a(G401), .O(gate124inter8));
  nand2 gate1214(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1215(.a(s_95), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1216(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1217(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1218(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1359(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1360(.a(gate126inter0), .b(s_116), .O(gate126inter1));
  and2  gate1361(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1362(.a(s_116), .O(gate126inter3));
  inv1  gate1363(.a(s_117), .O(gate126inter4));
  nand2 gate1364(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1365(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1366(.a(G404), .O(gate126inter7));
  inv1  gate1367(.a(G405), .O(gate126inter8));
  nand2 gate1368(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1369(.a(s_117), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1370(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1371(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1372(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1233(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1234(.a(gate129inter0), .b(s_98), .O(gate129inter1));
  and2  gate1235(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1236(.a(s_98), .O(gate129inter3));
  inv1  gate1237(.a(s_99), .O(gate129inter4));
  nand2 gate1238(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1239(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1240(.a(G410), .O(gate129inter7));
  inv1  gate1241(.a(G411), .O(gate129inter8));
  nand2 gate1242(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1243(.a(s_99), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1244(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1245(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1246(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate743(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate744(.a(gate133inter0), .b(s_28), .O(gate133inter1));
  and2  gate745(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate746(.a(s_28), .O(gate133inter3));
  inv1  gate747(.a(s_29), .O(gate133inter4));
  nand2 gate748(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate749(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate750(.a(G418), .O(gate133inter7));
  inv1  gate751(.a(G419), .O(gate133inter8));
  nand2 gate752(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate753(.a(s_29), .b(gate133inter3), .O(gate133inter10));
  nor2  gate754(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate755(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate756(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1401(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1402(.a(gate135inter0), .b(s_122), .O(gate135inter1));
  and2  gate1403(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1404(.a(s_122), .O(gate135inter3));
  inv1  gate1405(.a(s_123), .O(gate135inter4));
  nand2 gate1406(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1407(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1408(.a(G422), .O(gate135inter7));
  inv1  gate1409(.a(G423), .O(gate135inter8));
  nand2 gate1410(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1411(.a(s_123), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1412(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1413(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1414(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1583(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1584(.a(gate138inter0), .b(s_148), .O(gate138inter1));
  and2  gate1585(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1586(.a(s_148), .O(gate138inter3));
  inv1  gate1587(.a(s_149), .O(gate138inter4));
  nand2 gate1588(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1589(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1590(.a(G432), .O(gate138inter7));
  inv1  gate1591(.a(G435), .O(gate138inter8));
  nand2 gate1592(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1593(.a(s_149), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1594(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1595(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1596(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate757(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate758(.a(gate139inter0), .b(s_30), .O(gate139inter1));
  and2  gate759(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate760(.a(s_30), .O(gate139inter3));
  inv1  gate761(.a(s_31), .O(gate139inter4));
  nand2 gate762(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate763(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate764(.a(G438), .O(gate139inter7));
  inv1  gate765(.a(G441), .O(gate139inter8));
  nand2 gate766(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate767(.a(s_31), .b(gate139inter3), .O(gate139inter10));
  nor2  gate768(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate769(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate770(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2115(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2116(.a(gate143inter0), .b(s_224), .O(gate143inter1));
  and2  gate2117(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2118(.a(s_224), .O(gate143inter3));
  inv1  gate2119(.a(s_225), .O(gate143inter4));
  nand2 gate2120(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2121(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2122(.a(G462), .O(gate143inter7));
  inv1  gate2123(.a(G465), .O(gate143inter8));
  nand2 gate2124(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2125(.a(s_225), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2126(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2127(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2128(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate911(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate912(.a(gate147inter0), .b(s_52), .O(gate147inter1));
  and2  gate913(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate914(.a(s_52), .O(gate147inter3));
  inv1  gate915(.a(s_53), .O(gate147inter4));
  nand2 gate916(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate917(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate918(.a(G486), .O(gate147inter7));
  inv1  gate919(.a(G489), .O(gate147inter8));
  nand2 gate920(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate921(.a(s_53), .b(gate147inter3), .O(gate147inter10));
  nor2  gate922(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate923(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate924(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate869(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate870(.a(gate150inter0), .b(s_46), .O(gate150inter1));
  and2  gate871(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate872(.a(s_46), .O(gate150inter3));
  inv1  gate873(.a(s_47), .O(gate150inter4));
  nand2 gate874(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate875(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate876(.a(G504), .O(gate150inter7));
  inv1  gate877(.a(G507), .O(gate150inter8));
  nand2 gate878(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate879(.a(s_47), .b(gate150inter3), .O(gate150inter10));
  nor2  gate880(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate881(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate882(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2269(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2270(.a(gate151inter0), .b(s_246), .O(gate151inter1));
  and2  gate2271(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2272(.a(s_246), .O(gate151inter3));
  inv1  gate2273(.a(s_247), .O(gate151inter4));
  nand2 gate2274(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2275(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2276(.a(G510), .O(gate151inter7));
  inv1  gate2277(.a(G513), .O(gate151inter8));
  nand2 gate2278(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2279(.a(s_247), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2280(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2281(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2282(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2171(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2172(.a(gate152inter0), .b(s_232), .O(gate152inter1));
  and2  gate2173(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2174(.a(s_232), .O(gate152inter3));
  inv1  gate2175(.a(s_233), .O(gate152inter4));
  nand2 gate2176(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2177(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2178(.a(G516), .O(gate152inter7));
  inv1  gate2179(.a(G519), .O(gate152inter8));
  nand2 gate2180(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2181(.a(s_233), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2182(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2183(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2184(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1611(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1612(.a(gate156inter0), .b(s_152), .O(gate156inter1));
  and2  gate1613(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1614(.a(s_152), .O(gate156inter3));
  inv1  gate1615(.a(s_153), .O(gate156inter4));
  nand2 gate1616(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1617(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1618(.a(G435), .O(gate156inter7));
  inv1  gate1619(.a(G525), .O(gate156inter8));
  nand2 gate1620(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1621(.a(s_153), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1622(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1623(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1624(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate827(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate828(.a(gate160inter0), .b(s_40), .O(gate160inter1));
  and2  gate829(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate830(.a(s_40), .O(gate160inter3));
  inv1  gate831(.a(s_41), .O(gate160inter4));
  nand2 gate832(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate833(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate834(.a(G447), .O(gate160inter7));
  inv1  gate835(.a(G531), .O(gate160inter8));
  nand2 gate836(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate837(.a(s_41), .b(gate160inter3), .O(gate160inter10));
  nor2  gate838(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate839(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate840(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate2227(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2228(.a(gate161inter0), .b(s_240), .O(gate161inter1));
  and2  gate2229(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2230(.a(s_240), .O(gate161inter3));
  inv1  gate2231(.a(s_241), .O(gate161inter4));
  nand2 gate2232(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2233(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2234(.a(G450), .O(gate161inter7));
  inv1  gate2235(.a(G534), .O(gate161inter8));
  nand2 gate2236(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2237(.a(s_241), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2238(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2239(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2240(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2059(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2060(.a(gate167inter0), .b(s_216), .O(gate167inter1));
  and2  gate2061(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2062(.a(s_216), .O(gate167inter3));
  inv1  gate2063(.a(s_217), .O(gate167inter4));
  nand2 gate2064(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2065(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2066(.a(G468), .O(gate167inter7));
  inv1  gate2067(.a(G543), .O(gate167inter8));
  nand2 gate2068(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2069(.a(s_217), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2070(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2071(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2072(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1135(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1136(.a(gate168inter0), .b(s_84), .O(gate168inter1));
  and2  gate1137(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1138(.a(s_84), .O(gate168inter3));
  inv1  gate1139(.a(s_85), .O(gate168inter4));
  nand2 gate1140(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1141(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1142(.a(G471), .O(gate168inter7));
  inv1  gate1143(.a(G543), .O(gate168inter8));
  nand2 gate1144(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1145(.a(s_85), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1146(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1147(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1148(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1555(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1556(.a(gate171inter0), .b(s_144), .O(gate171inter1));
  and2  gate1557(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1558(.a(s_144), .O(gate171inter3));
  inv1  gate1559(.a(s_145), .O(gate171inter4));
  nand2 gate1560(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1561(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1562(.a(G480), .O(gate171inter7));
  inv1  gate1563(.a(G549), .O(gate171inter8));
  nand2 gate1564(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1565(.a(s_145), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1566(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1567(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1568(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1149(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1150(.a(gate177inter0), .b(s_86), .O(gate177inter1));
  and2  gate1151(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1152(.a(s_86), .O(gate177inter3));
  inv1  gate1153(.a(s_87), .O(gate177inter4));
  nand2 gate1154(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1155(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1156(.a(G498), .O(gate177inter7));
  inv1  gate1157(.a(G558), .O(gate177inter8));
  nand2 gate1158(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1159(.a(s_87), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1160(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1161(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1162(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2409(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2410(.a(gate187inter0), .b(s_266), .O(gate187inter1));
  and2  gate2411(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2412(.a(s_266), .O(gate187inter3));
  inv1  gate2413(.a(s_267), .O(gate187inter4));
  nand2 gate2414(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2415(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2416(.a(G574), .O(gate187inter7));
  inv1  gate2417(.a(G575), .O(gate187inter8));
  nand2 gate2418(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2419(.a(s_267), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2420(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2421(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2422(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2311(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2312(.a(gate189inter0), .b(s_252), .O(gate189inter1));
  and2  gate2313(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2314(.a(s_252), .O(gate189inter3));
  inv1  gate2315(.a(s_253), .O(gate189inter4));
  nand2 gate2316(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2317(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2318(.a(G578), .O(gate189inter7));
  inv1  gate2319(.a(G579), .O(gate189inter8));
  nand2 gate2320(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2321(.a(s_253), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2322(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2323(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2324(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1541(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1542(.a(gate194inter0), .b(s_142), .O(gate194inter1));
  and2  gate1543(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1544(.a(s_142), .O(gate194inter3));
  inv1  gate1545(.a(s_143), .O(gate194inter4));
  nand2 gate1546(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1547(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1548(.a(G588), .O(gate194inter7));
  inv1  gate1549(.a(G589), .O(gate194inter8));
  nand2 gate1550(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1551(.a(s_143), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1552(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1553(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1554(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2325(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2326(.a(gate195inter0), .b(s_254), .O(gate195inter1));
  and2  gate2327(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2328(.a(s_254), .O(gate195inter3));
  inv1  gate2329(.a(s_255), .O(gate195inter4));
  nand2 gate2330(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2331(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2332(.a(G590), .O(gate195inter7));
  inv1  gate2333(.a(G591), .O(gate195inter8));
  nand2 gate2334(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2335(.a(s_255), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2336(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2337(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2338(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1849(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1850(.a(gate196inter0), .b(s_186), .O(gate196inter1));
  and2  gate1851(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1852(.a(s_186), .O(gate196inter3));
  inv1  gate1853(.a(s_187), .O(gate196inter4));
  nand2 gate1854(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1855(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1856(.a(G592), .O(gate196inter7));
  inv1  gate1857(.a(G593), .O(gate196inter8));
  nand2 gate1858(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1859(.a(s_187), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1860(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1861(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1862(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate603(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate604(.a(gate199inter0), .b(s_8), .O(gate199inter1));
  and2  gate605(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate606(.a(s_8), .O(gate199inter3));
  inv1  gate607(.a(s_9), .O(gate199inter4));
  nand2 gate608(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate609(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate610(.a(G598), .O(gate199inter7));
  inv1  gate611(.a(G599), .O(gate199inter8));
  nand2 gate612(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate613(.a(s_9), .b(gate199inter3), .O(gate199inter10));
  nor2  gate614(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate615(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate616(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate813(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate814(.a(gate203inter0), .b(s_38), .O(gate203inter1));
  and2  gate815(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate816(.a(s_38), .O(gate203inter3));
  inv1  gate817(.a(s_39), .O(gate203inter4));
  nand2 gate818(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate819(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate820(.a(G602), .O(gate203inter7));
  inv1  gate821(.a(G612), .O(gate203inter8));
  nand2 gate822(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate823(.a(s_39), .b(gate203inter3), .O(gate203inter10));
  nor2  gate824(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate825(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate826(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1835(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1836(.a(gate204inter0), .b(s_184), .O(gate204inter1));
  and2  gate1837(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1838(.a(s_184), .O(gate204inter3));
  inv1  gate1839(.a(s_185), .O(gate204inter4));
  nand2 gate1840(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1841(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1842(.a(G607), .O(gate204inter7));
  inv1  gate1843(.a(G617), .O(gate204inter8));
  nand2 gate1844(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1845(.a(s_185), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1846(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1847(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1848(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2493(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2494(.a(gate206inter0), .b(s_278), .O(gate206inter1));
  and2  gate2495(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2496(.a(s_278), .O(gate206inter3));
  inv1  gate2497(.a(s_279), .O(gate206inter4));
  nand2 gate2498(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2499(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2500(.a(G632), .O(gate206inter7));
  inv1  gate2501(.a(G637), .O(gate206inter8));
  nand2 gate2502(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2503(.a(s_279), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2504(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2505(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2506(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1737(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1738(.a(gate207inter0), .b(s_170), .O(gate207inter1));
  and2  gate1739(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1740(.a(s_170), .O(gate207inter3));
  inv1  gate1741(.a(s_171), .O(gate207inter4));
  nand2 gate1742(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1743(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1744(.a(G622), .O(gate207inter7));
  inv1  gate1745(.a(G632), .O(gate207inter8));
  nand2 gate1746(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1747(.a(s_171), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1748(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1749(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1750(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2087(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2088(.a(gate208inter0), .b(s_220), .O(gate208inter1));
  and2  gate2089(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2090(.a(s_220), .O(gate208inter3));
  inv1  gate2091(.a(s_221), .O(gate208inter4));
  nand2 gate2092(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2093(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2094(.a(G627), .O(gate208inter7));
  inv1  gate2095(.a(G637), .O(gate208inter8));
  nand2 gate2096(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2097(.a(s_221), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2098(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2099(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2100(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2073(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2074(.a(gate212inter0), .b(s_218), .O(gate212inter1));
  and2  gate2075(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2076(.a(s_218), .O(gate212inter3));
  inv1  gate2077(.a(s_219), .O(gate212inter4));
  nand2 gate2078(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2079(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2080(.a(G617), .O(gate212inter7));
  inv1  gate2081(.a(G669), .O(gate212inter8));
  nand2 gate2082(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2083(.a(s_219), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2084(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2085(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2086(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate897(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate898(.a(gate216inter0), .b(s_50), .O(gate216inter1));
  and2  gate899(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate900(.a(s_50), .O(gate216inter3));
  inv1  gate901(.a(s_51), .O(gate216inter4));
  nand2 gate902(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate903(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate904(.a(G617), .O(gate216inter7));
  inv1  gate905(.a(G675), .O(gate216inter8));
  nand2 gate906(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate907(.a(s_51), .b(gate216inter3), .O(gate216inter10));
  nor2  gate908(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate909(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate910(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate729(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate730(.a(gate217inter0), .b(s_26), .O(gate217inter1));
  and2  gate731(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate732(.a(s_26), .O(gate217inter3));
  inv1  gate733(.a(s_27), .O(gate217inter4));
  nand2 gate734(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate735(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate736(.a(G622), .O(gate217inter7));
  inv1  gate737(.a(G678), .O(gate217inter8));
  nand2 gate738(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate739(.a(s_27), .b(gate217inter3), .O(gate217inter10));
  nor2  gate740(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate741(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate742(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate841(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate842(.a(gate221inter0), .b(s_42), .O(gate221inter1));
  and2  gate843(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate844(.a(s_42), .O(gate221inter3));
  inv1  gate845(.a(s_43), .O(gate221inter4));
  nand2 gate846(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate847(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate848(.a(G622), .O(gate221inter7));
  inv1  gate849(.a(G684), .O(gate221inter8));
  nand2 gate850(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate851(.a(s_43), .b(gate221inter3), .O(gate221inter10));
  nor2  gate852(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate853(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate854(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1429(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1430(.a(gate223inter0), .b(s_126), .O(gate223inter1));
  and2  gate1431(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1432(.a(s_126), .O(gate223inter3));
  inv1  gate1433(.a(s_127), .O(gate223inter4));
  nand2 gate1434(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1435(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1436(.a(G627), .O(gate223inter7));
  inv1  gate1437(.a(G687), .O(gate223inter8));
  nand2 gate1438(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1439(.a(s_127), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1440(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1441(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1442(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2339(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2340(.a(gate227inter0), .b(s_256), .O(gate227inter1));
  and2  gate2341(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2342(.a(s_256), .O(gate227inter3));
  inv1  gate2343(.a(s_257), .O(gate227inter4));
  nand2 gate2344(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2345(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2346(.a(G694), .O(gate227inter7));
  inv1  gate2347(.a(G695), .O(gate227inter8));
  nand2 gate2348(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2349(.a(s_257), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2350(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2351(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2352(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1821(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1822(.a(gate228inter0), .b(s_182), .O(gate228inter1));
  and2  gate1823(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1824(.a(s_182), .O(gate228inter3));
  inv1  gate1825(.a(s_183), .O(gate228inter4));
  nand2 gate1826(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1827(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1828(.a(G696), .O(gate228inter7));
  inv1  gate1829(.a(G697), .O(gate228inter8));
  nand2 gate1830(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1831(.a(s_183), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1832(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1833(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1834(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1653(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1654(.a(gate229inter0), .b(s_158), .O(gate229inter1));
  and2  gate1655(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1656(.a(s_158), .O(gate229inter3));
  inv1  gate1657(.a(s_159), .O(gate229inter4));
  nand2 gate1658(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1659(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1660(.a(G698), .O(gate229inter7));
  inv1  gate1661(.a(G699), .O(gate229inter8));
  nand2 gate1662(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1663(.a(s_159), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1664(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1665(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1666(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2297(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2298(.a(gate237inter0), .b(s_250), .O(gate237inter1));
  and2  gate2299(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2300(.a(s_250), .O(gate237inter3));
  inv1  gate2301(.a(s_251), .O(gate237inter4));
  nand2 gate2302(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2303(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2304(.a(G254), .O(gate237inter7));
  inv1  gate2305(.a(G706), .O(gate237inter8));
  nand2 gate2306(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2307(.a(s_251), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2308(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2309(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2310(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2423(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2424(.a(gate240inter0), .b(s_268), .O(gate240inter1));
  and2  gate2425(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2426(.a(s_268), .O(gate240inter3));
  inv1  gate2427(.a(s_269), .O(gate240inter4));
  nand2 gate2428(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2429(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2430(.a(G263), .O(gate240inter7));
  inv1  gate2431(.a(G715), .O(gate240inter8));
  nand2 gate2432(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2433(.a(s_269), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2434(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2435(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2436(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2017(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2018(.a(gate243inter0), .b(s_210), .O(gate243inter1));
  and2  gate2019(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2020(.a(s_210), .O(gate243inter3));
  inv1  gate2021(.a(s_211), .O(gate243inter4));
  nand2 gate2022(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2023(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2024(.a(G245), .O(gate243inter7));
  inv1  gate2025(.a(G733), .O(gate243inter8));
  nand2 gate2026(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2027(.a(s_211), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2028(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2029(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2030(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2381(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2382(.a(gate249inter0), .b(s_262), .O(gate249inter1));
  and2  gate2383(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2384(.a(s_262), .O(gate249inter3));
  inv1  gate2385(.a(s_263), .O(gate249inter4));
  nand2 gate2386(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2387(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2388(.a(G254), .O(gate249inter7));
  inv1  gate2389(.a(G742), .O(gate249inter8));
  nand2 gate2390(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2391(.a(s_263), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2392(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2393(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2394(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2479(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2480(.a(gate251inter0), .b(s_276), .O(gate251inter1));
  and2  gate2481(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2482(.a(s_276), .O(gate251inter3));
  inv1  gate2483(.a(s_277), .O(gate251inter4));
  nand2 gate2484(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2485(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2486(.a(G257), .O(gate251inter7));
  inv1  gate2487(.a(G745), .O(gate251inter8));
  nand2 gate2488(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2489(.a(s_277), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2490(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2491(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2492(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate995(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate996(.a(gate253inter0), .b(s_64), .O(gate253inter1));
  and2  gate997(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate998(.a(s_64), .O(gate253inter3));
  inv1  gate999(.a(s_65), .O(gate253inter4));
  nand2 gate1000(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1001(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1002(.a(G260), .O(gate253inter7));
  inv1  gate1003(.a(G748), .O(gate253inter8));
  nand2 gate1004(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1005(.a(s_65), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1006(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1007(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1008(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate925(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate926(.a(gate254inter0), .b(s_54), .O(gate254inter1));
  and2  gate927(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate928(.a(s_54), .O(gate254inter3));
  inv1  gate929(.a(s_55), .O(gate254inter4));
  nand2 gate930(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate931(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate932(.a(G712), .O(gate254inter7));
  inv1  gate933(.a(G748), .O(gate254inter8));
  nand2 gate934(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate935(.a(s_55), .b(gate254inter3), .O(gate254inter10));
  nor2  gate936(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate937(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate938(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1303(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1304(.a(gate260inter0), .b(s_108), .O(gate260inter1));
  and2  gate1305(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1306(.a(s_108), .O(gate260inter3));
  inv1  gate1307(.a(s_109), .O(gate260inter4));
  nand2 gate1308(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1309(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1310(.a(G760), .O(gate260inter7));
  inv1  gate1311(.a(G761), .O(gate260inter8));
  nand2 gate1312(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1313(.a(s_109), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1314(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1315(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1316(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2199(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2200(.a(gate261inter0), .b(s_236), .O(gate261inter1));
  and2  gate2201(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2202(.a(s_236), .O(gate261inter3));
  inv1  gate2203(.a(s_237), .O(gate261inter4));
  nand2 gate2204(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2205(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2206(.a(G762), .O(gate261inter7));
  inv1  gate2207(.a(G763), .O(gate261inter8));
  nand2 gate2208(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2209(.a(s_237), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2210(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2211(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2212(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate547(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate548(.a(gate263inter0), .b(s_0), .O(gate263inter1));
  and2  gate549(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate550(.a(s_0), .O(gate263inter3));
  inv1  gate551(.a(s_1), .O(gate263inter4));
  nand2 gate552(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate553(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate554(.a(G766), .O(gate263inter7));
  inv1  gate555(.a(G767), .O(gate263inter8));
  nand2 gate556(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate557(.a(s_1), .b(gate263inter3), .O(gate263inter10));
  nor2  gate558(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate559(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate560(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1065(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1066(.a(gate265inter0), .b(s_74), .O(gate265inter1));
  and2  gate1067(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1068(.a(s_74), .O(gate265inter3));
  inv1  gate1069(.a(s_75), .O(gate265inter4));
  nand2 gate1070(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1071(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1072(.a(G642), .O(gate265inter7));
  inv1  gate1073(.a(G770), .O(gate265inter8));
  nand2 gate1074(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1075(.a(s_75), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1076(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1077(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1078(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2129(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2130(.a(gate271inter0), .b(s_226), .O(gate271inter1));
  and2  gate2131(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2132(.a(s_226), .O(gate271inter3));
  inv1  gate2133(.a(s_227), .O(gate271inter4));
  nand2 gate2134(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2135(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2136(.a(G660), .O(gate271inter7));
  inv1  gate2137(.a(G788), .O(gate271inter8));
  nand2 gate2138(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2139(.a(s_227), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2140(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2141(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2142(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1317(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1318(.a(gate273inter0), .b(s_110), .O(gate273inter1));
  and2  gate1319(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1320(.a(s_110), .O(gate273inter3));
  inv1  gate1321(.a(s_111), .O(gate273inter4));
  nand2 gate1322(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1323(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1324(.a(G642), .O(gate273inter7));
  inv1  gate1325(.a(G794), .O(gate273inter8));
  nand2 gate1326(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1327(.a(s_111), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1328(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1329(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1330(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate883(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate884(.a(gate276inter0), .b(s_48), .O(gate276inter1));
  and2  gate885(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate886(.a(s_48), .O(gate276inter3));
  inv1  gate887(.a(s_49), .O(gate276inter4));
  nand2 gate888(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate889(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate890(.a(G773), .O(gate276inter7));
  inv1  gate891(.a(G797), .O(gate276inter8));
  nand2 gate892(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate893(.a(s_49), .b(gate276inter3), .O(gate276inter10));
  nor2  gate894(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate895(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate896(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1905(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1906(.a(gate278inter0), .b(s_194), .O(gate278inter1));
  and2  gate1907(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1908(.a(s_194), .O(gate278inter3));
  inv1  gate1909(.a(s_195), .O(gate278inter4));
  nand2 gate1910(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1911(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1912(.a(G776), .O(gate278inter7));
  inv1  gate1913(.a(G800), .O(gate278inter8));
  nand2 gate1914(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1915(.a(s_195), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1916(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1917(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1918(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate2241(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2242(.a(gate279inter0), .b(s_242), .O(gate279inter1));
  and2  gate2243(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2244(.a(s_242), .O(gate279inter3));
  inv1  gate2245(.a(s_243), .O(gate279inter4));
  nand2 gate2246(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2247(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2248(.a(G651), .O(gate279inter7));
  inv1  gate2249(.a(G803), .O(gate279inter8));
  nand2 gate2250(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2251(.a(s_243), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2252(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2253(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2254(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate2283(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2284(.a(gate280inter0), .b(s_248), .O(gate280inter1));
  and2  gate2285(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2286(.a(s_248), .O(gate280inter3));
  inv1  gate2287(.a(s_249), .O(gate280inter4));
  nand2 gate2288(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2289(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2290(.a(G779), .O(gate280inter7));
  inv1  gate2291(.a(G803), .O(gate280inter8));
  nand2 gate2292(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2293(.a(s_249), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2294(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2295(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2296(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1961(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1962(.a(gate284inter0), .b(s_202), .O(gate284inter1));
  and2  gate1963(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1964(.a(s_202), .O(gate284inter3));
  inv1  gate1965(.a(s_203), .O(gate284inter4));
  nand2 gate1966(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1967(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1968(.a(G785), .O(gate284inter7));
  inv1  gate1969(.a(G809), .O(gate284inter8));
  nand2 gate1970(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1971(.a(s_203), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1972(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1973(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1974(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate575(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate576(.a(gate286inter0), .b(s_4), .O(gate286inter1));
  and2  gate577(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate578(.a(s_4), .O(gate286inter3));
  inv1  gate579(.a(s_5), .O(gate286inter4));
  nand2 gate580(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate581(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate582(.a(G788), .O(gate286inter7));
  inv1  gate583(.a(G812), .O(gate286inter8));
  nand2 gate584(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate585(.a(s_5), .b(gate286inter3), .O(gate286inter10));
  nor2  gate586(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate587(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate588(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1681(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1682(.a(gate287inter0), .b(s_162), .O(gate287inter1));
  and2  gate1683(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1684(.a(s_162), .O(gate287inter3));
  inv1  gate1685(.a(s_163), .O(gate287inter4));
  nand2 gate1686(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1687(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1688(.a(G663), .O(gate287inter7));
  inv1  gate1689(.a(G815), .O(gate287inter8));
  nand2 gate1690(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1691(.a(s_163), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1692(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1693(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1694(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2451(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2452(.a(gate289inter0), .b(s_272), .O(gate289inter1));
  and2  gate2453(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2454(.a(s_272), .O(gate289inter3));
  inv1  gate2455(.a(s_273), .O(gate289inter4));
  nand2 gate2456(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2457(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2458(.a(G818), .O(gate289inter7));
  inv1  gate2459(.a(G819), .O(gate289inter8));
  nand2 gate2460(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2461(.a(s_273), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2462(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2463(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2464(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate2255(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2256(.a(gate290inter0), .b(s_244), .O(gate290inter1));
  and2  gate2257(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2258(.a(s_244), .O(gate290inter3));
  inv1  gate2259(.a(s_245), .O(gate290inter4));
  nand2 gate2260(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2261(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2262(.a(G820), .O(gate290inter7));
  inv1  gate2263(.a(G821), .O(gate290inter8));
  nand2 gate2264(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2265(.a(s_245), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2266(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2267(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2268(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1373(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1374(.a(gate296inter0), .b(s_118), .O(gate296inter1));
  and2  gate1375(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1376(.a(s_118), .O(gate296inter3));
  inv1  gate1377(.a(s_119), .O(gate296inter4));
  nand2 gate1378(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1379(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1380(.a(G826), .O(gate296inter7));
  inv1  gate1381(.a(G827), .O(gate296inter8));
  nand2 gate1382(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1383(.a(s_119), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1384(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1385(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1386(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2045(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2046(.a(gate394inter0), .b(s_214), .O(gate394inter1));
  and2  gate2047(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2048(.a(s_214), .O(gate394inter3));
  inv1  gate2049(.a(s_215), .O(gate394inter4));
  nand2 gate2050(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2051(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2052(.a(G8), .O(gate394inter7));
  inv1  gate2053(.a(G1057), .O(gate394inter8));
  nand2 gate2054(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2055(.a(s_215), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2056(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2057(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2058(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1023(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1024(.a(gate397inter0), .b(s_68), .O(gate397inter1));
  and2  gate1025(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1026(.a(s_68), .O(gate397inter3));
  inv1  gate1027(.a(s_69), .O(gate397inter4));
  nand2 gate1028(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1029(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1030(.a(G11), .O(gate397inter7));
  inv1  gate1031(.a(G1066), .O(gate397inter8));
  nand2 gate1032(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1033(.a(s_69), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1034(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1035(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1036(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1723(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1724(.a(gate400inter0), .b(s_168), .O(gate400inter1));
  and2  gate1725(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1726(.a(s_168), .O(gate400inter3));
  inv1  gate1727(.a(s_169), .O(gate400inter4));
  nand2 gate1728(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1729(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1730(.a(G14), .O(gate400inter7));
  inv1  gate1731(.a(G1075), .O(gate400inter8));
  nand2 gate1732(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1733(.a(s_169), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1734(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1735(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1736(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1471(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1472(.a(gate401inter0), .b(s_132), .O(gate401inter1));
  and2  gate1473(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1474(.a(s_132), .O(gate401inter3));
  inv1  gate1475(.a(s_133), .O(gate401inter4));
  nand2 gate1476(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1477(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1478(.a(G15), .O(gate401inter7));
  inv1  gate1479(.a(G1078), .O(gate401inter8));
  nand2 gate1480(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1481(.a(s_133), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1482(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1483(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1484(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1107(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1108(.a(gate405inter0), .b(s_80), .O(gate405inter1));
  and2  gate1109(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1110(.a(s_80), .O(gate405inter3));
  inv1  gate1111(.a(s_81), .O(gate405inter4));
  nand2 gate1112(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1113(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1114(.a(G19), .O(gate405inter7));
  inv1  gate1115(.a(G1090), .O(gate405inter8));
  nand2 gate1116(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1117(.a(s_81), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1118(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1119(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1120(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate855(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate856(.a(gate406inter0), .b(s_44), .O(gate406inter1));
  and2  gate857(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate858(.a(s_44), .O(gate406inter3));
  inv1  gate859(.a(s_45), .O(gate406inter4));
  nand2 gate860(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate861(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate862(.a(G20), .O(gate406inter7));
  inv1  gate863(.a(G1093), .O(gate406inter8));
  nand2 gate864(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate865(.a(s_45), .b(gate406inter3), .O(gate406inter10));
  nor2  gate866(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate867(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate868(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1807(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1808(.a(gate407inter0), .b(s_180), .O(gate407inter1));
  and2  gate1809(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1810(.a(s_180), .O(gate407inter3));
  inv1  gate1811(.a(s_181), .O(gate407inter4));
  nand2 gate1812(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1813(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1814(.a(G21), .O(gate407inter7));
  inv1  gate1815(.a(G1096), .O(gate407inter8));
  nand2 gate1816(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1817(.a(s_181), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1818(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1819(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1820(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate939(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate940(.a(gate411inter0), .b(s_56), .O(gate411inter1));
  and2  gate941(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate942(.a(s_56), .O(gate411inter3));
  inv1  gate943(.a(s_57), .O(gate411inter4));
  nand2 gate944(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate945(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate946(.a(G25), .O(gate411inter7));
  inv1  gate947(.a(G1108), .O(gate411inter8));
  nand2 gate948(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate949(.a(s_57), .b(gate411inter3), .O(gate411inter10));
  nor2  gate950(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate951(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate952(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1037(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1038(.a(gate413inter0), .b(s_70), .O(gate413inter1));
  and2  gate1039(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1040(.a(s_70), .O(gate413inter3));
  inv1  gate1041(.a(s_71), .O(gate413inter4));
  nand2 gate1042(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1043(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1044(.a(G27), .O(gate413inter7));
  inv1  gate1045(.a(G1114), .O(gate413inter8));
  nand2 gate1046(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1047(.a(s_71), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1048(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1049(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1050(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1499(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1500(.a(gate418inter0), .b(s_136), .O(gate418inter1));
  and2  gate1501(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1502(.a(s_136), .O(gate418inter3));
  inv1  gate1503(.a(s_137), .O(gate418inter4));
  nand2 gate1504(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1505(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1506(.a(G32), .O(gate418inter7));
  inv1  gate1507(.a(G1129), .O(gate418inter8));
  nand2 gate1508(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1509(.a(s_137), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1510(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1511(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1512(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2031(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2032(.a(gate421inter0), .b(s_212), .O(gate421inter1));
  and2  gate2033(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2034(.a(s_212), .O(gate421inter3));
  inv1  gate2035(.a(s_213), .O(gate421inter4));
  nand2 gate2036(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2037(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2038(.a(G2), .O(gate421inter7));
  inv1  gate2039(.a(G1135), .O(gate421inter8));
  nand2 gate2040(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2041(.a(s_213), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2042(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2043(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2044(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1569(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1570(.a(gate427inter0), .b(s_146), .O(gate427inter1));
  and2  gate1571(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1572(.a(s_146), .O(gate427inter3));
  inv1  gate1573(.a(s_147), .O(gate427inter4));
  nand2 gate1574(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1575(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1576(.a(G5), .O(gate427inter7));
  inv1  gate1577(.a(G1144), .O(gate427inter8));
  nand2 gate1578(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1579(.a(s_147), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1580(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1581(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1582(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1009(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1010(.a(gate429inter0), .b(s_66), .O(gate429inter1));
  and2  gate1011(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1012(.a(s_66), .O(gate429inter3));
  inv1  gate1013(.a(s_67), .O(gate429inter4));
  nand2 gate1014(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1015(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1016(.a(G6), .O(gate429inter7));
  inv1  gate1017(.a(G1147), .O(gate429inter8));
  nand2 gate1018(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1019(.a(s_67), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1020(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1021(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1022(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1177(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1178(.a(gate431inter0), .b(s_90), .O(gate431inter1));
  and2  gate1179(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1180(.a(s_90), .O(gate431inter3));
  inv1  gate1181(.a(s_91), .O(gate431inter4));
  nand2 gate1182(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1183(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1184(.a(G7), .O(gate431inter7));
  inv1  gate1185(.a(G1150), .O(gate431inter8));
  nand2 gate1186(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1187(.a(s_91), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1188(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1189(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1190(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate659(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate660(.a(gate432inter0), .b(s_16), .O(gate432inter1));
  and2  gate661(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate662(.a(s_16), .O(gate432inter3));
  inv1  gate663(.a(s_17), .O(gate432inter4));
  nand2 gate664(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate665(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate666(.a(G1054), .O(gate432inter7));
  inv1  gate667(.a(G1150), .O(gate432inter8));
  nand2 gate668(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate669(.a(s_17), .b(gate432inter3), .O(gate432inter10));
  nor2  gate670(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate671(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate672(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate799(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate800(.a(gate439inter0), .b(s_36), .O(gate439inter1));
  and2  gate801(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate802(.a(s_36), .O(gate439inter3));
  inv1  gate803(.a(s_37), .O(gate439inter4));
  nand2 gate804(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate805(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate806(.a(G11), .O(gate439inter7));
  inv1  gate807(.a(G1162), .O(gate439inter8));
  nand2 gate808(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate809(.a(s_37), .b(gate439inter3), .O(gate439inter10));
  nor2  gate810(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate811(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate812(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1219(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1220(.a(gate442inter0), .b(s_96), .O(gate442inter1));
  and2  gate1221(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1222(.a(s_96), .O(gate442inter3));
  inv1  gate1223(.a(s_97), .O(gate442inter4));
  nand2 gate1224(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1225(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1226(.a(G1069), .O(gate442inter7));
  inv1  gate1227(.a(G1165), .O(gate442inter8));
  nand2 gate1228(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1229(.a(s_97), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1230(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1231(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1232(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1667(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1668(.a(gate446inter0), .b(s_160), .O(gate446inter1));
  and2  gate1669(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1670(.a(s_160), .O(gate446inter3));
  inv1  gate1671(.a(s_161), .O(gate446inter4));
  nand2 gate1672(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1673(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1674(.a(G1075), .O(gate446inter7));
  inv1  gate1675(.a(G1171), .O(gate446inter8));
  nand2 gate1676(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1677(.a(s_161), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1678(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1679(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1680(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate617(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate618(.a(gate447inter0), .b(s_10), .O(gate447inter1));
  and2  gate619(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate620(.a(s_10), .O(gate447inter3));
  inv1  gate621(.a(s_11), .O(gate447inter4));
  nand2 gate622(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate623(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate624(.a(G15), .O(gate447inter7));
  inv1  gate625(.a(G1174), .O(gate447inter8));
  nand2 gate626(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate627(.a(s_11), .b(gate447inter3), .O(gate447inter10));
  nor2  gate628(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate629(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate630(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate2003(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2004(.a(gate449inter0), .b(s_208), .O(gate449inter1));
  and2  gate2005(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2006(.a(s_208), .O(gate449inter3));
  inv1  gate2007(.a(s_209), .O(gate449inter4));
  nand2 gate2008(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2009(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2010(.a(G16), .O(gate449inter7));
  inv1  gate2011(.a(G1177), .O(gate449inter8));
  nand2 gate2012(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2013(.a(s_209), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2014(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2015(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2016(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1457(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1458(.a(gate450inter0), .b(s_130), .O(gate450inter1));
  and2  gate1459(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1460(.a(s_130), .O(gate450inter3));
  inv1  gate1461(.a(s_131), .O(gate450inter4));
  nand2 gate1462(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1463(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1464(.a(G1081), .O(gate450inter7));
  inv1  gate1465(.a(G1177), .O(gate450inter8));
  nand2 gate1466(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1467(.a(s_131), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1468(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1469(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1470(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1947(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1948(.a(gate452inter0), .b(s_200), .O(gate452inter1));
  and2  gate1949(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1950(.a(s_200), .O(gate452inter3));
  inv1  gate1951(.a(s_201), .O(gate452inter4));
  nand2 gate1952(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1953(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1954(.a(G1084), .O(gate452inter7));
  inv1  gate1955(.a(G1180), .O(gate452inter8));
  nand2 gate1956(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1957(.a(s_201), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1958(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1959(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1960(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate589(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate590(.a(gate463inter0), .b(s_6), .O(gate463inter1));
  and2  gate591(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate592(.a(s_6), .O(gate463inter3));
  inv1  gate593(.a(s_7), .O(gate463inter4));
  nand2 gate594(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate595(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate596(.a(G23), .O(gate463inter7));
  inv1  gate597(.a(G1198), .O(gate463inter8));
  nand2 gate598(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate599(.a(s_7), .b(gate463inter3), .O(gate463inter10));
  nor2  gate600(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate601(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate602(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate645(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate646(.a(gate466inter0), .b(s_14), .O(gate466inter1));
  and2  gate647(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate648(.a(s_14), .O(gate466inter3));
  inv1  gate649(.a(s_15), .O(gate466inter4));
  nand2 gate650(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate651(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate652(.a(G1105), .O(gate466inter7));
  inv1  gate653(.a(G1201), .O(gate466inter8));
  nand2 gate654(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate655(.a(s_15), .b(gate466inter3), .O(gate466inter10));
  nor2  gate656(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate657(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate658(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1345(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1346(.a(gate471inter0), .b(s_114), .O(gate471inter1));
  and2  gate1347(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1348(.a(s_114), .O(gate471inter3));
  inv1  gate1349(.a(s_115), .O(gate471inter4));
  nand2 gate1350(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1351(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1352(.a(G27), .O(gate471inter7));
  inv1  gate1353(.a(G1210), .O(gate471inter8));
  nand2 gate1354(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1355(.a(s_115), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1356(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1357(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1358(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate687(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate688(.a(gate474inter0), .b(s_20), .O(gate474inter1));
  and2  gate689(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate690(.a(s_20), .O(gate474inter3));
  inv1  gate691(.a(s_21), .O(gate474inter4));
  nand2 gate692(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate693(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate694(.a(G1117), .O(gate474inter7));
  inv1  gate695(.a(G1213), .O(gate474inter8));
  nand2 gate696(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate697(.a(s_21), .b(gate474inter3), .O(gate474inter10));
  nor2  gate698(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate699(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate700(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate673(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate674(.a(gate476inter0), .b(s_18), .O(gate476inter1));
  and2  gate675(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate676(.a(s_18), .O(gate476inter3));
  inv1  gate677(.a(s_19), .O(gate476inter4));
  nand2 gate678(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate679(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate680(.a(G1120), .O(gate476inter7));
  inv1  gate681(.a(G1216), .O(gate476inter8));
  nand2 gate682(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate683(.a(s_19), .b(gate476inter3), .O(gate476inter10));
  nor2  gate684(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate685(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate686(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1387(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1388(.a(gate478inter0), .b(s_120), .O(gate478inter1));
  and2  gate1389(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1390(.a(s_120), .O(gate478inter3));
  inv1  gate1391(.a(s_121), .O(gate478inter4));
  nand2 gate1392(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1393(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1394(.a(G1123), .O(gate478inter7));
  inv1  gate1395(.a(G1219), .O(gate478inter8));
  nand2 gate1396(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1397(.a(s_121), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1398(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1399(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1400(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1513(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1514(.a(gate479inter0), .b(s_138), .O(gate479inter1));
  and2  gate1515(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1516(.a(s_138), .O(gate479inter3));
  inv1  gate1517(.a(s_139), .O(gate479inter4));
  nand2 gate1518(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1519(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1520(.a(G31), .O(gate479inter7));
  inv1  gate1521(.a(G1222), .O(gate479inter8));
  nand2 gate1522(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1523(.a(s_139), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1524(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1525(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1526(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate981(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate982(.a(gate493inter0), .b(s_62), .O(gate493inter1));
  and2  gate983(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate984(.a(s_62), .O(gate493inter3));
  inv1  gate985(.a(s_63), .O(gate493inter4));
  nand2 gate986(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate987(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate988(.a(G1248), .O(gate493inter7));
  inv1  gate989(.a(G1249), .O(gate493inter8));
  nand2 gate990(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate991(.a(s_63), .b(gate493inter3), .O(gate493inter10));
  nor2  gate992(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate993(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate994(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate2143(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2144(.a(gate495inter0), .b(s_228), .O(gate495inter1));
  and2  gate2145(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2146(.a(s_228), .O(gate495inter3));
  inv1  gate2147(.a(s_229), .O(gate495inter4));
  nand2 gate2148(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2149(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2150(.a(G1252), .O(gate495inter7));
  inv1  gate2151(.a(G1253), .O(gate495inter8));
  nand2 gate2152(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2153(.a(s_229), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2154(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2155(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2156(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1415(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1416(.a(gate497inter0), .b(s_124), .O(gate497inter1));
  and2  gate1417(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1418(.a(s_124), .O(gate497inter3));
  inv1  gate1419(.a(s_125), .O(gate497inter4));
  nand2 gate1420(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1421(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1422(.a(G1256), .O(gate497inter7));
  inv1  gate1423(.a(G1257), .O(gate497inter8));
  nand2 gate1424(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1425(.a(s_125), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1426(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1427(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1428(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1891(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1892(.a(gate498inter0), .b(s_192), .O(gate498inter1));
  and2  gate1893(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1894(.a(s_192), .O(gate498inter3));
  inv1  gate1895(.a(s_193), .O(gate498inter4));
  nand2 gate1896(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1897(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1898(.a(G1258), .O(gate498inter7));
  inv1  gate1899(.a(G1259), .O(gate498inter8));
  nand2 gate1900(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1901(.a(s_193), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1902(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1903(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1904(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1877(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1878(.a(gate503inter0), .b(s_190), .O(gate503inter1));
  and2  gate1879(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1880(.a(s_190), .O(gate503inter3));
  inv1  gate1881(.a(s_191), .O(gate503inter4));
  nand2 gate1882(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1883(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1884(.a(G1268), .O(gate503inter7));
  inv1  gate1885(.a(G1269), .O(gate503inter8));
  nand2 gate1886(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1887(.a(s_191), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1888(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1889(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1890(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2367(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2368(.a(gate504inter0), .b(s_260), .O(gate504inter1));
  and2  gate2369(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2370(.a(s_260), .O(gate504inter3));
  inv1  gate2371(.a(s_261), .O(gate504inter4));
  nand2 gate2372(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2373(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2374(.a(G1270), .O(gate504inter7));
  inv1  gate2375(.a(G1271), .O(gate504inter8));
  nand2 gate2376(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2377(.a(s_261), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2378(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2379(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2380(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1779(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1780(.a(gate506inter0), .b(s_176), .O(gate506inter1));
  and2  gate1781(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1782(.a(s_176), .O(gate506inter3));
  inv1  gate1783(.a(s_177), .O(gate506inter4));
  nand2 gate1784(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1785(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1786(.a(G1274), .O(gate506inter7));
  inv1  gate1787(.a(G1275), .O(gate506inter8));
  nand2 gate1788(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1789(.a(s_177), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1790(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1791(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1792(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2353(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2354(.a(gate509inter0), .b(s_258), .O(gate509inter1));
  and2  gate2355(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2356(.a(s_258), .O(gate509inter3));
  inv1  gate2357(.a(s_259), .O(gate509inter4));
  nand2 gate2358(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2359(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2360(.a(G1280), .O(gate509inter7));
  inv1  gate2361(.a(G1281), .O(gate509inter8));
  nand2 gate2362(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2363(.a(s_259), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2364(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2365(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2366(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule