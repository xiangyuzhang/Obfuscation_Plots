module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate743(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate744(.a(gate11inter0), .b(s_28), .O(gate11inter1));
  and2  gate745(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate746(.a(s_28), .O(gate11inter3));
  inv1  gate747(.a(s_29), .O(gate11inter4));
  nand2 gate748(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate749(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate750(.a(G5), .O(gate11inter7));
  inv1  gate751(.a(G6), .O(gate11inter8));
  nand2 gate752(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate753(.a(s_29), .b(gate11inter3), .O(gate11inter10));
  nor2  gate754(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate755(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate756(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1303(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1304(.a(gate14inter0), .b(s_108), .O(gate14inter1));
  and2  gate1305(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1306(.a(s_108), .O(gate14inter3));
  inv1  gate1307(.a(s_109), .O(gate14inter4));
  nand2 gate1308(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1309(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1310(.a(G11), .O(gate14inter7));
  inv1  gate1311(.a(G12), .O(gate14inter8));
  nand2 gate1312(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1313(.a(s_109), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1314(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1315(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1316(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate869(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate870(.a(gate15inter0), .b(s_46), .O(gate15inter1));
  and2  gate871(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate872(.a(s_46), .O(gate15inter3));
  inv1  gate873(.a(s_47), .O(gate15inter4));
  nand2 gate874(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate875(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate876(.a(G13), .O(gate15inter7));
  inv1  gate877(.a(G14), .O(gate15inter8));
  nand2 gate878(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate879(.a(s_47), .b(gate15inter3), .O(gate15inter10));
  nor2  gate880(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate881(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate882(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1205(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1206(.a(gate16inter0), .b(s_94), .O(gate16inter1));
  and2  gate1207(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1208(.a(s_94), .O(gate16inter3));
  inv1  gate1209(.a(s_95), .O(gate16inter4));
  nand2 gate1210(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1211(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1212(.a(G15), .O(gate16inter7));
  inv1  gate1213(.a(G16), .O(gate16inter8));
  nand2 gate1214(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1215(.a(s_95), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1216(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1217(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1218(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1191(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1192(.a(gate19inter0), .b(s_92), .O(gate19inter1));
  and2  gate1193(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1194(.a(s_92), .O(gate19inter3));
  inv1  gate1195(.a(s_93), .O(gate19inter4));
  nand2 gate1196(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1197(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1198(.a(G21), .O(gate19inter7));
  inv1  gate1199(.a(G22), .O(gate19inter8));
  nand2 gate1200(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1201(.a(s_93), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1202(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1203(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1204(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1723(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1724(.a(gate23inter0), .b(s_168), .O(gate23inter1));
  and2  gate1725(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1726(.a(s_168), .O(gate23inter3));
  inv1  gate1727(.a(s_169), .O(gate23inter4));
  nand2 gate1728(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1729(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1730(.a(G29), .O(gate23inter7));
  inv1  gate1731(.a(G30), .O(gate23inter8));
  nand2 gate1732(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1733(.a(s_169), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1734(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1735(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1736(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1667(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1668(.a(gate24inter0), .b(s_160), .O(gate24inter1));
  and2  gate1669(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1670(.a(s_160), .O(gate24inter3));
  inv1  gate1671(.a(s_161), .O(gate24inter4));
  nand2 gate1672(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1673(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1674(.a(G31), .O(gate24inter7));
  inv1  gate1675(.a(G32), .O(gate24inter8));
  nand2 gate1676(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1677(.a(s_161), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1678(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1679(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1680(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1695(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1696(.a(gate25inter0), .b(s_164), .O(gate25inter1));
  and2  gate1697(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1698(.a(s_164), .O(gate25inter3));
  inv1  gate1699(.a(s_165), .O(gate25inter4));
  nand2 gate1700(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1701(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1702(.a(G1), .O(gate25inter7));
  inv1  gate1703(.a(G5), .O(gate25inter8));
  nand2 gate1704(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1705(.a(s_165), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1706(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1707(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1708(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1485(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1486(.a(gate27inter0), .b(s_134), .O(gate27inter1));
  and2  gate1487(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1488(.a(s_134), .O(gate27inter3));
  inv1  gate1489(.a(s_135), .O(gate27inter4));
  nand2 gate1490(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1491(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1492(.a(G2), .O(gate27inter7));
  inv1  gate1493(.a(G6), .O(gate27inter8));
  nand2 gate1494(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1495(.a(s_135), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1496(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1497(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1498(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate645(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate646(.a(gate31inter0), .b(s_14), .O(gate31inter1));
  and2  gate647(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate648(.a(s_14), .O(gate31inter3));
  inv1  gate649(.a(s_15), .O(gate31inter4));
  nand2 gate650(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate651(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate652(.a(G4), .O(gate31inter7));
  inv1  gate653(.a(G8), .O(gate31inter8));
  nand2 gate654(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate655(.a(s_15), .b(gate31inter3), .O(gate31inter10));
  nor2  gate656(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate657(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate658(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1905(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1906(.a(gate39inter0), .b(s_194), .O(gate39inter1));
  and2  gate1907(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1908(.a(s_194), .O(gate39inter3));
  inv1  gate1909(.a(s_195), .O(gate39inter4));
  nand2 gate1910(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1911(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1912(.a(G20), .O(gate39inter7));
  inv1  gate1913(.a(G24), .O(gate39inter8));
  nand2 gate1914(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1915(.a(s_195), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1916(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1917(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1918(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate925(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate926(.a(gate41inter0), .b(s_54), .O(gate41inter1));
  and2  gate927(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate928(.a(s_54), .O(gate41inter3));
  inv1  gate929(.a(s_55), .O(gate41inter4));
  nand2 gate930(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate931(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate932(.a(G1), .O(gate41inter7));
  inv1  gate933(.a(G266), .O(gate41inter8));
  nand2 gate934(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate935(.a(s_55), .b(gate41inter3), .O(gate41inter10));
  nor2  gate936(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate937(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate938(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate799(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate800(.a(gate44inter0), .b(s_36), .O(gate44inter1));
  and2  gate801(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate802(.a(s_36), .O(gate44inter3));
  inv1  gate803(.a(s_37), .O(gate44inter4));
  nand2 gate804(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate805(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate806(.a(G4), .O(gate44inter7));
  inv1  gate807(.a(G269), .O(gate44inter8));
  nand2 gate808(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate809(.a(s_37), .b(gate44inter3), .O(gate44inter10));
  nor2  gate810(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate811(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate812(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1877(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1878(.a(gate45inter0), .b(s_190), .O(gate45inter1));
  and2  gate1879(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1880(.a(s_190), .O(gate45inter3));
  inv1  gate1881(.a(s_191), .O(gate45inter4));
  nand2 gate1882(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1883(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1884(.a(G5), .O(gate45inter7));
  inv1  gate1885(.a(G272), .O(gate45inter8));
  nand2 gate1886(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1887(.a(s_191), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1888(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1889(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1890(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1779(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1780(.a(gate51inter0), .b(s_176), .O(gate51inter1));
  and2  gate1781(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1782(.a(s_176), .O(gate51inter3));
  inv1  gate1783(.a(s_177), .O(gate51inter4));
  nand2 gate1784(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1785(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1786(.a(G11), .O(gate51inter7));
  inv1  gate1787(.a(G281), .O(gate51inter8));
  nand2 gate1788(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1789(.a(s_177), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1790(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1791(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1792(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1261(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1262(.a(gate59inter0), .b(s_102), .O(gate59inter1));
  and2  gate1263(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1264(.a(s_102), .O(gate59inter3));
  inv1  gate1265(.a(s_103), .O(gate59inter4));
  nand2 gate1266(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1267(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1268(.a(G19), .O(gate59inter7));
  inv1  gate1269(.a(G293), .O(gate59inter8));
  nand2 gate1270(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1271(.a(s_103), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1272(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1273(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1274(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1247(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1248(.a(gate60inter0), .b(s_100), .O(gate60inter1));
  and2  gate1249(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1250(.a(s_100), .O(gate60inter3));
  inv1  gate1251(.a(s_101), .O(gate60inter4));
  nand2 gate1252(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1253(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1254(.a(G20), .O(gate60inter7));
  inv1  gate1255(.a(G293), .O(gate60inter8));
  nand2 gate1256(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1257(.a(s_101), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1258(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1259(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1260(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1121(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1122(.a(gate70inter0), .b(s_82), .O(gate70inter1));
  and2  gate1123(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1124(.a(s_82), .O(gate70inter3));
  inv1  gate1125(.a(s_83), .O(gate70inter4));
  nand2 gate1126(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1127(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1128(.a(G30), .O(gate70inter7));
  inv1  gate1129(.a(G308), .O(gate70inter8));
  nand2 gate1130(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1131(.a(s_83), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1132(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1133(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1134(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate701(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate702(.a(gate71inter0), .b(s_22), .O(gate71inter1));
  and2  gate703(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate704(.a(s_22), .O(gate71inter3));
  inv1  gate705(.a(s_23), .O(gate71inter4));
  nand2 gate706(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate707(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate708(.a(G31), .O(gate71inter7));
  inv1  gate709(.a(G311), .O(gate71inter8));
  nand2 gate710(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate711(.a(s_23), .b(gate71inter3), .O(gate71inter10));
  nor2  gate712(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate713(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate714(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1765(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1766(.a(gate72inter0), .b(s_174), .O(gate72inter1));
  and2  gate1767(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1768(.a(s_174), .O(gate72inter3));
  inv1  gate1769(.a(s_175), .O(gate72inter4));
  nand2 gate1770(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1771(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1772(.a(G32), .O(gate72inter7));
  inv1  gate1773(.a(G311), .O(gate72inter8));
  nand2 gate1774(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1775(.a(s_175), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1776(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1777(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1778(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1499(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1500(.a(gate78inter0), .b(s_136), .O(gate78inter1));
  and2  gate1501(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1502(.a(s_136), .O(gate78inter3));
  inv1  gate1503(.a(s_137), .O(gate78inter4));
  nand2 gate1504(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1505(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1506(.a(G6), .O(gate78inter7));
  inv1  gate1507(.a(G320), .O(gate78inter8));
  nand2 gate1508(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1509(.a(s_137), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1510(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1511(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1512(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate687(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate688(.a(gate81inter0), .b(s_20), .O(gate81inter1));
  and2  gate689(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate690(.a(s_20), .O(gate81inter3));
  inv1  gate691(.a(s_21), .O(gate81inter4));
  nand2 gate692(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate693(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate694(.a(G3), .O(gate81inter7));
  inv1  gate695(.a(G326), .O(gate81inter8));
  nand2 gate696(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate697(.a(s_21), .b(gate81inter3), .O(gate81inter10));
  nor2  gate698(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate699(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate700(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1653(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1654(.a(gate84inter0), .b(s_158), .O(gate84inter1));
  and2  gate1655(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1656(.a(s_158), .O(gate84inter3));
  inv1  gate1657(.a(s_159), .O(gate84inter4));
  nand2 gate1658(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1659(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1660(.a(G15), .O(gate84inter7));
  inv1  gate1661(.a(G329), .O(gate84inter8));
  nand2 gate1662(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1663(.a(s_159), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1664(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1665(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1666(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate813(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate814(.a(gate85inter0), .b(s_38), .O(gate85inter1));
  and2  gate815(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate816(.a(s_38), .O(gate85inter3));
  inv1  gate817(.a(s_39), .O(gate85inter4));
  nand2 gate818(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate819(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate820(.a(G4), .O(gate85inter7));
  inv1  gate821(.a(G332), .O(gate85inter8));
  nand2 gate822(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate823(.a(s_39), .b(gate85inter3), .O(gate85inter10));
  nor2  gate824(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate825(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate826(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1107(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1108(.a(gate88inter0), .b(s_80), .O(gate88inter1));
  and2  gate1109(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1110(.a(s_80), .O(gate88inter3));
  inv1  gate1111(.a(s_81), .O(gate88inter4));
  nand2 gate1112(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1113(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1114(.a(G16), .O(gate88inter7));
  inv1  gate1115(.a(G335), .O(gate88inter8));
  nand2 gate1116(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1117(.a(s_81), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1118(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1119(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1120(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1527(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1528(.a(gate90inter0), .b(s_140), .O(gate90inter1));
  and2  gate1529(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1530(.a(s_140), .O(gate90inter3));
  inv1  gate1531(.a(s_141), .O(gate90inter4));
  nand2 gate1532(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1533(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1534(.a(G21), .O(gate90inter7));
  inv1  gate1535(.a(G338), .O(gate90inter8));
  nand2 gate1536(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1537(.a(s_141), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1538(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1539(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1540(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate911(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate912(.a(gate96inter0), .b(s_52), .O(gate96inter1));
  and2  gate913(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate914(.a(s_52), .O(gate96inter3));
  inv1  gate915(.a(s_53), .O(gate96inter4));
  nand2 gate916(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate917(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate918(.a(G30), .O(gate96inter7));
  inv1  gate919(.a(G347), .O(gate96inter8));
  nand2 gate920(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate921(.a(s_53), .b(gate96inter3), .O(gate96inter10));
  nor2  gate922(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate923(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate924(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1863(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1864(.a(gate101inter0), .b(s_188), .O(gate101inter1));
  and2  gate1865(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1866(.a(s_188), .O(gate101inter3));
  inv1  gate1867(.a(s_189), .O(gate101inter4));
  nand2 gate1868(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1869(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1870(.a(G20), .O(gate101inter7));
  inv1  gate1871(.a(G356), .O(gate101inter8));
  nand2 gate1872(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1873(.a(s_189), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1874(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1875(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1876(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1933(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1934(.a(gate110inter0), .b(s_198), .O(gate110inter1));
  and2  gate1935(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1936(.a(s_198), .O(gate110inter3));
  inv1  gate1937(.a(s_199), .O(gate110inter4));
  nand2 gate1938(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1939(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1940(.a(G372), .O(gate110inter7));
  inv1  gate1941(.a(G373), .O(gate110inter8));
  nand2 gate1942(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1943(.a(s_199), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1944(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1945(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1946(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate547(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate548(.a(gate120inter0), .b(s_0), .O(gate120inter1));
  and2  gate549(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate550(.a(s_0), .O(gate120inter3));
  inv1  gate551(.a(s_1), .O(gate120inter4));
  nand2 gate552(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate553(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate554(.a(G392), .O(gate120inter7));
  inv1  gate555(.a(G393), .O(gate120inter8));
  nand2 gate556(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate557(.a(s_1), .b(gate120inter3), .O(gate120inter10));
  nor2  gate558(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate559(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate560(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate967(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate968(.a(gate123inter0), .b(s_60), .O(gate123inter1));
  and2  gate969(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate970(.a(s_60), .O(gate123inter3));
  inv1  gate971(.a(s_61), .O(gate123inter4));
  nand2 gate972(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate973(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate974(.a(G398), .O(gate123inter7));
  inv1  gate975(.a(G399), .O(gate123inter8));
  nand2 gate976(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate977(.a(s_61), .b(gate123inter3), .O(gate123inter10));
  nor2  gate978(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate979(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate980(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate659(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate660(.a(gate127inter0), .b(s_16), .O(gate127inter1));
  and2  gate661(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate662(.a(s_16), .O(gate127inter3));
  inv1  gate663(.a(s_17), .O(gate127inter4));
  nand2 gate664(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate665(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate666(.a(G406), .O(gate127inter7));
  inv1  gate667(.a(G407), .O(gate127inter8));
  nand2 gate668(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate669(.a(s_17), .b(gate127inter3), .O(gate127inter10));
  nor2  gate670(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate671(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate672(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate617(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate618(.a(gate129inter0), .b(s_10), .O(gate129inter1));
  and2  gate619(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate620(.a(s_10), .O(gate129inter3));
  inv1  gate621(.a(s_11), .O(gate129inter4));
  nand2 gate622(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate623(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate624(.a(G410), .O(gate129inter7));
  inv1  gate625(.a(G411), .O(gate129inter8));
  nand2 gate626(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate627(.a(s_11), .b(gate129inter3), .O(gate129inter10));
  nor2  gate628(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate629(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate630(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate589(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate590(.a(gate138inter0), .b(s_6), .O(gate138inter1));
  and2  gate591(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate592(.a(s_6), .O(gate138inter3));
  inv1  gate593(.a(s_7), .O(gate138inter4));
  nand2 gate594(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate595(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate596(.a(G432), .O(gate138inter7));
  inv1  gate597(.a(G435), .O(gate138inter8));
  nand2 gate598(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate599(.a(s_7), .b(gate138inter3), .O(gate138inter10));
  nor2  gate600(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate601(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate602(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1737(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1738(.a(gate139inter0), .b(s_170), .O(gate139inter1));
  and2  gate1739(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1740(.a(s_170), .O(gate139inter3));
  inv1  gate1741(.a(s_171), .O(gate139inter4));
  nand2 gate1742(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1743(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1744(.a(G438), .O(gate139inter7));
  inv1  gate1745(.a(G441), .O(gate139inter8));
  nand2 gate1746(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1747(.a(s_171), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1748(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1749(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1750(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1093(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1094(.a(gate141inter0), .b(s_78), .O(gate141inter1));
  and2  gate1095(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1096(.a(s_78), .O(gate141inter3));
  inv1  gate1097(.a(s_79), .O(gate141inter4));
  nand2 gate1098(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1099(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1100(.a(G450), .O(gate141inter7));
  inv1  gate1101(.a(G453), .O(gate141inter8));
  nand2 gate1102(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1103(.a(s_79), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1104(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1105(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1106(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1163(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1164(.a(gate145inter0), .b(s_88), .O(gate145inter1));
  and2  gate1165(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1166(.a(s_88), .O(gate145inter3));
  inv1  gate1167(.a(s_89), .O(gate145inter4));
  nand2 gate1168(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1169(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1170(.a(G474), .O(gate145inter7));
  inv1  gate1171(.a(G477), .O(gate145inter8));
  nand2 gate1172(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1173(.a(s_89), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1174(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1175(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1176(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate883(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate884(.a(gate146inter0), .b(s_48), .O(gate146inter1));
  and2  gate885(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate886(.a(s_48), .O(gate146inter3));
  inv1  gate887(.a(s_49), .O(gate146inter4));
  nand2 gate888(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate889(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate890(.a(G480), .O(gate146inter7));
  inv1  gate891(.a(G483), .O(gate146inter8));
  nand2 gate892(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate893(.a(s_49), .b(gate146inter3), .O(gate146inter10));
  nor2  gate894(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate895(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate896(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1597(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1598(.a(gate147inter0), .b(s_150), .O(gate147inter1));
  and2  gate1599(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1600(.a(s_150), .O(gate147inter3));
  inv1  gate1601(.a(s_151), .O(gate147inter4));
  nand2 gate1602(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1603(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1604(.a(G486), .O(gate147inter7));
  inv1  gate1605(.a(G489), .O(gate147inter8));
  nand2 gate1606(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1607(.a(s_151), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1608(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1609(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1610(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1079(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1080(.a(gate165inter0), .b(s_76), .O(gate165inter1));
  and2  gate1081(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1082(.a(s_76), .O(gate165inter3));
  inv1  gate1083(.a(s_77), .O(gate165inter4));
  nand2 gate1084(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1085(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1086(.a(G462), .O(gate165inter7));
  inv1  gate1087(.a(G540), .O(gate165inter8));
  nand2 gate1088(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1089(.a(s_77), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1090(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1091(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1092(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1457(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1458(.a(gate166inter0), .b(s_130), .O(gate166inter1));
  and2  gate1459(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1460(.a(s_130), .O(gate166inter3));
  inv1  gate1461(.a(s_131), .O(gate166inter4));
  nand2 gate1462(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1463(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1464(.a(G465), .O(gate166inter7));
  inv1  gate1465(.a(G540), .O(gate166inter8));
  nand2 gate1466(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1467(.a(s_131), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1468(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1469(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1470(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1387(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1388(.a(gate185inter0), .b(s_120), .O(gate185inter1));
  and2  gate1389(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1390(.a(s_120), .O(gate185inter3));
  inv1  gate1391(.a(s_121), .O(gate185inter4));
  nand2 gate1392(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1393(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1394(.a(G570), .O(gate185inter7));
  inv1  gate1395(.a(G571), .O(gate185inter8));
  nand2 gate1396(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1397(.a(s_121), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1398(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1399(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1400(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1611(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1612(.a(gate190inter0), .b(s_152), .O(gate190inter1));
  and2  gate1613(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1614(.a(s_152), .O(gate190inter3));
  inv1  gate1615(.a(s_153), .O(gate190inter4));
  nand2 gate1616(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1617(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1618(.a(G580), .O(gate190inter7));
  inv1  gate1619(.a(G581), .O(gate190inter8));
  nand2 gate1620(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1621(.a(s_153), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1622(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1623(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1624(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1415(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1416(.a(gate191inter0), .b(s_124), .O(gate191inter1));
  and2  gate1417(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1418(.a(s_124), .O(gate191inter3));
  inv1  gate1419(.a(s_125), .O(gate191inter4));
  nand2 gate1420(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1421(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1422(.a(G582), .O(gate191inter7));
  inv1  gate1423(.a(G583), .O(gate191inter8));
  nand2 gate1424(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1425(.a(s_125), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1426(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1427(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1428(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1947(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1948(.a(gate197inter0), .b(s_200), .O(gate197inter1));
  and2  gate1949(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1950(.a(s_200), .O(gate197inter3));
  inv1  gate1951(.a(s_201), .O(gate197inter4));
  nand2 gate1952(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1953(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1954(.a(G594), .O(gate197inter7));
  inv1  gate1955(.a(G595), .O(gate197inter8));
  nand2 gate1956(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1957(.a(s_201), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1958(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1959(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1960(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate715(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate716(.a(gate208inter0), .b(s_24), .O(gate208inter1));
  and2  gate717(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate718(.a(s_24), .O(gate208inter3));
  inv1  gate719(.a(s_25), .O(gate208inter4));
  nand2 gate720(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate721(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate722(.a(G627), .O(gate208inter7));
  inv1  gate723(.a(G637), .O(gate208inter8));
  nand2 gate724(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate725(.a(s_25), .b(gate208inter3), .O(gate208inter10));
  nor2  gate726(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate727(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate728(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1891(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1892(.a(gate222inter0), .b(s_192), .O(gate222inter1));
  and2  gate1893(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1894(.a(s_192), .O(gate222inter3));
  inv1  gate1895(.a(s_193), .O(gate222inter4));
  nand2 gate1896(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1897(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1898(.a(G632), .O(gate222inter7));
  inv1  gate1899(.a(G684), .O(gate222inter8));
  nand2 gate1900(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1901(.a(s_193), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1902(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1903(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1904(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1233(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1234(.a(gate227inter0), .b(s_98), .O(gate227inter1));
  and2  gate1235(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1236(.a(s_98), .O(gate227inter3));
  inv1  gate1237(.a(s_99), .O(gate227inter4));
  nand2 gate1238(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1239(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1240(.a(G694), .O(gate227inter7));
  inv1  gate1241(.a(G695), .O(gate227inter8));
  nand2 gate1242(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1243(.a(s_99), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1244(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1245(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1246(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1835(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1836(.a(gate230inter0), .b(s_184), .O(gate230inter1));
  and2  gate1837(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1838(.a(s_184), .O(gate230inter3));
  inv1  gate1839(.a(s_185), .O(gate230inter4));
  nand2 gate1840(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1841(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1842(.a(G700), .O(gate230inter7));
  inv1  gate1843(.a(G701), .O(gate230inter8));
  nand2 gate1844(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1845(.a(s_185), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1846(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1847(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1848(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate827(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate828(.a(gate233inter0), .b(s_40), .O(gate233inter1));
  and2  gate829(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate830(.a(s_40), .O(gate233inter3));
  inv1  gate831(.a(s_41), .O(gate233inter4));
  nand2 gate832(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate833(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate834(.a(G242), .O(gate233inter7));
  inv1  gate835(.a(G718), .O(gate233inter8));
  nand2 gate836(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate837(.a(s_41), .b(gate233inter3), .O(gate233inter10));
  nor2  gate838(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate839(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate840(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1541(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1542(.a(gate234inter0), .b(s_142), .O(gate234inter1));
  and2  gate1543(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1544(.a(s_142), .O(gate234inter3));
  inv1  gate1545(.a(s_143), .O(gate234inter4));
  nand2 gate1546(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1547(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1548(.a(G245), .O(gate234inter7));
  inv1  gate1549(.a(G721), .O(gate234inter8));
  nand2 gate1550(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1551(.a(s_143), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1552(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1553(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1554(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate561(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate562(.a(gate238inter0), .b(s_2), .O(gate238inter1));
  and2  gate563(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate564(.a(s_2), .O(gate238inter3));
  inv1  gate565(.a(s_3), .O(gate238inter4));
  nand2 gate566(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate567(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate568(.a(G257), .O(gate238inter7));
  inv1  gate569(.a(G709), .O(gate238inter8));
  nand2 gate570(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate571(.a(s_3), .b(gate238inter3), .O(gate238inter10));
  nor2  gate572(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate573(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate574(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1709(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1710(.a(gate249inter0), .b(s_166), .O(gate249inter1));
  and2  gate1711(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1712(.a(s_166), .O(gate249inter3));
  inv1  gate1713(.a(s_167), .O(gate249inter4));
  nand2 gate1714(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1715(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1716(.a(G254), .O(gate249inter7));
  inv1  gate1717(.a(G742), .O(gate249inter8));
  nand2 gate1718(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1719(.a(s_167), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1720(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1721(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1722(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate939(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate940(.a(gate251inter0), .b(s_56), .O(gate251inter1));
  and2  gate941(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate942(.a(s_56), .O(gate251inter3));
  inv1  gate943(.a(s_57), .O(gate251inter4));
  nand2 gate944(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate945(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate946(.a(G257), .O(gate251inter7));
  inv1  gate947(.a(G745), .O(gate251inter8));
  nand2 gate948(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate949(.a(s_57), .b(gate251inter3), .O(gate251inter10));
  nor2  gate950(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate951(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate952(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1513(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1514(.a(gate254inter0), .b(s_138), .O(gate254inter1));
  and2  gate1515(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1516(.a(s_138), .O(gate254inter3));
  inv1  gate1517(.a(s_139), .O(gate254inter4));
  nand2 gate1518(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1519(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1520(.a(G712), .O(gate254inter7));
  inv1  gate1521(.a(G748), .O(gate254inter8));
  nand2 gate1522(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1523(.a(s_139), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1524(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1525(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1526(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1821(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1822(.a(gate258inter0), .b(s_182), .O(gate258inter1));
  and2  gate1823(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1824(.a(s_182), .O(gate258inter3));
  inv1  gate1825(.a(s_183), .O(gate258inter4));
  nand2 gate1826(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1827(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1828(.a(G756), .O(gate258inter7));
  inv1  gate1829(.a(G757), .O(gate258inter8));
  nand2 gate1830(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1831(.a(s_183), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1832(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1833(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1834(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1471(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1472(.a(gate261inter0), .b(s_132), .O(gate261inter1));
  and2  gate1473(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1474(.a(s_132), .O(gate261inter3));
  inv1  gate1475(.a(s_133), .O(gate261inter4));
  nand2 gate1476(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1477(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1478(.a(G762), .O(gate261inter7));
  inv1  gate1479(.a(G763), .O(gate261inter8));
  nand2 gate1480(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1481(.a(s_133), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1482(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1483(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1484(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1807(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1808(.a(gate266inter0), .b(s_180), .O(gate266inter1));
  and2  gate1809(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1810(.a(s_180), .O(gate266inter3));
  inv1  gate1811(.a(s_181), .O(gate266inter4));
  nand2 gate1812(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1813(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1814(.a(G645), .O(gate266inter7));
  inv1  gate1815(.a(G773), .O(gate266inter8));
  nand2 gate1816(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1817(.a(s_181), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1818(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1819(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1820(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1583(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1584(.a(gate269inter0), .b(s_148), .O(gate269inter1));
  and2  gate1585(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1586(.a(s_148), .O(gate269inter3));
  inv1  gate1587(.a(s_149), .O(gate269inter4));
  nand2 gate1588(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1589(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1590(.a(G654), .O(gate269inter7));
  inv1  gate1591(.a(G782), .O(gate269inter8));
  nand2 gate1592(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1593(.a(s_149), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1594(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1595(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1596(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1849(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1850(.a(gate276inter0), .b(s_186), .O(gate276inter1));
  and2  gate1851(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1852(.a(s_186), .O(gate276inter3));
  inv1  gate1853(.a(s_187), .O(gate276inter4));
  nand2 gate1854(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1855(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1856(.a(G773), .O(gate276inter7));
  inv1  gate1857(.a(G797), .O(gate276inter8));
  nand2 gate1858(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1859(.a(s_187), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1860(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1861(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1862(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1429(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1430(.a(gate277inter0), .b(s_126), .O(gate277inter1));
  and2  gate1431(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1432(.a(s_126), .O(gate277inter3));
  inv1  gate1433(.a(s_127), .O(gate277inter4));
  nand2 gate1434(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1435(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1436(.a(G648), .O(gate277inter7));
  inv1  gate1437(.a(G800), .O(gate277inter8));
  nand2 gate1438(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1439(.a(s_127), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1440(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1441(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1442(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate897(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate898(.a(gate285inter0), .b(s_50), .O(gate285inter1));
  and2  gate899(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate900(.a(s_50), .O(gate285inter3));
  inv1  gate901(.a(s_51), .O(gate285inter4));
  nand2 gate902(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate903(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate904(.a(G660), .O(gate285inter7));
  inv1  gate905(.a(G812), .O(gate285inter8));
  nand2 gate906(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate907(.a(s_51), .b(gate285inter3), .O(gate285inter10));
  nor2  gate908(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate909(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate910(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1051(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1052(.a(gate287inter0), .b(s_72), .O(gate287inter1));
  and2  gate1053(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1054(.a(s_72), .O(gate287inter3));
  inv1  gate1055(.a(s_73), .O(gate287inter4));
  nand2 gate1056(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1057(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1058(.a(G663), .O(gate287inter7));
  inv1  gate1059(.a(G815), .O(gate287inter8));
  nand2 gate1060(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1061(.a(s_73), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1062(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1063(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1064(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1009(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1010(.a(gate290inter0), .b(s_66), .O(gate290inter1));
  and2  gate1011(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1012(.a(s_66), .O(gate290inter3));
  inv1  gate1013(.a(s_67), .O(gate290inter4));
  nand2 gate1014(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1015(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1016(.a(G820), .O(gate290inter7));
  inv1  gate1017(.a(G821), .O(gate290inter8));
  nand2 gate1018(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1019(.a(s_67), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1020(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1021(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1022(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1289(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1290(.a(gate291inter0), .b(s_106), .O(gate291inter1));
  and2  gate1291(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1292(.a(s_106), .O(gate291inter3));
  inv1  gate1293(.a(s_107), .O(gate291inter4));
  nand2 gate1294(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1295(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1296(.a(G822), .O(gate291inter7));
  inv1  gate1297(.a(G823), .O(gate291inter8));
  nand2 gate1298(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1299(.a(s_107), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1300(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1301(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1302(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate841(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate842(.a(gate293inter0), .b(s_42), .O(gate293inter1));
  and2  gate843(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate844(.a(s_42), .O(gate293inter3));
  inv1  gate845(.a(s_43), .O(gate293inter4));
  nand2 gate846(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate847(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate848(.a(G828), .O(gate293inter7));
  inv1  gate849(.a(G829), .O(gate293inter8));
  nand2 gate850(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate851(.a(s_43), .b(gate293inter3), .O(gate293inter10));
  nor2  gate852(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate853(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate854(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1149(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1150(.a(gate294inter0), .b(s_86), .O(gate294inter1));
  and2  gate1151(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1152(.a(s_86), .O(gate294inter3));
  inv1  gate1153(.a(s_87), .O(gate294inter4));
  nand2 gate1154(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1155(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1156(.a(G832), .O(gate294inter7));
  inv1  gate1157(.a(G833), .O(gate294inter8));
  nand2 gate1158(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1159(.a(s_87), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1160(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1161(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1162(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1023(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1024(.a(gate389inter0), .b(s_68), .O(gate389inter1));
  and2  gate1025(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1026(.a(s_68), .O(gate389inter3));
  inv1  gate1027(.a(s_69), .O(gate389inter4));
  nand2 gate1028(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1029(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1030(.a(G3), .O(gate389inter7));
  inv1  gate1031(.a(G1042), .O(gate389inter8));
  nand2 gate1032(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1033(.a(s_69), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1034(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1035(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1036(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1569(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1570(.a(gate392inter0), .b(s_146), .O(gate392inter1));
  and2  gate1571(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1572(.a(s_146), .O(gate392inter3));
  inv1  gate1573(.a(s_147), .O(gate392inter4));
  nand2 gate1574(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1575(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1576(.a(G6), .O(gate392inter7));
  inv1  gate1577(.a(G1051), .O(gate392inter8));
  nand2 gate1578(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1579(.a(s_147), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1580(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1581(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1582(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1681(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1682(.a(gate393inter0), .b(s_162), .O(gate393inter1));
  and2  gate1683(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1684(.a(s_162), .O(gate393inter3));
  inv1  gate1685(.a(s_163), .O(gate393inter4));
  nand2 gate1686(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1687(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1688(.a(G7), .O(gate393inter7));
  inv1  gate1689(.a(G1054), .O(gate393inter8));
  nand2 gate1690(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1691(.a(s_163), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1692(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1693(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1694(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1317(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1318(.a(gate395inter0), .b(s_110), .O(gate395inter1));
  and2  gate1319(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1320(.a(s_110), .O(gate395inter3));
  inv1  gate1321(.a(s_111), .O(gate395inter4));
  nand2 gate1322(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1323(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1324(.a(G9), .O(gate395inter7));
  inv1  gate1325(.a(G1060), .O(gate395inter8));
  nand2 gate1326(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1327(.a(s_111), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1328(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1329(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1330(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1793(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1794(.a(gate399inter0), .b(s_178), .O(gate399inter1));
  and2  gate1795(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1796(.a(s_178), .O(gate399inter3));
  inv1  gate1797(.a(s_179), .O(gate399inter4));
  nand2 gate1798(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1799(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1800(.a(G13), .O(gate399inter7));
  inv1  gate1801(.a(G1072), .O(gate399inter8));
  nand2 gate1802(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1803(.a(s_179), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1804(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1805(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1806(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate673(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate674(.a(gate405inter0), .b(s_18), .O(gate405inter1));
  and2  gate675(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate676(.a(s_18), .O(gate405inter3));
  inv1  gate677(.a(s_19), .O(gate405inter4));
  nand2 gate678(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate679(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate680(.a(G19), .O(gate405inter7));
  inv1  gate681(.a(G1090), .O(gate405inter8));
  nand2 gate682(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate683(.a(s_19), .b(gate405inter3), .O(gate405inter10));
  nor2  gate684(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate685(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate686(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate631(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate632(.a(gate411inter0), .b(s_12), .O(gate411inter1));
  and2  gate633(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate634(.a(s_12), .O(gate411inter3));
  inv1  gate635(.a(s_13), .O(gate411inter4));
  nand2 gate636(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate637(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate638(.a(G25), .O(gate411inter7));
  inv1  gate639(.a(G1108), .O(gate411inter8));
  nand2 gate640(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate641(.a(s_13), .b(gate411inter3), .O(gate411inter10));
  nor2  gate642(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate643(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate644(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1373(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1374(.a(gate413inter0), .b(s_118), .O(gate413inter1));
  and2  gate1375(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1376(.a(s_118), .O(gate413inter3));
  inv1  gate1377(.a(s_119), .O(gate413inter4));
  nand2 gate1378(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1379(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1380(.a(G27), .O(gate413inter7));
  inv1  gate1381(.a(G1114), .O(gate413inter8));
  nand2 gate1382(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1383(.a(s_119), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1384(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1385(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1386(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1359(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1360(.a(gate414inter0), .b(s_116), .O(gate414inter1));
  and2  gate1361(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1362(.a(s_116), .O(gate414inter3));
  inv1  gate1363(.a(s_117), .O(gate414inter4));
  nand2 gate1364(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1365(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1366(.a(G28), .O(gate414inter7));
  inv1  gate1367(.a(G1117), .O(gate414inter8));
  nand2 gate1368(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1369(.a(s_117), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1370(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1371(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1372(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1275(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1276(.a(gate416inter0), .b(s_104), .O(gate416inter1));
  and2  gate1277(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1278(.a(s_104), .O(gate416inter3));
  inv1  gate1279(.a(s_105), .O(gate416inter4));
  nand2 gate1280(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1281(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1282(.a(G30), .O(gate416inter7));
  inv1  gate1283(.a(G1123), .O(gate416inter8));
  nand2 gate1284(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1285(.a(s_105), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1286(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1287(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1288(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate995(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate996(.a(gate418inter0), .b(s_64), .O(gate418inter1));
  and2  gate997(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate998(.a(s_64), .O(gate418inter3));
  inv1  gate999(.a(s_65), .O(gate418inter4));
  nand2 gate1000(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1001(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1002(.a(G32), .O(gate418inter7));
  inv1  gate1003(.a(G1129), .O(gate418inter8));
  nand2 gate1004(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1005(.a(s_65), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1006(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1007(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1008(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1443(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1444(.a(gate422inter0), .b(s_128), .O(gate422inter1));
  and2  gate1445(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1446(.a(s_128), .O(gate422inter3));
  inv1  gate1447(.a(s_129), .O(gate422inter4));
  nand2 gate1448(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1449(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1450(.a(G1039), .O(gate422inter7));
  inv1  gate1451(.a(G1135), .O(gate422inter8));
  nand2 gate1452(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1453(.a(s_129), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1454(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1455(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1456(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1639(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1640(.a(gate429inter0), .b(s_156), .O(gate429inter1));
  and2  gate1641(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1642(.a(s_156), .O(gate429inter3));
  inv1  gate1643(.a(s_157), .O(gate429inter4));
  nand2 gate1644(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1645(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1646(.a(G6), .O(gate429inter7));
  inv1  gate1647(.a(G1147), .O(gate429inter8));
  nand2 gate1648(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1649(.a(s_157), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1650(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1651(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1652(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate981(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate982(.a(gate431inter0), .b(s_62), .O(gate431inter1));
  and2  gate983(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate984(.a(s_62), .O(gate431inter3));
  inv1  gate985(.a(s_63), .O(gate431inter4));
  nand2 gate986(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate987(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate988(.a(G7), .O(gate431inter7));
  inv1  gate989(.a(G1150), .O(gate431inter8));
  nand2 gate990(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate991(.a(s_63), .b(gate431inter3), .O(gate431inter10));
  nor2  gate992(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate993(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate994(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1177(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1178(.a(gate434inter0), .b(s_90), .O(gate434inter1));
  and2  gate1179(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1180(.a(s_90), .O(gate434inter3));
  inv1  gate1181(.a(s_91), .O(gate434inter4));
  nand2 gate1182(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1183(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1184(.a(G1057), .O(gate434inter7));
  inv1  gate1185(.a(G1153), .O(gate434inter8));
  nand2 gate1186(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1187(.a(s_91), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1188(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1189(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1190(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1751(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1752(.a(gate443inter0), .b(s_172), .O(gate443inter1));
  and2  gate1753(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1754(.a(s_172), .O(gate443inter3));
  inv1  gate1755(.a(s_173), .O(gate443inter4));
  nand2 gate1756(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1757(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1758(.a(G13), .O(gate443inter7));
  inv1  gate1759(.a(G1168), .O(gate443inter8));
  nand2 gate1760(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1761(.a(s_173), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1762(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1763(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1764(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1345(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1346(.a(gate444inter0), .b(s_114), .O(gate444inter1));
  and2  gate1347(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1348(.a(s_114), .O(gate444inter3));
  inv1  gate1349(.a(s_115), .O(gate444inter4));
  nand2 gate1350(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1351(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1352(.a(G1072), .O(gate444inter7));
  inv1  gate1353(.a(G1168), .O(gate444inter8));
  nand2 gate1354(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1355(.a(s_115), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1356(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1357(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1358(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate757(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate758(.a(gate457inter0), .b(s_30), .O(gate457inter1));
  and2  gate759(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate760(.a(s_30), .O(gate457inter3));
  inv1  gate761(.a(s_31), .O(gate457inter4));
  nand2 gate762(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate763(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate764(.a(G20), .O(gate457inter7));
  inv1  gate765(.a(G1189), .O(gate457inter8));
  nand2 gate766(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate767(.a(s_31), .b(gate457inter3), .O(gate457inter10));
  nor2  gate768(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate769(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate770(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate603(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate604(.a(gate458inter0), .b(s_8), .O(gate458inter1));
  and2  gate605(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate606(.a(s_8), .O(gate458inter3));
  inv1  gate607(.a(s_9), .O(gate458inter4));
  nand2 gate608(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate609(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate610(.a(G1093), .O(gate458inter7));
  inv1  gate611(.a(G1189), .O(gate458inter8));
  nand2 gate612(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate613(.a(s_9), .b(gate458inter3), .O(gate458inter10));
  nor2  gate614(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate615(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate616(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1135(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1136(.a(gate459inter0), .b(s_84), .O(gate459inter1));
  and2  gate1137(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1138(.a(s_84), .O(gate459inter3));
  inv1  gate1139(.a(s_85), .O(gate459inter4));
  nand2 gate1140(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1141(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1142(.a(G21), .O(gate459inter7));
  inv1  gate1143(.a(G1192), .O(gate459inter8));
  nand2 gate1144(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1145(.a(s_85), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1146(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1147(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1148(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1625(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1626(.a(gate461inter0), .b(s_154), .O(gate461inter1));
  and2  gate1627(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1628(.a(s_154), .O(gate461inter3));
  inv1  gate1629(.a(s_155), .O(gate461inter4));
  nand2 gate1630(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1631(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1632(.a(G22), .O(gate461inter7));
  inv1  gate1633(.a(G1195), .O(gate461inter8));
  nand2 gate1634(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1635(.a(s_155), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1636(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1637(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1638(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1065(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1066(.a(gate465inter0), .b(s_74), .O(gate465inter1));
  and2  gate1067(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1068(.a(s_74), .O(gate465inter3));
  inv1  gate1069(.a(s_75), .O(gate465inter4));
  nand2 gate1070(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1071(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1072(.a(G24), .O(gate465inter7));
  inv1  gate1073(.a(G1201), .O(gate465inter8));
  nand2 gate1074(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1075(.a(s_75), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1076(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1077(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1078(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1919(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1920(.a(gate471inter0), .b(s_196), .O(gate471inter1));
  and2  gate1921(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1922(.a(s_196), .O(gate471inter3));
  inv1  gate1923(.a(s_197), .O(gate471inter4));
  nand2 gate1924(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1925(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1926(.a(G27), .O(gate471inter7));
  inv1  gate1927(.a(G1210), .O(gate471inter8));
  nand2 gate1928(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1929(.a(s_197), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1930(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1931(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1932(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1037(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1038(.a(gate476inter0), .b(s_70), .O(gate476inter1));
  and2  gate1039(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1040(.a(s_70), .O(gate476inter3));
  inv1  gate1041(.a(s_71), .O(gate476inter4));
  nand2 gate1042(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1043(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1044(.a(G1120), .O(gate476inter7));
  inv1  gate1045(.a(G1216), .O(gate476inter8));
  nand2 gate1046(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1047(.a(s_71), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1048(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1049(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1050(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1219(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1220(.a(gate481inter0), .b(s_96), .O(gate481inter1));
  and2  gate1221(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1222(.a(s_96), .O(gate481inter3));
  inv1  gate1223(.a(s_97), .O(gate481inter4));
  nand2 gate1224(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1225(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1226(.a(G32), .O(gate481inter7));
  inv1  gate1227(.a(G1225), .O(gate481inter8));
  nand2 gate1228(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1229(.a(s_97), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1230(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1231(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1232(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate1555(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1556(.a(gate482inter0), .b(s_144), .O(gate482inter1));
  and2  gate1557(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1558(.a(s_144), .O(gate482inter3));
  inv1  gate1559(.a(s_145), .O(gate482inter4));
  nand2 gate1560(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1561(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1562(.a(G1129), .O(gate482inter7));
  inv1  gate1563(.a(G1225), .O(gate482inter8));
  nand2 gate1564(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1565(.a(s_145), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1566(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1567(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1568(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate575(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate576(.a(gate483inter0), .b(s_4), .O(gate483inter1));
  and2  gate577(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate578(.a(s_4), .O(gate483inter3));
  inv1  gate579(.a(s_5), .O(gate483inter4));
  nand2 gate580(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate581(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate582(.a(G1228), .O(gate483inter7));
  inv1  gate583(.a(G1229), .O(gate483inter8));
  nand2 gate584(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate585(.a(s_5), .b(gate483inter3), .O(gate483inter10));
  nor2  gate586(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate587(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate588(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1401(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1402(.a(gate486inter0), .b(s_122), .O(gate486inter1));
  and2  gate1403(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1404(.a(s_122), .O(gate486inter3));
  inv1  gate1405(.a(s_123), .O(gate486inter4));
  nand2 gate1406(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1407(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1408(.a(G1234), .O(gate486inter7));
  inv1  gate1409(.a(G1235), .O(gate486inter8));
  nand2 gate1410(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1411(.a(s_123), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1412(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1413(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1414(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate785(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate786(.a(gate495inter0), .b(s_34), .O(gate495inter1));
  and2  gate787(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate788(.a(s_34), .O(gate495inter3));
  inv1  gate789(.a(s_35), .O(gate495inter4));
  nand2 gate790(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate791(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate792(.a(G1252), .O(gate495inter7));
  inv1  gate793(.a(G1253), .O(gate495inter8));
  nand2 gate794(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate795(.a(s_35), .b(gate495inter3), .O(gate495inter10));
  nor2  gate796(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate797(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate798(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate953(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate954(.a(gate500inter0), .b(s_58), .O(gate500inter1));
  and2  gate955(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate956(.a(s_58), .O(gate500inter3));
  inv1  gate957(.a(s_59), .O(gate500inter4));
  nand2 gate958(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate959(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate960(.a(G1262), .O(gate500inter7));
  inv1  gate961(.a(G1263), .O(gate500inter8));
  nand2 gate962(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate963(.a(s_59), .b(gate500inter3), .O(gate500inter10));
  nor2  gate964(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate965(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate966(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1331(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1332(.a(gate501inter0), .b(s_112), .O(gate501inter1));
  and2  gate1333(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1334(.a(s_112), .O(gate501inter3));
  inv1  gate1335(.a(s_113), .O(gate501inter4));
  nand2 gate1336(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1337(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1338(.a(G1264), .O(gate501inter7));
  inv1  gate1339(.a(G1265), .O(gate501inter8));
  nand2 gate1340(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1341(.a(s_113), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1342(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1343(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1344(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate771(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate772(.a(gate503inter0), .b(s_32), .O(gate503inter1));
  and2  gate773(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate774(.a(s_32), .O(gate503inter3));
  inv1  gate775(.a(s_33), .O(gate503inter4));
  nand2 gate776(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate777(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate778(.a(G1268), .O(gate503inter7));
  inv1  gate779(.a(G1269), .O(gate503inter8));
  nand2 gate780(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate781(.a(s_33), .b(gate503inter3), .O(gate503inter10));
  nor2  gate782(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate783(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate784(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate855(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate856(.a(gate507inter0), .b(s_44), .O(gate507inter1));
  and2  gate857(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate858(.a(s_44), .O(gate507inter3));
  inv1  gate859(.a(s_45), .O(gate507inter4));
  nand2 gate860(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate861(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate862(.a(G1276), .O(gate507inter7));
  inv1  gate863(.a(G1277), .O(gate507inter8));
  nand2 gate864(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate865(.a(s_45), .b(gate507inter3), .O(gate507inter10));
  nor2  gate866(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate867(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate868(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate729(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate730(.a(gate512inter0), .b(s_26), .O(gate512inter1));
  and2  gate731(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate732(.a(s_26), .O(gate512inter3));
  inv1  gate733(.a(s_27), .O(gate512inter4));
  nand2 gate734(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate735(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate736(.a(G1286), .O(gate512inter7));
  inv1  gate737(.a(G1287), .O(gate512inter8));
  nand2 gate738(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate739(.a(s_27), .b(gate512inter3), .O(gate512inter10));
  nor2  gate740(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate741(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate742(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule