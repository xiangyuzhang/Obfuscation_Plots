module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );

  xor2  gate245(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate246(.a(gate25inter0), .b(s_12), .O(gate25inter1));
  and2  gate247(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate248(.a(s_12), .O(gate25inter3));
  inv1  gate249(.a(s_13), .O(gate25inter4));
  nand2 gate250(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate251(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate252(.a(N134), .O(gate25inter7));
  inv1  gate253(.a(N56), .O(gate25inter8));
  nand2 gate254(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate255(.a(s_13), .b(gate25inter3), .O(gate25inter10));
  nor2  gate256(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate257(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate258(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate217(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate218(.a(gate28inter0), .b(s_8), .O(gate28inter1));
  and2  gate219(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate220(.a(s_8), .O(gate28inter3));
  inv1  gate221(.a(s_9), .O(gate28inter4));
  nand2 gate222(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate223(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate224(.a(N146), .O(gate28inter7));
  inv1  gate225(.a(N95), .O(gate28inter8));
  nand2 gate226(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate227(.a(s_9), .b(gate28inter3), .O(gate28inter10));
  nor2  gate228(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate229(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate230(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate189(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate190(.a(gate32inter0), .b(s_4), .O(gate32inter1));
  and2  gate191(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate192(.a(s_4), .O(gate32inter3));
  inv1  gate193(.a(s_5), .O(gate32inter4));
  nand2 gate194(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate195(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate196(.a(N34), .O(gate32inter7));
  inv1  gate197(.a(N127), .O(gate32inter8));
  nand2 gate198(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate199(.a(s_5), .b(gate32inter3), .O(gate32inter10));
  nor2  gate200(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate201(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate202(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );

  xor2  gate273(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate274(.a(gate35inter0), .b(s_16), .O(gate35inter1));
  and2  gate275(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate276(.a(s_16), .O(gate35inter3));
  inv1  gate277(.a(s_17), .O(gate35inter4));
  nand2 gate278(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate279(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate280(.a(N53), .O(gate35inter7));
  inv1  gate281(.a(N131), .O(gate35inter8));
  nand2 gate282(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate283(.a(s_17), .b(gate35inter3), .O(gate35inter10));
  nor2  gate284(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate285(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate286(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );

  xor2  gate175(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate176(.a(gate44inter0), .b(s_2), .O(gate44inter1));
  and2  gate177(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate178(.a(s_2), .O(gate44inter3));
  inv1  gate179(.a(s_3), .O(gate44inter4));
  nand2 gate180(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate181(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate182(.a(N112), .O(gate44inter7));
  inv1  gate183(.a(N151), .O(gate44inter8));
  nand2 gate184(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate185(.a(s_3), .b(gate44inter3), .O(gate44inter10));
  nor2  gate186(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate187(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate188(.a(gate44inter12), .b(gate44inter1), .O(N197));
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate315(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate316(.a(gate50inter0), .b(s_22), .O(gate50inter1));
  and2  gate317(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate318(.a(s_22), .O(gate50inter3));
  inv1  gate319(.a(s_23), .O(gate50inter4));
  nand2 gate320(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate321(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate322(.a(N203), .O(gate50inter7));
  inv1  gate323(.a(N154), .O(gate50inter8));
  nand2 gate324(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate325(.a(s_23), .b(gate50inter3), .O(gate50inter10));
  nor2  gate326(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate327(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate328(.a(gate50inter12), .b(gate50inter1), .O(N224));
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );

  xor2  gate343(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate344(.a(gate54inter0), .b(s_26), .O(gate54inter1));
  and2  gate345(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate346(.a(s_26), .O(gate54inter3));
  inv1  gate347(.a(s_27), .O(gate54inter4));
  nand2 gate348(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate349(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate350(.a(N203), .O(gate54inter7));
  inv1  gate351(.a(N168), .O(gate54inter8));
  nand2 gate352(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate353(.a(s_27), .b(gate54inter3), .O(gate54inter10));
  nor2  gate354(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate355(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate356(.a(gate54inter12), .b(gate54inter1), .O(N236));
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate371(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate372(.a(gate70inter0), .b(s_30), .O(gate70inter1));
  and2  gate373(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate374(.a(s_30), .O(gate70inter3));
  inv1  gate375(.a(s_31), .O(gate70inter4));
  nand2 gate376(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate377(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate378(.a(N227), .O(gate70inter7));
  inv1  gate379(.a(N183), .O(gate70inter8));
  nand2 gate380(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate381(.a(s_31), .b(gate70inter3), .O(gate70inter10));
  nor2  gate382(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate383(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate384(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate259(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate260(.a(gate75inter0), .b(s_14), .O(gate75inter1));
  and2  gate261(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate262(.a(s_14), .O(gate75inter3));
  inv1  gate263(.a(s_15), .O(gate75inter4));
  nand2 gate264(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate265(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate266(.a(N243), .O(gate75inter7));
  inv1  gate267(.a(N193), .O(gate75inter8));
  nand2 gate268(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate269(.a(s_15), .b(gate75inter3), .O(gate75inter10));
  nor2  gate270(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate271(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate272(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );

  xor2  gate329(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate330(.a(gate79inter0), .b(s_24), .O(gate79inter1));
  and2  gate331(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate332(.a(s_24), .O(gate79inter3));
  inv1  gate333(.a(s_25), .O(gate79inter4));
  nand2 gate334(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate335(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate336(.a(N230), .O(gate79inter7));
  inv1  gate337(.a(N186), .O(gate79inter8));
  nand2 gate338(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate339(.a(s_25), .b(gate79inter3), .O(gate79inter10));
  nor2  gate340(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate341(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate342(.a(gate79inter12), .b(gate79inter1), .O(N289));
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate161(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate162(.a(gate111inter0), .b(s_0), .O(gate111inter1));
  and2  gate163(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate164(.a(s_0), .O(gate111inter3));
  inv1  gate165(.a(s_1), .O(gate111inter4));
  nand2 gate166(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate167(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate168(.a(N319), .O(gate111inter7));
  inv1  gate169(.a(N60), .O(gate111inter8));
  nand2 gate170(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate171(.a(s_1), .b(gate111inter3), .O(gate111inter10));
  nor2  gate172(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate173(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate174(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate357(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate358(.a(gate115inter0), .b(s_28), .O(gate115inter1));
  and2  gate359(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate360(.a(s_28), .O(gate115inter3));
  inv1  gate361(.a(s_29), .O(gate115inter4));
  nand2 gate362(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate363(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate364(.a(N319), .O(gate115inter7));
  inv1  gate365(.a(N99), .O(gate115inter8));
  nand2 gate366(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate367(.a(s_29), .b(gate115inter3), .O(gate115inter10));
  nor2  gate368(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate369(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate370(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );

  xor2  gate203(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate204(.a(gate122inter0), .b(s_6), .O(gate122inter1));
  and2  gate205(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate206(.a(s_6), .O(gate122inter3));
  inv1  gate207(.a(s_7), .O(gate122inter4));
  nand2 gate208(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate209(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate210(.a(N337), .O(gate122inter7));
  inv1  gate211(.a(N305), .O(gate122inter8));
  nand2 gate212(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate213(.a(s_7), .b(gate122inter3), .O(gate122inter10));
  nor2  gate214(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate215(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate216(.a(gate122inter12), .b(gate122inter1), .O(N353));

  xor2  gate301(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate302(.a(gate123inter0), .b(s_20), .O(gate123inter1));
  and2  gate303(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate304(.a(s_20), .O(gate123inter3));
  inv1  gate305(.a(s_21), .O(gate123inter4));
  nand2 gate306(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate307(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate308(.a(N339), .O(gate123inter7));
  inv1  gate309(.a(N306), .O(gate123inter8));
  nand2 gate310(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate311(.a(s_21), .b(gate123inter3), .O(gate123inter10));
  nor2  gate312(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate313(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate314(.a(gate123inter12), .b(gate123inter1), .O(N354));
nand2 gate124( .a(N341), .b(N307), .O(N355) );

  xor2  gate231(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate232(.a(gate125inter0), .b(s_10), .O(gate125inter1));
  and2  gate233(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate234(.a(s_10), .O(gate125inter3));
  inv1  gate235(.a(s_11), .O(gate125inter4));
  nand2 gate236(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate237(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate238(.a(N343), .O(gate125inter7));
  inv1  gate239(.a(N308), .O(gate125inter8));
  nand2 gate240(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate241(.a(s_11), .b(gate125inter3), .O(gate125inter10));
  nor2  gate242(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate243(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate244(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );

  xor2  gate287(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate288(.a(gate154inter0), .b(s_18), .O(gate154inter1));
  and2  gate289(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate290(.a(s_18), .O(gate154inter3));
  inv1  gate291(.a(s_19), .O(gate154inter4));
  nand2 gate292(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate293(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate294(.a(N386), .O(gate154inter7));
  inv1  gate295(.a(N417), .O(gate154inter8));
  nand2 gate296(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate297(.a(s_19), .b(gate154inter3), .O(gate154inter10));
  nor2  gate298(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate299(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate300(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule