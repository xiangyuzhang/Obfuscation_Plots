module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12;

  xor2  gate231(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate232(.a(gate1inter0), .b(s_4), .O(gate1inter1));
  and2  gate233(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate234(.a(s_4), .O(gate1inter3));
  inv1  gate235(.a(s_5), .O(gate1inter4));
  nand2 gate236(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate237(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate238(.a(N1), .O(gate1inter7));
  inv1  gate239(.a(N5), .O(gate1inter8));
  nand2 gate240(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate241(.a(s_5), .b(gate1inter3), .O(gate1inter10));
  nor2  gate242(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate243(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate244(.a(gate1inter12), .b(gate1inter1), .O(N250));
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );

  xor2  gate203(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate204(.a(gate5inter0), .b(s_0), .O(gate5inter1));
  and2  gate205(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate206(.a(s_0), .O(gate5inter3));
  inv1  gate207(.a(s_1), .O(gate5inter4));
  nand2 gate208(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate209(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate210(.a(N33), .O(gate5inter7));
  inv1  gate211(.a(N37), .O(gate5inter8));
  nand2 gate212(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate213(.a(s_1), .b(gate5inter3), .O(gate5inter10));
  nor2  gate214(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate215(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate216(.a(gate5inter12), .b(gate5inter1), .O(N254));
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate273(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate274(.a(gate8inter0), .b(s_10), .O(gate8inter1));
  and2  gate275(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate276(.a(s_10), .O(gate8inter3));
  inv1  gate277(.a(s_11), .O(gate8inter4));
  nand2 gate278(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate279(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate280(.a(N57), .O(gate8inter7));
  inv1  gate281(.a(N61), .O(gate8inter8));
  nand2 gate282(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate283(.a(s_11), .b(gate8inter3), .O(gate8inter10));
  nor2  gate284(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate285(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate286(.a(gate8inter12), .b(gate8inter1), .O(N257));
xor2 gate9( .a(N65), .b(N69), .O(N258) );

  xor2  gate371(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate372(.a(gate10inter0), .b(s_24), .O(gate10inter1));
  and2  gate373(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate374(.a(s_24), .O(gate10inter3));
  inv1  gate375(.a(s_25), .O(gate10inter4));
  nand2 gate376(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate377(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate378(.a(N73), .O(gate10inter7));
  inv1  gate379(.a(N77), .O(gate10inter8));
  nand2 gate380(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate381(.a(s_25), .b(gate10inter3), .O(gate10inter10));
  nor2  gate382(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate383(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate384(.a(gate10inter12), .b(gate10inter1), .O(N259));
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );

  xor2  gate329(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate330(.a(gate28inter0), .b(s_18), .O(gate28inter1));
  and2  gate331(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate332(.a(s_18), .O(gate28inter3));
  inv1  gate333(.a(s_19), .O(gate28inter4));
  nand2 gate334(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate335(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate336(.a(N37), .O(gate28inter7));
  inv1  gate337(.a(N53), .O(gate28inter8));
  nand2 gate338(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate339(.a(s_19), .b(gate28inter3), .O(gate28inter10));
  nor2  gate340(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate341(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate342(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate553(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate554(.a(gate30inter0), .b(s_50), .O(gate30inter1));
  and2  gate555(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate556(.a(s_50), .O(gate30inter3));
  inv1  gate557(.a(s_51), .O(gate30inter4));
  nand2 gate558(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate559(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate560(.a(N41), .O(gate30inter7));
  inv1  gate561(.a(N57), .O(gate30inter8));
  nand2 gate562(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate563(.a(s_51), .b(gate30inter3), .O(gate30inter10));
  nor2  gate564(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate565(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate566(.a(gate30inter12), .b(gate30inter1), .O(N279));

  xor2  gate483(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate484(.a(gate31inter0), .b(s_40), .O(gate31inter1));
  and2  gate485(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate486(.a(s_40), .O(gate31inter3));
  inv1  gate487(.a(s_41), .O(gate31inter4));
  nand2 gate488(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate489(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate490(.a(N13), .O(gate31inter7));
  inv1  gate491(.a(N29), .O(gate31inter8));
  nand2 gate492(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate493(.a(s_41), .b(gate31inter3), .O(gate31inter10));
  nor2  gate494(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate495(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate496(.a(gate31inter12), .b(gate31inter1), .O(N280));
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );

  xor2  gate315(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate316(.a(gate36inter0), .b(s_16), .O(gate36inter1));
  and2  gate317(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate318(.a(s_16), .O(gate36inter3));
  inv1  gate319(.a(s_17), .O(gate36inter4));
  nand2 gate320(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate321(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate322(.a(N101), .O(gate36inter7));
  inv1  gate323(.a(N117), .O(gate36inter8));
  nand2 gate324(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate325(.a(s_17), .b(gate36inter3), .O(gate36inter10));
  nor2  gate326(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate327(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate328(.a(gate36inter12), .b(gate36inter1), .O(N285));
xor2 gate37( .a(N73), .b(N89), .O(N286) );

  xor2  gate567(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate568(.a(gate38inter0), .b(s_52), .O(gate38inter1));
  and2  gate569(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate570(.a(s_52), .O(gate38inter3));
  inv1  gate571(.a(s_53), .O(gate38inter4));
  nand2 gate572(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate573(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate574(.a(N105), .O(gate38inter7));
  inv1  gate575(.a(N121), .O(gate38inter8));
  nand2 gate576(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate577(.a(s_53), .b(gate38inter3), .O(gate38inter10));
  nor2  gate578(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate579(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate580(.a(gate38inter12), .b(gate38inter1), .O(N287));
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );

  xor2  gate259(.a(N257), .b(N256), .O(gate44inter0));
  nand2 gate260(.a(gate44inter0), .b(s_8), .O(gate44inter1));
  and2  gate261(.a(N257), .b(N256), .O(gate44inter2));
  inv1  gate262(.a(s_8), .O(gate44inter3));
  inv1  gate263(.a(s_9), .O(gate44inter4));
  nand2 gate264(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate265(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate266(.a(N256), .O(gate44inter7));
  inv1  gate267(.a(N257), .O(gate44inter8));
  nand2 gate268(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate269(.a(s_9), .b(gate44inter3), .O(gate44inter10));
  nor2  gate270(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate271(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate272(.a(gate44inter12), .b(gate44inter1), .O(N299));

  xor2  gate595(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate596(.a(gate45inter0), .b(s_56), .O(gate45inter1));
  and2  gate597(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate598(.a(s_56), .O(gate45inter3));
  inv1  gate599(.a(s_57), .O(gate45inter4));
  nand2 gate600(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate601(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate602(.a(N258), .O(gate45inter7));
  inv1  gate603(.a(N259), .O(gate45inter8));
  nand2 gate604(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate605(.a(s_57), .b(gate45inter3), .O(gate45inter10));
  nor2  gate606(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate607(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate608(.a(gate45inter12), .b(gate45inter1), .O(N302));

  xor2  gate511(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate512(.a(gate46inter0), .b(s_44), .O(gate46inter1));
  and2  gate513(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate514(.a(s_44), .O(gate46inter3));
  inv1  gate515(.a(s_45), .O(gate46inter4));
  nand2 gate516(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate517(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate518(.a(N260), .O(gate46inter7));
  inv1  gate519(.a(N261), .O(gate46inter8));
  nand2 gate520(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate521(.a(s_45), .b(gate46inter3), .O(gate46inter10));
  nor2  gate522(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate523(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate524(.a(gate46inter12), .b(gate46inter1), .O(N305));

  xor2  gate343(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate344(.a(gate47inter0), .b(s_20), .O(gate47inter1));
  and2  gate345(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate346(.a(s_20), .O(gate47inter3));
  inv1  gate347(.a(s_21), .O(gate47inter4));
  nand2 gate348(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate349(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate350(.a(N262), .O(gate47inter7));
  inv1  gate351(.a(N263), .O(gate47inter8));
  nand2 gate352(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate353(.a(s_21), .b(gate47inter3), .O(gate47inter10));
  nor2  gate354(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate355(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate356(.a(gate47inter12), .b(gate47inter1), .O(N308));

  xor2  gate399(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate400(.a(gate48inter0), .b(s_28), .O(gate48inter1));
  and2  gate401(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate402(.a(s_28), .O(gate48inter3));
  inv1  gate403(.a(s_29), .O(gate48inter4));
  nand2 gate404(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate405(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate406(.a(N264), .O(gate48inter7));
  inv1  gate407(.a(N265), .O(gate48inter8));
  nand2 gate408(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate409(.a(s_29), .b(gate48inter3), .O(gate48inter10));
  nor2  gate410(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate411(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate412(.a(gate48inter12), .b(gate48inter1), .O(N311));
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate609(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate610(.a(gate50inter0), .b(s_58), .O(gate50inter1));
  and2  gate611(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate612(.a(s_58), .O(gate50inter3));
  inv1  gate613(.a(s_59), .O(gate50inter4));
  nand2 gate614(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate615(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate616(.a(N276), .O(gate50inter7));
  inv1  gate617(.a(N277), .O(gate50inter8));
  nand2 gate618(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate619(.a(s_59), .b(gate50inter3), .O(gate50inter10));
  nor2  gate620(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate621(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate622(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );

  xor2  gate413(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate414(.a(gate66inter0), .b(s_30), .O(gate66inter1));
  and2  gate415(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate416(.a(s_30), .O(gate66inter3));
  inv1  gate417(.a(s_31), .O(gate66inter4));
  nand2 gate418(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate419(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate420(.a(N267), .O(gate66inter7));
  inv1  gate421(.a(N343), .O(gate66inter8));
  nand2 gate422(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate423(.a(s_31), .b(gate66inter3), .O(gate66inter10));
  nor2  gate424(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate425(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate426(.a(gate66inter12), .b(gate66inter1), .O(N347));
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate539(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate540(.a(gate70inter0), .b(s_48), .O(gate70inter1));
  and2  gate541(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate542(.a(s_48), .O(gate70inter3));
  inv1  gate543(.a(s_49), .O(gate70inter4));
  nand2 gate544(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate545(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate546(.a(N271), .O(gate70inter7));
  inv1  gate547(.a(N339), .O(gate70inter8));
  nand2 gate548(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate549(.a(s_49), .b(gate70inter3), .O(gate70inter10));
  nor2  gate550(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate551(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate552(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );

  xor2  gate581(.a(N341), .b(N273), .O(gate72inter0));
  nand2 gate582(.a(gate72inter0), .b(s_54), .O(gate72inter1));
  and2  gate583(.a(N341), .b(N273), .O(gate72inter2));
  inv1  gate584(.a(s_54), .O(gate72inter3));
  inv1  gate585(.a(s_55), .O(gate72inter4));
  nand2 gate586(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate587(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate588(.a(N273), .O(gate72inter7));
  inv1  gate589(.a(N341), .O(gate72inter8));
  nand2 gate590(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate591(.a(s_55), .b(gate72inter3), .O(gate72inter10));
  nor2  gate592(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate593(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate594(.a(gate72inter12), .b(gate72inter1), .O(N353));

  xor2  gate525(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate526(.a(gate73inter0), .b(s_46), .O(gate73inter1));
  and2  gate527(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate528(.a(s_46), .O(gate73inter3));
  inv1  gate529(.a(s_47), .O(gate73inter4));
  nand2 gate530(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate531(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate532(.a(N314), .O(gate73inter7));
  inv1  gate533(.a(N346), .O(gate73inter8));
  nand2 gate534(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate535(.a(s_47), .b(gate73inter3), .O(gate73inter10));
  nor2  gate536(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate537(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate538(.a(gate73inter12), .b(gate73inter1), .O(N354));
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );

  xor2  gate301(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate302(.a(gate78inter0), .b(s_14), .O(gate78inter1));
  and2  gate303(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate304(.a(s_14), .O(gate78inter3));
  inv1  gate305(.a(s_15), .O(gate78inter4));
  nand2 gate306(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate307(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate308(.a(N319), .O(gate78inter7));
  inv1  gate309(.a(N351), .O(gate78inter8));
  nand2 gate310(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate311(.a(s_15), .b(gate78inter3), .O(gate78inter10));
  nor2  gate312(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate313(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate314(.a(gate78inter12), .b(gate78inter1), .O(N419));
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate427(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate428(.a(gate80inter0), .b(s_32), .O(gate80inter1));
  and2  gate429(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate430(.a(s_32), .O(gate80inter3));
  inv1  gate431(.a(s_33), .O(gate80inter4));
  nand2 gate432(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate433(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate434(.a(N321), .O(gate80inter7));
  inv1  gate435(.a(N353), .O(gate80inter8));
  nand2 gate436(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate437(.a(s_33), .b(gate80inter3), .O(gate80inter10));
  nor2  gate438(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate439(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate440(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate287(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate288(.a(gate172inter0), .b(s_12), .O(gate172inter1));
  and2  gate289(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate290(.a(s_12), .O(gate172inter3));
  inv1  gate291(.a(s_13), .O(gate172inter4));
  nand2 gate292(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate293(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate294(.a(N5), .O(gate172inter7));
  inv1  gate295(.a(N693), .O(gate172inter8));
  nand2 gate296(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate297(.a(s_13), .b(gate172inter3), .O(gate172inter10));
  nor2  gate298(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate299(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate300(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate497(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate498(.a(gate177inter0), .b(s_42), .O(gate177inter1));
  and2  gate499(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate500(.a(s_42), .O(gate177inter3));
  inv1  gate501(.a(s_43), .O(gate177inter4));
  nand2 gate502(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate503(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate504(.a(N25), .O(gate177inter7));
  inv1  gate505(.a(N698), .O(gate177inter8));
  nand2 gate506(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate507(.a(s_43), .b(gate177inter3), .O(gate177inter10));
  nor2  gate508(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate509(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate510(.a(gate177inter12), .b(gate177inter1), .O(N730));

  xor2  gate357(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate358(.a(gate178inter0), .b(s_22), .O(gate178inter1));
  and2  gate359(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate360(.a(s_22), .O(gate178inter3));
  inv1  gate361(.a(s_23), .O(gate178inter4));
  nand2 gate362(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate363(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate364(.a(N29), .O(gate178inter7));
  inv1  gate365(.a(N699), .O(gate178inter8));
  nand2 gate366(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate367(.a(s_23), .b(gate178inter3), .O(gate178inter10));
  nor2  gate368(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate369(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate370(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );

  xor2  gate623(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate624(.a(gate182inter0), .b(s_60), .O(gate182inter1));
  and2  gate625(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate626(.a(s_60), .O(gate182inter3));
  inv1  gate627(.a(s_61), .O(gate182inter4));
  nand2 gate628(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate629(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate630(.a(N45), .O(gate182inter7));
  inv1  gate631(.a(N703), .O(gate182inter8));
  nand2 gate632(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate633(.a(s_61), .b(gate182inter3), .O(gate182inter10));
  nor2  gate634(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate635(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate636(.a(gate182inter12), .b(gate182inter1), .O(N735));
xor2 gate183( .a(N49), .b(N704), .O(N736) );

  xor2  gate455(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate456(.a(gate184inter0), .b(s_36), .O(gate184inter1));
  and2  gate457(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate458(.a(s_36), .O(gate184inter3));
  inv1  gate459(.a(s_37), .O(gate184inter4));
  nand2 gate460(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate461(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate462(.a(N53), .O(gate184inter7));
  inv1  gate463(.a(N705), .O(gate184inter8));
  nand2 gate464(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate465(.a(s_37), .b(gate184inter3), .O(gate184inter10));
  nor2  gate466(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate467(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate468(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );

  xor2  gate385(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate386(.a(gate191inter0), .b(s_26), .O(gate191inter1));
  and2  gate387(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate388(.a(s_26), .O(gate191inter3));
  inv1  gate389(.a(s_27), .O(gate191inter4));
  nand2 gate390(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate391(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate392(.a(N81), .O(gate191inter7));
  inv1  gate393(.a(N712), .O(gate191inter8));
  nand2 gate394(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate395(.a(s_27), .b(gate191inter3), .O(gate191inter10));
  nor2  gate396(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate397(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate398(.a(gate191inter12), .b(gate191inter1), .O(N744));
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );

  xor2  gate469(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate470(.a(gate196inter0), .b(s_38), .O(gate196inter1));
  and2  gate471(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate472(.a(s_38), .O(gate196inter3));
  inv1  gate473(.a(s_39), .O(gate196inter4));
  nand2 gate474(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate475(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate476(.a(N101), .O(gate196inter7));
  inv1  gate477(.a(N717), .O(gate196inter8));
  nand2 gate478(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate479(.a(s_39), .b(gate196inter3), .O(gate196inter10));
  nor2  gate480(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate481(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate482(.a(gate196inter12), .b(gate196inter1), .O(N749));
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );

  xor2  gate245(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate246(.a(gate199inter0), .b(s_6), .O(gate199inter1));
  and2  gate247(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate248(.a(s_6), .O(gate199inter3));
  inv1  gate249(.a(s_7), .O(gate199inter4));
  nand2 gate250(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate251(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate252(.a(N113), .O(gate199inter7));
  inv1  gate253(.a(N720), .O(gate199inter8));
  nand2 gate254(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate255(.a(s_7), .b(gate199inter3), .O(gate199inter10));
  nor2  gate256(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate257(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate258(.a(gate199inter12), .b(gate199inter1), .O(N752));

  xor2  gate217(.a(N721), .b(N117), .O(gate200inter0));
  nand2 gate218(.a(gate200inter0), .b(s_2), .O(gate200inter1));
  and2  gate219(.a(N721), .b(N117), .O(gate200inter2));
  inv1  gate220(.a(s_2), .O(gate200inter3));
  inv1  gate221(.a(s_3), .O(gate200inter4));
  nand2 gate222(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate223(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate224(.a(N117), .O(gate200inter7));
  inv1  gate225(.a(N721), .O(gate200inter8));
  nand2 gate226(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate227(.a(s_3), .b(gate200inter3), .O(gate200inter10));
  nor2  gate228(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate229(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate230(.a(gate200inter12), .b(gate200inter1), .O(N753));

  xor2  gate441(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate442(.a(gate201inter0), .b(s_34), .O(gate201inter1));
  and2  gate443(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate444(.a(s_34), .O(gate201inter3));
  inv1  gate445(.a(s_35), .O(gate201inter4));
  nand2 gate446(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate447(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate448(.a(N121), .O(gate201inter7));
  inv1  gate449(.a(N722), .O(gate201inter8));
  nand2 gate450(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate451(.a(s_35), .b(gate201inter3), .O(gate201inter10));
  nor2  gate452(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate453(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate454(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule