module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381, s_382, s_383, s_384, s_385, s_386, s_387, s_388, s_389, s_390, s_391;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate3235(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate3236(.a(gate9inter0), .b(s_384), .O(gate9inter1));
  and2  gate3237(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate3238(.a(s_384), .O(gate9inter3));
  inv1  gate3239(.a(s_385), .O(gate9inter4));
  nand2 gate3240(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate3241(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate3242(.a(G1), .O(gate9inter7));
  inv1  gate3243(.a(G2), .O(gate9inter8));
  nand2 gate3244(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate3245(.a(s_385), .b(gate9inter3), .O(gate9inter10));
  nor2  gate3246(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate3247(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate3248(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1065(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1066(.a(gate10inter0), .b(s_74), .O(gate10inter1));
  and2  gate1067(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1068(.a(s_74), .O(gate10inter3));
  inv1  gate1069(.a(s_75), .O(gate10inter4));
  nand2 gate1070(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1071(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1072(.a(G3), .O(gate10inter7));
  inv1  gate1073(.a(G4), .O(gate10inter8));
  nand2 gate1074(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1075(.a(s_75), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1076(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1077(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1078(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2101(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2102(.a(gate12inter0), .b(s_222), .O(gate12inter1));
  and2  gate2103(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2104(.a(s_222), .O(gate12inter3));
  inv1  gate2105(.a(s_223), .O(gate12inter4));
  nand2 gate2106(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2107(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2108(.a(G7), .O(gate12inter7));
  inv1  gate2109(.a(G8), .O(gate12inter8));
  nand2 gate2110(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2111(.a(s_223), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2112(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2113(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2114(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1625(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1626(.a(gate16inter0), .b(s_154), .O(gate16inter1));
  and2  gate1627(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1628(.a(s_154), .O(gate16inter3));
  inv1  gate1629(.a(s_155), .O(gate16inter4));
  nand2 gate1630(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1631(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1632(.a(G15), .O(gate16inter7));
  inv1  gate1633(.a(G16), .O(gate16inter8));
  nand2 gate1634(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1635(.a(s_155), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1636(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1637(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1638(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate3249(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate3250(.a(gate17inter0), .b(s_386), .O(gate17inter1));
  and2  gate3251(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate3252(.a(s_386), .O(gate17inter3));
  inv1  gate3253(.a(s_387), .O(gate17inter4));
  nand2 gate3254(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate3255(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate3256(.a(G17), .O(gate17inter7));
  inv1  gate3257(.a(G18), .O(gate17inter8));
  nand2 gate3258(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate3259(.a(s_387), .b(gate17inter3), .O(gate17inter10));
  nor2  gate3260(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate3261(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate3262(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2283(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2284(.a(gate21inter0), .b(s_248), .O(gate21inter1));
  and2  gate2285(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2286(.a(s_248), .O(gate21inter3));
  inv1  gate2287(.a(s_249), .O(gate21inter4));
  nand2 gate2288(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2289(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2290(.a(G25), .O(gate21inter7));
  inv1  gate2291(.a(G26), .O(gate21inter8));
  nand2 gate2292(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2293(.a(s_249), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2294(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2295(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2296(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2003(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2004(.a(gate22inter0), .b(s_208), .O(gate22inter1));
  and2  gate2005(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2006(.a(s_208), .O(gate22inter3));
  inv1  gate2007(.a(s_209), .O(gate22inter4));
  nand2 gate2008(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2009(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2010(.a(G27), .O(gate22inter7));
  inv1  gate2011(.a(G28), .O(gate22inter8));
  nand2 gate2012(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2013(.a(s_209), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2014(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2015(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2016(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1541(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1542(.a(gate27inter0), .b(s_142), .O(gate27inter1));
  and2  gate1543(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1544(.a(s_142), .O(gate27inter3));
  inv1  gate1545(.a(s_143), .O(gate27inter4));
  nand2 gate1546(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1547(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1548(.a(G2), .O(gate27inter7));
  inv1  gate1549(.a(G6), .O(gate27inter8));
  nand2 gate1550(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1551(.a(s_143), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1552(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1553(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1554(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate2633(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2634(.a(gate28inter0), .b(s_298), .O(gate28inter1));
  and2  gate2635(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2636(.a(s_298), .O(gate28inter3));
  inv1  gate2637(.a(s_299), .O(gate28inter4));
  nand2 gate2638(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2639(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2640(.a(G10), .O(gate28inter7));
  inv1  gate2641(.a(G14), .O(gate28inter8));
  nand2 gate2642(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2643(.a(s_299), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2644(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2645(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2646(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate547(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate548(.a(gate30inter0), .b(s_0), .O(gate30inter1));
  and2  gate549(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate550(.a(s_0), .O(gate30inter3));
  inv1  gate551(.a(s_1), .O(gate30inter4));
  nand2 gate552(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate553(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate554(.a(G11), .O(gate30inter7));
  inv1  gate555(.a(G15), .O(gate30inter8));
  nand2 gate556(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate557(.a(s_1), .b(gate30inter3), .O(gate30inter10));
  nor2  gate558(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate559(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate560(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate883(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate884(.a(gate33inter0), .b(s_48), .O(gate33inter1));
  and2  gate885(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate886(.a(s_48), .O(gate33inter3));
  inv1  gate887(.a(s_49), .O(gate33inter4));
  nand2 gate888(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate889(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate890(.a(G17), .O(gate33inter7));
  inv1  gate891(.a(G21), .O(gate33inter8));
  nand2 gate892(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate893(.a(s_49), .b(gate33inter3), .O(gate33inter10));
  nor2  gate894(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate895(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate896(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2787(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2788(.a(gate34inter0), .b(s_320), .O(gate34inter1));
  and2  gate2789(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2790(.a(s_320), .O(gate34inter3));
  inv1  gate2791(.a(s_321), .O(gate34inter4));
  nand2 gate2792(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2793(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2794(.a(G25), .O(gate34inter7));
  inv1  gate2795(.a(G29), .O(gate34inter8));
  nand2 gate2796(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2797(.a(s_321), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2798(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2799(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2800(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1513(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1514(.a(gate35inter0), .b(s_138), .O(gate35inter1));
  and2  gate1515(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1516(.a(s_138), .O(gate35inter3));
  inv1  gate1517(.a(s_139), .O(gate35inter4));
  nand2 gate1518(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1519(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1520(.a(G18), .O(gate35inter7));
  inv1  gate1521(.a(G22), .O(gate35inter8));
  nand2 gate1522(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1523(.a(s_139), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1524(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1525(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1526(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1877(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1878(.a(gate36inter0), .b(s_190), .O(gate36inter1));
  and2  gate1879(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1880(.a(s_190), .O(gate36inter3));
  inv1  gate1881(.a(s_191), .O(gate36inter4));
  nand2 gate1882(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1883(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1884(.a(G26), .O(gate36inter7));
  inv1  gate1885(.a(G30), .O(gate36inter8));
  nand2 gate1886(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1887(.a(s_191), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1888(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1889(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1890(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2395(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2396(.a(gate38inter0), .b(s_264), .O(gate38inter1));
  and2  gate2397(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2398(.a(s_264), .O(gate38inter3));
  inv1  gate2399(.a(s_265), .O(gate38inter4));
  nand2 gate2400(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2401(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2402(.a(G27), .O(gate38inter7));
  inv1  gate2403(.a(G31), .O(gate38inter8));
  nand2 gate2404(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2405(.a(s_265), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2406(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2407(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2408(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate2129(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2130(.a(gate45inter0), .b(s_226), .O(gate45inter1));
  and2  gate2131(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2132(.a(s_226), .O(gate45inter3));
  inv1  gate2133(.a(s_227), .O(gate45inter4));
  nand2 gate2134(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2135(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2136(.a(G5), .O(gate45inter7));
  inv1  gate2137(.a(G272), .O(gate45inter8));
  nand2 gate2138(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2139(.a(s_227), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2140(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2141(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2142(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate841(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate842(.a(gate46inter0), .b(s_42), .O(gate46inter1));
  and2  gate843(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate844(.a(s_42), .O(gate46inter3));
  inv1  gate845(.a(s_43), .O(gate46inter4));
  nand2 gate846(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate847(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate848(.a(G6), .O(gate46inter7));
  inv1  gate849(.a(G272), .O(gate46inter8));
  nand2 gate850(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate851(.a(s_43), .b(gate46inter3), .O(gate46inter10));
  nor2  gate852(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate853(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate854(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1653(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1654(.a(gate47inter0), .b(s_158), .O(gate47inter1));
  and2  gate1655(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1656(.a(s_158), .O(gate47inter3));
  inv1  gate1657(.a(s_159), .O(gate47inter4));
  nand2 gate1658(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1659(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1660(.a(G7), .O(gate47inter7));
  inv1  gate1661(.a(G275), .O(gate47inter8));
  nand2 gate1662(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1663(.a(s_159), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1664(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1665(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1666(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2521(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2522(.a(gate49inter0), .b(s_282), .O(gate49inter1));
  and2  gate2523(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2524(.a(s_282), .O(gate49inter3));
  inv1  gate2525(.a(s_283), .O(gate49inter4));
  nand2 gate2526(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2527(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2528(.a(G9), .O(gate49inter7));
  inv1  gate2529(.a(G278), .O(gate49inter8));
  nand2 gate2530(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2531(.a(s_283), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2532(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2533(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2534(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2409(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2410(.a(gate50inter0), .b(s_266), .O(gate50inter1));
  and2  gate2411(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2412(.a(s_266), .O(gate50inter3));
  inv1  gate2413(.a(s_267), .O(gate50inter4));
  nand2 gate2414(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2415(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2416(.a(G10), .O(gate50inter7));
  inv1  gate2417(.a(G278), .O(gate50inter8));
  nand2 gate2418(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2419(.a(s_267), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2420(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2421(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2422(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1695(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1696(.a(gate52inter0), .b(s_164), .O(gate52inter1));
  and2  gate1697(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1698(.a(s_164), .O(gate52inter3));
  inv1  gate1699(.a(s_165), .O(gate52inter4));
  nand2 gate1700(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1701(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1702(.a(G12), .O(gate52inter7));
  inv1  gate1703(.a(G281), .O(gate52inter8));
  nand2 gate1704(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1705(.a(s_165), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1706(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1707(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1708(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1051(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1052(.a(gate53inter0), .b(s_72), .O(gate53inter1));
  and2  gate1053(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1054(.a(s_72), .O(gate53inter3));
  inv1  gate1055(.a(s_73), .O(gate53inter4));
  nand2 gate1056(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1057(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1058(.a(G13), .O(gate53inter7));
  inv1  gate1059(.a(G284), .O(gate53inter8));
  nand2 gate1060(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1061(.a(s_73), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1062(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1063(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1064(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1037(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1038(.a(gate54inter0), .b(s_70), .O(gate54inter1));
  and2  gate1039(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1040(.a(s_70), .O(gate54inter3));
  inv1  gate1041(.a(s_71), .O(gate54inter4));
  nand2 gate1042(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1043(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1044(.a(G14), .O(gate54inter7));
  inv1  gate1045(.a(G284), .O(gate54inter8));
  nand2 gate1046(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1047(.a(s_71), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1048(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1049(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1050(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1149(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1150(.a(gate55inter0), .b(s_86), .O(gate55inter1));
  and2  gate1151(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1152(.a(s_86), .O(gate55inter3));
  inv1  gate1153(.a(s_87), .O(gate55inter4));
  nand2 gate1154(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1155(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1156(.a(G15), .O(gate55inter7));
  inv1  gate1157(.a(G287), .O(gate55inter8));
  nand2 gate1158(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1159(.a(s_87), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1160(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1161(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1162(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate2955(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2956(.a(gate57inter0), .b(s_344), .O(gate57inter1));
  and2  gate2957(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2958(.a(s_344), .O(gate57inter3));
  inv1  gate2959(.a(s_345), .O(gate57inter4));
  nand2 gate2960(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2961(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2962(.a(G17), .O(gate57inter7));
  inv1  gate2963(.a(G290), .O(gate57inter8));
  nand2 gate2964(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2965(.a(s_345), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2966(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2967(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2968(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2507(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2508(.a(gate59inter0), .b(s_280), .O(gate59inter1));
  and2  gate2509(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2510(.a(s_280), .O(gate59inter3));
  inv1  gate2511(.a(s_281), .O(gate59inter4));
  nand2 gate2512(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2513(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2514(.a(G19), .O(gate59inter7));
  inv1  gate2515(.a(G293), .O(gate59inter8));
  nand2 gate2516(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2517(.a(s_281), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2518(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2519(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2520(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2913(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2914(.a(gate62inter0), .b(s_338), .O(gate62inter1));
  and2  gate2915(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2916(.a(s_338), .O(gate62inter3));
  inv1  gate2917(.a(s_339), .O(gate62inter4));
  nand2 gate2918(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2919(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2920(.a(G22), .O(gate62inter7));
  inv1  gate2921(.a(G296), .O(gate62inter8));
  nand2 gate2922(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2923(.a(s_339), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2924(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2925(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2926(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2535(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2536(.a(gate64inter0), .b(s_284), .O(gate64inter1));
  and2  gate2537(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2538(.a(s_284), .O(gate64inter3));
  inv1  gate2539(.a(s_285), .O(gate64inter4));
  nand2 gate2540(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2541(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2542(.a(G24), .O(gate64inter7));
  inv1  gate2543(.a(G299), .O(gate64inter8));
  nand2 gate2544(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2545(.a(s_285), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2546(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2547(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2548(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1331(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1332(.a(gate66inter0), .b(s_112), .O(gate66inter1));
  and2  gate1333(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1334(.a(s_112), .O(gate66inter3));
  inv1  gate1335(.a(s_113), .O(gate66inter4));
  nand2 gate1336(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1337(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1338(.a(G26), .O(gate66inter7));
  inv1  gate1339(.a(G302), .O(gate66inter8));
  nand2 gate1340(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1341(.a(s_113), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1342(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1343(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1344(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1415(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1416(.a(gate71inter0), .b(s_124), .O(gate71inter1));
  and2  gate1417(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1418(.a(s_124), .O(gate71inter3));
  inv1  gate1419(.a(s_125), .O(gate71inter4));
  nand2 gate1420(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1421(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1422(.a(G31), .O(gate71inter7));
  inv1  gate1423(.a(G311), .O(gate71inter8));
  nand2 gate1424(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1425(.a(s_125), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1426(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1427(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1428(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1135(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1136(.a(gate73inter0), .b(s_84), .O(gate73inter1));
  and2  gate1137(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1138(.a(s_84), .O(gate73inter3));
  inv1  gate1139(.a(s_85), .O(gate73inter4));
  nand2 gate1140(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1141(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1142(.a(G1), .O(gate73inter7));
  inv1  gate1143(.a(G314), .O(gate73inter8));
  nand2 gate1144(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1145(.a(s_85), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1146(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1147(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1148(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1555(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1556(.a(gate74inter0), .b(s_144), .O(gate74inter1));
  and2  gate1557(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1558(.a(s_144), .O(gate74inter3));
  inv1  gate1559(.a(s_145), .O(gate74inter4));
  nand2 gate1560(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1561(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1562(.a(G5), .O(gate74inter7));
  inv1  gate1563(.a(G314), .O(gate74inter8));
  nand2 gate1564(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1565(.a(s_145), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1566(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1567(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1568(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate2325(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2326(.a(gate75inter0), .b(s_254), .O(gate75inter1));
  and2  gate2327(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2328(.a(s_254), .O(gate75inter3));
  inv1  gate2329(.a(s_255), .O(gate75inter4));
  nand2 gate2330(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2331(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2332(.a(G9), .O(gate75inter7));
  inv1  gate2333(.a(G317), .O(gate75inter8));
  nand2 gate2334(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2335(.a(s_255), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2336(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2337(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2338(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1247(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1248(.a(gate79inter0), .b(s_100), .O(gate79inter1));
  and2  gate1249(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1250(.a(s_100), .O(gate79inter3));
  inv1  gate1251(.a(s_101), .O(gate79inter4));
  nand2 gate1252(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1253(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1254(.a(G10), .O(gate79inter7));
  inv1  gate1255(.a(G323), .O(gate79inter8));
  nand2 gate1256(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1257(.a(s_101), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1258(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1259(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1260(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate981(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate982(.a(gate80inter0), .b(s_62), .O(gate80inter1));
  and2  gate983(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate984(.a(s_62), .O(gate80inter3));
  inv1  gate985(.a(s_63), .O(gate80inter4));
  nand2 gate986(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate987(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate988(.a(G14), .O(gate80inter7));
  inv1  gate989(.a(G323), .O(gate80inter8));
  nand2 gate990(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate991(.a(s_63), .b(gate80inter3), .O(gate80inter10));
  nor2  gate992(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate993(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate994(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1401(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1402(.a(gate82inter0), .b(s_122), .O(gate82inter1));
  and2  gate1403(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1404(.a(s_122), .O(gate82inter3));
  inv1  gate1405(.a(s_123), .O(gate82inter4));
  nand2 gate1406(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1407(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1408(.a(G7), .O(gate82inter7));
  inv1  gate1409(.a(G326), .O(gate82inter8));
  nand2 gate1410(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1411(.a(s_123), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1412(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1413(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1414(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate645(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate646(.a(gate86inter0), .b(s_14), .O(gate86inter1));
  and2  gate647(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate648(.a(s_14), .O(gate86inter3));
  inv1  gate649(.a(s_15), .O(gate86inter4));
  nand2 gate650(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate651(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate652(.a(G8), .O(gate86inter7));
  inv1  gate653(.a(G332), .O(gate86inter8));
  nand2 gate654(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate655(.a(s_15), .b(gate86inter3), .O(gate86inter10));
  nor2  gate656(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate657(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate658(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1527(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1528(.a(gate87inter0), .b(s_140), .O(gate87inter1));
  and2  gate1529(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1530(.a(s_140), .O(gate87inter3));
  inv1  gate1531(.a(s_141), .O(gate87inter4));
  nand2 gate1532(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1533(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1534(.a(G12), .O(gate87inter7));
  inv1  gate1535(.a(G335), .O(gate87inter8));
  nand2 gate1536(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1537(.a(s_141), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1538(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1539(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1540(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2731(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2732(.a(gate90inter0), .b(s_312), .O(gate90inter1));
  and2  gate2733(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2734(.a(s_312), .O(gate90inter3));
  inv1  gate2735(.a(s_313), .O(gate90inter4));
  nand2 gate2736(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2737(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2738(.a(G21), .O(gate90inter7));
  inv1  gate2739(.a(G338), .O(gate90inter8));
  nand2 gate2740(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2741(.a(s_313), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2742(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2743(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2744(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate3179(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate3180(.a(gate94inter0), .b(s_376), .O(gate94inter1));
  and2  gate3181(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate3182(.a(s_376), .O(gate94inter3));
  inv1  gate3183(.a(s_377), .O(gate94inter4));
  nand2 gate3184(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate3185(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate3186(.a(G22), .O(gate94inter7));
  inv1  gate3187(.a(G344), .O(gate94inter8));
  nand2 gate3188(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate3189(.a(s_377), .b(gate94inter3), .O(gate94inter10));
  nor2  gate3190(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate3191(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate3192(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate3137(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate3138(.a(gate95inter0), .b(s_370), .O(gate95inter1));
  and2  gate3139(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate3140(.a(s_370), .O(gate95inter3));
  inv1  gate3141(.a(s_371), .O(gate95inter4));
  nand2 gate3142(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate3143(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate3144(.a(G26), .O(gate95inter7));
  inv1  gate3145(.a(G347), .O(gate95inter8));
  nand2 gate3146(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate3147(.a(s_371), .b(gate95inter3), .O(gate95inter10));
  nor2  gate3148(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate3149(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate3150(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate659(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate660(.a(gate96inter0), .b(s_16), .O(gate96inter1));
  and2  gate661(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate662(.a(s_16), .O(gate96inter3));
  inv1  gate663(.a(s_17), .O(gate96inter4));
  nand2 gate664(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate665(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate666(.a(G30), .O(gate96inter7));
  inv1  gate667(.a(G347), .O(gate96inter8));
  nand2 gate668(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate669(.a(s_17), .b(gate96inter3), .O(gate96inter10));
  nor2  gate670(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate671(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate672(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2983(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2984(.a(gate97inter0), .b(s_348), .O(gate97inter1));
  and2  gate2985(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2986(.a(s_348), .O(gate97inter3));
  inv1  gate2987(.a(s_349), .O(gate97inter4));
  nand2 gate2988(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2989(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2990(.a(G19), .O(gate97inter7));
  inv1  gate2991(.a(G350), .O(gate97inter8));
  nand2 gate2992(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2993(.a(s_349), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2994(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2995(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2996(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1989(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1990(.a(gate99inter0), .b(s_206), .O(gate99inter1));
  and2  gate1991(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1992(.a(s_206), .O(gate99inter3));
  inv1  gate1993(.a(s_207), .O(gate99inter4));
  nand2 gate1994(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1995(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1996(.a(G27), .O(gate99inter7));
  inv1  gate1997(.a(G353), .O(gate99inter8));
  nand2 gate1998(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1999(.a(s_207), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2000(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2001(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2002(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2241(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2242(.a(gate102inter0), .b(s_242), .O(gate102inter1));
  and2  gate2243(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2244(.a(s_242), .O(gate102inter3));
  inv1  gate2245(.a(s_243), .O(gate102inter4));
  nand2 gate2246(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2247(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2248(.a(G24), .O(gate102inter7));
  inv1  gate2249(.a(G356), .O(gate102inter8));
  nand2 gate2250(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2251(.a(s_243), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2252(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2253(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2254(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate3067(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate3068(.a(gate105inter0), .b(s_360), .O(gate105inter1));
  and2  gate3069(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate3070(.a(s_360), .O(gate105inter3));
  inv1  gate3071(.a(s_361), .O(gate105inter4));
  nand2 gate3072(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate3073(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate3074(.a(G362), .O(gate105inter7));
  inv1  gate3075(.a(G363), .O(gate105inter8));
  nand2 gate3076(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate3077(.a(s_361), .b(gate105inter3), .O(gate105inter10));
  nor2  gate3078(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate3079(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate3080(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1387(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1388(.a(gate108inter0), .b(s_120), .O(gate108inter1));
  and2  gate1389(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1390(.a(s_120), .O(gate108inter3));
  inv1  gate1391(.a(s_121), .O(gate108inter4));
  nand2 gate1392(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1393(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1394(.a(G368), .O(gate108inter7));
  inv1  gate1395(.a(G369), .O(gate108inter8));
  nand2 gate1396(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1397(.a(s_121), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1398(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1399(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1400(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1709(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1710(.a(gate109inter0), .b(s_166), .O(gate109inter1));
  and2  gate1711(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1712(.a(s_166), .O(gate109inter3));
  inv1  gate1713(.a(s_167), .O(gate109inter4));
  nand2 gate1714(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1715(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1716(.a(G370), .O(gate109inter7));
  inv1  gate1717(.a(G371), .O(gate109inter8));
  nand2 gate1718(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1719(.a(s_167), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1720(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1721(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1722(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate995(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate996(.a(gate110inter0), .b(s_64), .O(gate110inter1));
  and2  gate997(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate998(.a(s_64), .O(gate110inter3));
  inv1  gate999(.a(s_65), .O(gate110inter4));
  nand2 gate1000(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1001(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1002(.a(G372), .O(gate110inter7));
  inv1  gate1003(.a(G373), .O(gate110inter8));
  nand2 gate1004(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1005(.a(s_65), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1006(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1007(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1008(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2871(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2872(.a(gate112inter0), .b(s_332), .O(gate112inter1));
  and2  gate2873(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2874(.a(s_332), .O(gate112inter3));
  inv1  gate2875(.a(s_333), .O(gate112inter4));
  nand2 gate2876(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2877(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2878(.a(G376), .O(gate112inter7));
  inv1  gate2879(.a(G377), .O(gate112inter8));
  nand2 gate2880(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2881(.a(s_333), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2882(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2883(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2884(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate589(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate590(.a(gate115inter0), .b(s_6), .O(gate115inter1));
  and2  gate591(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate592(.a(s_6), .O(gate115inter3));
  inv1  gate593(.a(s_7), .O(gate115inter4));
  nand2 gate594(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate595(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate596(.a(G382), .O(gate115inter7));
  inv1  gate597(.a(G383), .O(gate115inter8));
  nand2 gate598(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate599(.a(s_7), .b(gate115inter3), .O(gate115inter10));
  nor2  gate600(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate601(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate602(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1443(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1444(.a(gate120inter0), .b(s_128), .O(gate120inter1));
  and2  gate1445(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1446(.a(s_128), .O(gate120inter3));
  inv1  gate1447(.a(s_129), .O(gate120inter4));
  nand2 gate1448(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1449(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1450(.a(G392), .O(gate120inter7));
  inv1  gate1451(.a(G393), .O(gate120inter8));
  nand2 gate1452(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1453(.a(s_129), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1454(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1455(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1456(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2451(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2452(.a(gate125inter0), .b(s_272), .O(gate125inter1));
  and2  gate2453(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2454(.a(s_272), .O(gate125inter3));
  inv1  gate2455(.a(s_273), .O(gate125inter4));
  nand2 gate2456(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2457(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2458(.a(G402), .O(gate125inter7));
  inv1  gate2459(.a(G403), .O(gate125inter8));
  nand2 gate2460(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2461(.a(s_273), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2462(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2463(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2464(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate785(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate786(.a(gate128inter0), .b(s_34), .O(gate128inter1));
  and2  gate787(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate788(.a(s_34), .O(gate128inter3));
  inv1  gate789(.a(s_35), .O(gate128inter4));
  nand2 gate790(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate791(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate792(.a(G408), .O(gate128inter7));
  inv1  gate793(.a(G409), .O(gate128inter8));
  nand2 gate794(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate795(.a(s_35), .b(gate128inter3), .O(gate128inter10));
  nor2  gate796(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate797(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate798(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate3095(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate3096(.a(gate130inter0), .b(s_364), .O(gate130inter1));
  and2  gate3097(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate3098(.a(s_364), .O(gate130inter3));
  inv1  gate3099(.a(s_365), .O(gate130inter4));
  nand2 gate3100(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate3101(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate3102(.a(G412), .O(gate130inter7));
  inv1  gate3103(.a(G413), .O(gate130inter8));
  nand2 gate3104(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate3105(.a(s_365), .b(gate130inter3), .O(gate130inter10));
  nor2  gate3106(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate3107(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate3108(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate3109(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate3110(.a(gate131inter0), .b(s_366), .O(gate131inter1));
  and2  gate3111(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate3112(.a(s_366), .O(gate131inter3));
  inv1  gate3113(.a(s_367), .O(gate131inter4));
  nand2 gate3114(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate3115(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate3116(.a(G414), .O(gate131inter7));
  inv1  gate3117(.a(G415), .O(gate131inter8));
  nand2 gate3118(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate3119(.a(s_367), .b(gate131inter3), .O(gate131inter10));
  nor2  gate3120(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate3121(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate3122(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate3151(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate3152(.a(gate132inter0), .b(s_372), .O(gate132inter1));
  and2  gate3153(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate3154(.a(s_372), .O(gate132inter3));
  inv1  gate3155(.a(s_373), .O(gate132inter4));
  nand2 gate3156(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate3157(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate3158(.a(G416), .O(gate132inter7));
  inv1  gate3159(.a(G417), .O(gate132inter8));
  nand2 gate3160(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate3161(.a(s_373), .b(gate132inter3), .O(gate132inter10));
  nor2  gate3162(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate3163(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate3164(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1807(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1808(.a(gate133inter0), .b(s_180), .O(gate133inter1));
  and2  gate1809(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1810(.a(s_180), .O(gate133inter3));
  inv1  gate1811(.a(s_181), .O(gate133inter4));
  nand2 gate1812(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1813(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1814(.a(G418), .O(gate133inter7));
  inv1  gate1815(.a(G419), .O(gate133inter8));
  nand2 gate1816(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1817(.a(s_181), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1818(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1819(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1820(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate2087(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2088(.a(gate134inter0), .b(s_220), .O(gate134inter1));
  and2  gate2089(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2090(.a(s_220), .O(gate134inter3));
  inv1  gate2091(.a(s_221), .O(gate134inter4));
  nand2 gate2092(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2093(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2094(.a(G420), .O(gate134inter7));
  inv1  gate2095(.a(G421), .O(gate134inter8));
  nand2 gate2096(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2097(.a(s_221), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2098(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2099(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2100(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2311(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2312(.a(gate140inter0), .b(s_252), .O(gate140inter1));
  and2  gate2313(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2314(.a(s_252), .O(gate140inter3));
  inv1  gate2315(.a(s_253), .O(gate140inter4));
  nand2 gate2316(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2317(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2318(.a(G444), .O(gate140inter7));
  inv1  gate2319(.a(G447), .O(gate140inter8));
  nand2 gate2320(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2321(.a(s_253), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2322(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2323(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2324(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate799(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate800(.a(gate141inter0), .b(s_36), .O(gate141inter1));
  and2  gate801(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate802(.a(s_36), .O(gate141inter3));
  inv1  gate803(.a(s_37), .O(gate141inter4));
  nand2 gate804(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate805(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate806(.a(G450), .O(gate141inter7));
  inv1  gate807(.a(G453), .O(gate141inter8));
  nand2 gate808(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate809(.a(s_37), .b(gate141inter3), .O(gate141inter10));
  nor2  gate810(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate811(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate812(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2745(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2746(.a(gate144inter0), .b(s_314), .O(gate144inter1));
  and2  gate2747(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2748(.a(s_314), .O(gate144inter3));
  inv1  gate2749(.a(s_315), .O(gate144inter4));
  nand2 gate2750(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2751(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2752(.a(G468), .O(gate144inter7));
  inv1  gate2753(.a(G471), .O(gate144inter8));
  nand2 gate2754(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2755(.a(s_315), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2756(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2757(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2758(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate561(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate562(.a(gate146inter0), .b(s_2), .O(gate146inter1));
  and2  gate563(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate564(.a(s_2), .O(gate146inter3));
  inv1  gate565(.a(s_3), .O(gate146inter4));
  nand2 gate566(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate567(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate568(.a(G480), .O(gate146inter7));
  inv1  gate569(.a(G483), .O(gate146inter8));
  nand2 gate570(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate571(.a(s_3), .b(gate146inter3), .O(gate146inter10));
  nor2  gate572(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate573(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate574(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2801(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2802(.a(gate148inter0), .b(s_322), .O(gate148inter1));
  and2  gate2803(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2804(.a(s_322), .O(gate148inter3));
  inv1  gate2805(.a(s_323), .O(gate148inter4));
  nand2 gate2806(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2807(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2808(.a(G492), .O(gate148inter7));
  inv1  gate2809(.a(G495), .O(gate148inter8));
  nand2 gate2810(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2811(.a(s_323), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2812(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2813(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2814(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate2227(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2228(.a(gate149inter0), .b(s_240), .O(gate149inter1));
  and2  gate2229(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2230(.a(s_240), .O(gate149inter3));
  inv1  gate2231(.a(s_241), .O(gate149inter4));
  nand2 gate2232(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2233(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2234(.a(G498), .O(gate149inter7));
  inv1  gate2235(.a(G501), .O(gate149inter8));
  nand2 gate2236(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2237(.a(s_241), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2238(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2239(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2240(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2703(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2704(.a(gate150inter0), .b(s_308), .O(gate150inter1));
  and2  gate2705(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2706(.a(s_308), .O(gate150inter3));
  inv1  gate2707(.a(s_309), .O(gate150inter4));
  nand2 gate2708(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2709(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2710(.a(G504), .O(gate150inter7));
  inv1  gate2711(.a(G507), .O(gate150inter8));
  nand2 gate2712(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2713(.a(s_309), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2714(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2715(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2716(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate939(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate940(.a(gate151inter0), .b(s_56), .O(gate151inter1));
  and2  gate941(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate942(.a(s_56), .O(gate151inter3));
  inv1  gate943(.a(s_57), .O(gate151inter4));
  nand2 gate944(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate945(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate946(.a(G510), .O(gate151inter7));
  inv1  gate947(.a(G513), .O(gate151inter8));
  nand2 gate948(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate949(.a(s_57), .b(gate151inter3), .O(gate151inter10));
  nor2  gate950(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate951(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate952(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1317(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1318(.a(gate153inter0), .b(s_110), .O(gate153inter1));
  and2  gate1319(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1320(.a(s_110), .O(gate153inter3));
  inv1  gate1321(.a(s_111), .O(gate153inter4));
  nand2 gate1322(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1323(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1324(.a(G426), .O(gate153inter7));
  inv1  gate1325(.a(G522), .O(gate153inter8));
  nand2 gate1326(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1327(.a(s_111), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1328(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1329(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1330(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate3277(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate3278(.a(gate154inter0), .b(s_390), .O(gate154inter1));
  and2  gate3279(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate3280(.a(s_390), .O(gate154inter3));
  inv1  gate3281(.a(s_391), .O(gate154inter4));
  nand2 gate3282(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate3283(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate3284(.a(G429), .O(gate154inter7));
  inv1  gate3285(.a(G522), .O(gate154inter8));
  nand2 gate3286(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate3287(.a(s_391), .b(gate154inter3), .O(gate154inter10));
  nor2  gate3288(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate3289(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate3290(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2255(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2256(.a(gate155inter0), .b(s_244), .O(gate155inter1));
  and2  gate2257(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2258(.a(s_244), .O(gate155inter3));
  inv1  gate2259(.a(s_245), .O(gate155inter4));
  nand2 gate2260(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2261(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2262(.a(G432), .O(gate155inter7));
  inv1  gate2263(.a(G525), .O(gate155inter8));
  nand2 gate2264(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2265(.a(s_245), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2266(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2267(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2268(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2857(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2858(.a(gate156inter0), .b(s_330), .O(gate156inter1));
  and2  gate2859(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2860(.a(s_330), .O(gate156inter3));
  inv1  gate2861(.a(s_331), .O(gate156inter4));
  nand2 gate2862(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2863(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2864(.a(G435), .O(gate156inter7));
  inv1  gate2865(.a(G525), .O(gate156inter8));
  nand2 gate2866(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2867(.a(s_331), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2868(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2869(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2870(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2773(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2774(.a(gate161inter0), .b(s_318), .O(gate161inter1));
  and2  gate2775(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2776(.a(s_318), .O(gate161inter3));
  inv1  gate2777(.a(s_319), .O(gate161inter4));
  nand2 gate2778(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2779(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2780(.a(G450), .O(gate161inter7));
  inv1  gate2781(.a(G534), .O(gate161inter8));
  nand2 gate2782(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2783(.a(s_319), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2784(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2785(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2786(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate2143(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2144(.a(gate163inter0), .b(s_228), .O(gate163inter1));
  and2  gate2145(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2146(.a(s_228), .O(gate163inter3));
  inv1  gate2147(.a(s_229), .O(gate163inter4));
  nand2 gate2148(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2149(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2150(.a(G456), .O(gate163inter7));
  inv1  gate2151(.a(G537), .O(gate163inter8));
  nand2 gate2152(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2153(.a(s_229), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2154(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2155(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2156(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1429(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1430(.a(gate164inter0), .b(s_126), .O(gate164inter1));
  and2  gate1431(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1432(.a(s_126), .O(gate164inter3));
  inv1  gate1433(.a(s_127), .O(gate164inter4));
  nand2 gate1434(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1435(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1436(.a(G459), .O(gate164inter7));
  inv1  gate1437(.a(G537), .O(gate164inter8));
  nand2 gate1438(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1439(.a(s_127), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1440(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1441(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1442(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2619(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2620(.a(gate168inter0), .b(s_296), .O(gate168inter1));
  and2  gate2621(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2622(.a(s_296), .O(gate168inter3));
  inv1  gate2623(.a(s_297), .O(gate168inter4));
  nand2 gate2624(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2625(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2626(.a(G471), .O(gate168inter7));
  inv1  gate2627(.a(G543), .O(gate168inter8));
  nand2 gate2628(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2629(.a(s_297), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2630(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2631(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2632(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1597(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1598(.a(gate169inter0), .b(s_150), .O(gate169inter1));
  and2  gate1599(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1600(.a(s_150), .O(gate169inter3));
  inv1  gate1601(.a(s_151), .O(gate169inter4));
  nand2 gate1602(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1603(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1604(.a(G474), .O(gate169inter7));
  inv1  gate1605(.a(G546), .O(gate169inter8));
  nand2 gate1606(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1607(.a(s_151), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1608(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1609(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1610(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate575(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate576(.a(gate170inter0), .b(s_4), .O(gate170inter1));
  and2  gate577(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate578(.a(s_4), .O(gate170inter3));
  inv1  gate579(.a(s_5), .O(gate170inter4));
  nand2 gate580(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate581(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate582(.a(G477), .O(gate170inter7));
  inv1  gate583(.a(G546), .O(gate170inter8));
  nand2 gate584(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate585(.a(s_5), .b(gate170inter3), .O(gate170inter10));
  nor2  gate586(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate587(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate588(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1107(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1108(.a(gate176inter0), .b(s_80), .O(gate176inter1));
  and2  gate1109(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1110(.a(s_80), .O(gate176inter3));
  inv1  gate1111(.a(s_81), .O(gate176inter4));
  nand2 gate1112(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1113(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1114(.a(G495), .O(gate176inter7));
  inv1  gate1115(.a(G555), .O(gate176inter8));
  nand2 gate1116(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1117(.a(s_81), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1118(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1119(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1120(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2689(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2690(.a(gate179inter0), .b(s_306), .O(gate179inter1));
  and2  gate2691(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2692(.a(s_306), .O(gate179inter3));
  inv1  gate2693(.a(s_307), .O(gate179inter4));
  nand2 gate2694(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2695(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2696(.a(G504), .O(gate179inter7));
  inv1  gate2697(.a(G561), .O(gate179inter8));
  nand2 gate2698(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2699(.a(s_307), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2700(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2701(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2702(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1499(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1500(.a(gate180inter0), .b(s_136), .O(gate180inter1));
  and2  gate1501(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1502(.a(s_136), .O(gate180inter3));
  inv1  gate1503(.a(s_137), .O(gate180inter4));
  nand2 gate1504(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1505(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1506(.a(G507), .O(gate180inter7));
  inv1  gate1507(.a(G561), .O(gate180inter8));
  nand2 gate1508(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1509(.a(s_137), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1510(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1511(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1512(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate2339(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2340(.a(gate181inter0), .b(s_256), .O(gate181inter1));
  and2  gate2341(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2342(.a(s_256), .O(gate181inter3));
  inv1  gate2343(.a(s_257), .O(gate181inter4));
  nand2 gate2344(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2345(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2346(.a(G510), .O(gate181inter7));
  inv1  gate2347(.a(G564), .O(gate181inter8));
  nand2 gate2348(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2349(.a(s_257), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2350(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2351(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2352(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate3263(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate3264(.a(gate184inter0), .b(s_388), .O(gate184inter1));
  and2  gate3265(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate3266(.a(s_388), .O(gate184inter3));
  inv1  gate3267(.a(s_389), .O(gate184inter4));
  nand2 gate3268(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate3269(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate3270(.a(G519), .O(gate184inter7));
  inv1  gate3271(.a(G567), .O(gate184inter8));
  nand2 gate3272(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate3273(.a(s_389), .b(gate184inter3), .O(gate184inter10));
  nor2  gate3274(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate3275(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate3276(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate3039(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate3040(.a(gate188inter0), .b(s_356), .O(gate188inter1));
  and2  gate3041(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate3042(.a(s_356), .O(gate188inter3));
  inv1  gate3043(.a(s_357), .O(gate188inter4));
  nand2 gate3044(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate3045(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate3046(.a(G576), .O(gate188inter7));
  inv1  gate3047(.a(G577), .O(gate188inter8));
  nand2 gate3048(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate3049(.a(s_357), .b(gate188inter3), .O(gate188inter10));
  nor2  gate3050(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate3051(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate3052(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1261(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1262(.a(gate189inter0), .b(s_102), .O(gate189inter1));
  and2  gate1263(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1264(.a(s_102), .O(gate189inter3));
  inv1  gate1265(.a(s_103), .O(gate189inter4));
  nand2 gate1266(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1267(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1268(.a(G578), .O(gate189inter7));
  inv1  gate1269(.a(G579), .O(gate189inter8));
  nand2 gate1270(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1271(.a(s_103), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1272(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1273(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1274(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1947(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1948(.a(gate190inter0), .b(s_200), .O(gate190inter1));
  and2  gate1949(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1950(.a(s_200), .O(gate190inter3));
  inv1  gate1951(.a(s_201), .O(gate190inter4));
  nand2 gate1952(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1953(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1954(.a(G580), .O(gate190inter7));
  inv1  gate1955(.a(G581), .O(gate190inter8));
  nand2 gate1956(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1957(.a(s_201), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1958(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1959(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1960(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate687(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate688(.a(gate193inter0), .b(s_20), .O(gate193inter1));
  and2  gate689(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate690(.a(s_20), .O(gate193inter3));
  inv1  gate691(.a(s_21), .O(gate193inter4));
  nand2 gate692(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate693(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate694(.a(G586), .O(gate193inter7));
  inv1  gate695(.a(G587), .O(gate193inter8));
  nand2 gate696(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate697(.a(s_21), .b(gate193inter3), .O(gate193inter10));
  nor2  gate698(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate699(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate700(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2675(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2676(.a(gate195inter0), .b(s_304), .O(gate195inter1));
  and2  gate2677(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2678(.a(s_304), .O(gate195inter3));
  inv1  gate2679(.a(s_305), .O(gate195inter4));
  nand2 gate2680(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2681(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2682(.a(G590), .O(gate195inter7));
  inv1  gate2683(.a(G591), .O(gate195inter8));
  nand2 gate2684(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2685(.a(s_305), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2686(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2687(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2688(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate631(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate632(.a(gate196inter0), .b(s_12), .O(gate196inter1));
  and2  gate633(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate634(.a(s_12), .O(gate196inter3));
  inv1  gate635(.a(s_13), .O(gate196inter4));
  nand2 gate636(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate637(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate638(.a(G592), .O(gate196inter7));
  inv1  gate639(.a(G593), .O(gate196inter8));
  nand2 gate640(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate641(.a(s_13), .b(gate196inter3), .O(gate196inter10));
  nor2  gate642(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate643(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate644(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2059(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2060(.a(gate198inter0), .b(s_216), .O(gate198inter1));
  and2  gate2061(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2062(.a(s_216), .O(gate198inter3));
  inv1  gate2063(.a(s_217), .O(gate198inter4));
  nand2 gate2064(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2065(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2066(.a(G596), .O(gate198inter7));
  inv1  gate2067(.a(G597), .O(gate198inter8));
  nand2 gate2068(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2069(.a(s_217), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2070(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2071(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2072(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1961(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1962(.a(gate199inter0), .b(s_202), .O(gate199inter1));
  and2  gate1963(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1964(.a(s_202), .O(gate199inter3));
  inv1  gate1965(.a(s_203), .O(gate199inter4));
  nand2 gate1966(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1967(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1968(.a(G598), .O(gate199inter7));
  inv1  gate1969(.a(G599), .O(gate199inter8));
  nand2 gate1970(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1971(.a(s_203), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1972(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1973(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1974(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate617(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate618(.a(gate200inter0), .b(s_10), .O(gate200inter1));
  and2  gate619(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate620(.a(s_10), .O(gate200inter3));
  inv1  gate621(.a(s_11), .O(gate200inter4));
  nand2 gate622(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate623(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate624(.a(G600), .O(gate200inter7));
  inv1  gate625(.a(G601), .O(gate200inter8));
  nand2 gate626(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate627(.a(s_11), .b(gate200inter3), .O(gate200inter10));
  nor2  gate628(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate629(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate630(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1485(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1486(.a(gate203inter0), .b(s_134), .O(gate203inter1));
  and2  gate1487(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1488(.a(s_134), .O(gate203inter3));
  inv1  gate1489(.a(s_135), .O(gate203inter4));
  nand2 gate1490(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1491(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1492(.a(G602), .O(gate203inter7));
  inv1  gate1493(.a(G612), .O(gate203inter8));
  nand2 gate1494(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1495(.a(s_135), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1496(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1497(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1498(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1289(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1290(.a(gate205inter0), .b(s_106), .O(gate205inter1));
  and2  gate1291(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1292(.a(s_106), .O(gate205inter3));
  inv1  gate1293(.a(s_107), .O(gate205inter4));
  nand2 gate1294(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1295(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1296(.a(G622), .O(gate205inter7));
  inv1  gate1297(.a(G627), .O(gate205inter8));
  nand2 gate1298(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1299(.a(s_107), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1300(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1301(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1302(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1765(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1766(.a(gate206inter0), .b(s_174), .O(gate206inter1));
  and2  gate1767(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1768(.a(s_174), .O(gate206inter3));
  inv1  gate1769(.a(s_175), .O(gate206inter4));
  nand2 gate1770(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1771(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1772(.a(G632), .O(gate206inter7));
  inv1  gate1773(.a(G637), .O(gate206inter8));
  nand2 gate1774(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1775(.a(s_175), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1776(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1777(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1778(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1793(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1794(.a(gate208inter0), .b(s_178), .O(gate208inter1));
  and2  gate1795(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1796(.a(s_178), .O(gate208inter3));
  inv1  gate1797(.a(s_179), .O(gate208inter4));
  nand2 gate1798(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1799(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1800(.a(G627), .O(gate208inter7));
  inv1  gate1801(.a(G637), .O(gate208inter8));
  nand2 gate1802(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1803(.a(s_179), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1804(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1805(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1806(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2577(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2578(.a(gate209inter0), .b(s_290), .O(gate209inter1));
  and2  gate2579(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2580(.a(s_290), .O(gate209inter3));
  inv1  gate2581(.a(s_291), .O(gate209inter4));
  nand2 gate2582(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2583(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2584(.a(G602), .O(gate209inter7));
  inv1  gate2585(.a(G666), .O(gate209inter8));
  nand2 gate2586(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2587(.a(s_291), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2588(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2589(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2590(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1023(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1024(.a(gate212inter0), .b(s_68), .O(gate212inter1));
  and2  gate1025(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1026(.a(s_68), .O(gate212inter3));
  inv1  gate1027(.a(s_69), .O(gate212inter4));
  nand2 gate1028(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1029(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1030(.a(G617), .O(gate212inter7));
  inv1  gate1031(.a(G669), .O(gate212inter8));
  nand2 gate1032(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1033(.a(s_69), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1034(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1035(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1036(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1779(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1780(.a(gate214inter0), .b(s_176), .O(gate214inter1));
  and2  gate1781(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1782(.a(s_176), .O(gate214inter3));
  inv1  gate1783(.a(s_177), .O(gate214inter4));
  nand2 gate1784(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1785(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1786(.a(G612), .O(gate214inter7));
  inv1  gate1787(.a(G672), .O(gate214inter8));
  nand2 gate1788(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1789(.a(s_177), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1790(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1791(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1792(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2591(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2592(.a(gate215inter0), .b(s_292), .O(gate215inter1));
  and2  gate2593(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2594(.a(s_292), .O(gate215inter3));
  inv1  gate2595(.a(s_293), .O(gate215inter4));
  nand2 gate2596(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2597(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2598(.a(G607), .O(gate215inter7));
  inv1  gate2599(.a(G675), .O(gate215inter8));
  nand2 gate2600(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2601(.a(s_293), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2602(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2603(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2604(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate967(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate968(.a(gate216inter0), .b(s_60), .O(gate216inter1));
  and2  gate969(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate970(.a(s_60), .O(gate216inter3));
  inv1  gate971(.a(s_61), .O(gate216inter4));
  nand2 gate972(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate973(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate974(.a(G617), .O(gate216inter7));
  inv1  gate975(.a(G675), .O(gate216inter8));
  nand2 gate976(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate977(.a(s_61), .b(gate216inter3), .O(gate216inter10));
  nor2  gate978(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate979(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate980(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate3025(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate3026(.a(gate217inter0), .b(s_354), .O(gate217inter1));
  and2  gate3027(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate3028(.a(s_354), .O(gate217inter3));
  inv1  gate3029(.a(s_355), .O(gate217inter4));
  nand2 gate3030(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate3031(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate3032(.a(G622), .O(gate217inter7));
  inv1  gate3033(.a(G678), .O(gate217inter8));
  nand2 gate3034(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate3035(.a(s_355), .b(gate217inter3), .O(gate217inter10));
  nor2  gate3036(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate3037(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate3038(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2017(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2018(.a(gate220inter0), .b(s_210), .O(gate220inter1));
  and2  gate2019(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2020(.a(s_210), .O(gate220inter3));
  inv1  gate2021(.a(s_211), .O(gate220inter4));
  nand2 gate2022(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2023(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2024(.a(G637), .O(gate220inter7));
  inv1  gate2025(.a(G681), .O(gate220inter8));
  nand2 gate2026(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2027(.a(s_211), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2028(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2029(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2030(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1933(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1934(.a(gate221inter0), .b(s_198), .O(gate221inter1));
  and2  gate1935(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1936(.a(s_198), .O(gate221inter3));
  inv1  gate1937(.a(s_199), .O(gate221inter4));
  nand2 gate1938(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1939(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1940(.a(G622), .O(gate221inter7));
  inv1  gate1941(.a(G684), .O(gate221inter8));
  nand2 gate1942(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1943(.a(s_199), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1944(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1945(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1946(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1737(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1738(.a(gate229inter0), .b(s_170), .O(gate229inter1));
  and2  gate1739(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1740(.a(s_170), .O(gate229inter3));
  inv1  gate1741(.a(s_171), .O(gate229inter4));
  nand2 gate1742(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1743(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1744(.a(G698), .O(gate229inter7));
  inv1  gate1745(.a(G699), .O(gate229inter8));
  nand2 gate1746(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1747(.a(s_171), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1748(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1749(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1750(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2549(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2550(.a(gate231inter0), .b(s_286), .O(gate231inter1));
  and2  gate2551(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2552(.a(s_286), .O(gate231inter3));
  inv1  gate2553(.a(s_287), .O(gate231inter4));
  nand2 gate2554(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2555(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2556(.a(G702), .O(gate231inter7));
  inv1  gate2557(.a(G703), .O(gate231inter8));
  nand2 gate2558(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2559(.a(s_287), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2560(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2561(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2562(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1751(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1752(.a(gate234inter0), .b(s_172), .O(gate234inter1));
  and2  gate1753(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1754(.a(s_172), .O(gate234inter3));
  inv1  gate1755(.a(s_173), .O(gate234inter4));
  nand2 gate1756(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1757(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1758(.a(G245), .O(gate234inter7));
  inv1  gate1759(.a(G721), .O(gate234inter8));
  nand2 gate1760(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1761(.a(s_173), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1762(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1763(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1764(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate925(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate926(.a(gate236inter0), .b(s_54), .O(gate236inter1));
  and2  gate927(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate928(.a(s_54), .O(gate236inter3));
  inv1  gate929(.a(s_55), .O(gate236inter4));
  nand2 gate930(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate931(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate932(.a(G251), .O(gate236inter7));
  inv1  gate933(.a(G727), .O(gate236inter8));
  nand2 gate934(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate935(.a(s_55), .b(gate236inter3), .O(gate236inter10));
  nor2  gate936(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate937(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate938(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1975(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1976(.a(gate237inter0), .b(s_204), .O(gate237inter1));
  and2  gate1977(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1978(.a(s_204), .O(gate237inter3));
  inv1  gate1979(.a(s_205), .O(gate237inter4));
  nand2 gate1980(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1981(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1982(.a(G254), .O(gate237inter7));
  inv1  gate1983(.a(G706), .O(gate237inter8));
  nand2 gate1984(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1985(.a(s_205), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1986(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1987(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1988(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate2031(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate2032(.a(gate238inter0), .b(s_212), .O(gate238inter1));
  and2  gate2033(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate2034(.a(s_212), .O(gate238inter3));
  inv1  gate2035(.a(s_213), .O(gate238inter4));
  nand2 gate2036(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate2037(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate2038(.a(G257), .O(gate238inter7));
  inv1  gate2039(.a(G709), .O(gate238inter8));
  nand2 gate2040(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate2041(.a(s_213), .b(gate238inter3), .O(gate238inter10));
  nor2  gate2042(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate2043(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate2044(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2269(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2270(.a(gate242inter0), .b(s_246), .O(gate242inter1));
  and2  gate2271(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2272(.a(s_246), .O(gate242inter3));
  inv1  gate2273(.a(s_247), .O(gate242inter4));
  nand2 gate2274(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2275(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2276(.a(G718), .O(gate242inter7));
  inv1  gate2277(.a(G730), .O(gate242inter8));
  nand2 gate2278(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2279(.a(s_247), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2280(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2281(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2282(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate603(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate604(.a(gate244inter0), .b(s_8), .O(gate244inter1));
  and2  gate605(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate606(.a(s_8), .O(gate244inter3));
  inv1  gate607(.a(s_9), .O(gate244inter4));
  nand2 gate608(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate609(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate610(.a(G721), .O(gate244inter7));
  inv1  gate611(.a(G733), .O(gate244inter8));
  nand2 gate612(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate613(.a(s_9), .b(gate244inter3), .O(gate244inter10));
  nor2  gate614(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate615(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate616(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2661(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2662(.a(gate246inter0), .b(s_302), .O(gate246inter1));
  and2  gate2663(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2664(.a(s_302), .O(gate246inter3));
  inv1  gate2665(.a(s_303), .O(gate246inter4));
  nand2 gate2666(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2667(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2668(.a(G724), .O(gate246inter7));
  inv1  gate2669(.a(G736), .O(gate246inter8));
  nand2 gate2670(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2671(.a(s_303), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2672(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2673(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2674(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate3193(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate3194(.a(gate247inter0), .b(s_378), .O(gate247inter1));
  and2  gate3195(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate3196(.a(s_378), .O(gate247inter3));
  inv1  gate3197(.a(s_379), .O(gate247inter4));
  nand2 gate3198(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate3199(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate3200(.a(G251), .O(gate247inter7));
  inv1  gate3201(.a(G739), .O(gate247inter8));
  nand2 gate3202(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate3203(.a(s_379), .b(gate247inter3), .O(gate247inter10));
  nor2  gate3204(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate3205(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate3206(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2185(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2186(.a(gate249inter0), .b(s_234), .O(gate249inter1));
  and2  gate2187(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2188(.a(s_234), .O(gate249inter3));
  inv1  gate2189(.a(s_235), .O(gate249inter4));
  nand2 gate2190(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2191(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2192(.a(G254), .O(gate249inter7));
  inv1  gate2193(.a(G742), .O(gate249inter8));
  nand2 gate2194(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2195(.a(s_235), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2196(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2197(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2198(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2563(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2564(.a(gate252inter0), .b(s_288), .O(gate252inter1));
  and2  gate2565(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2566(.a(s_288), .O(gate252inter3));
  inv1  gate2567(.a(s_289), .O(gate252inter4));
  nand2 gate2568(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2569(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2570(.a(G709), .O(gate252inter7));
  inv1  gate2571(.a(G745), .O(gate252inter8));
  nand2 gate2572(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2573(.a(s_289), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2574(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2575(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2576(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate2367(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2368(.a(gate253inter0), .b(s_260), .O(gate253inter1));
  and2  gate2369(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2370(.a(s_260), .O(gate253inter3));
  inv1  gate2371(.a(s_261), .O(gate253inter4));
  nand2 gate2372(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2373(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2374(.a(G260), .O(gate253inter7));
  inv1  gate2375(.a(G748), .O(gate253inter8));
  nand2 gate2376(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2377(.a(s_261), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2378(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2379(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2380(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1863(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1864(.a(gate254inter0), .b(s_188), .O(gate254inter1));
  and2  gate1865(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1866(.a(s_188), .O(gate254inter3));
  inv1  gate1867(.a(s_189), .O(gate254inter4));
  nand2 gate1868(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1869(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1870(.a(G712), .O(gate254inter7));
  inv1  gate1871(.a(G748), .O(gate254inter8));
  nand2 gate1872(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1873(.a(s_189), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1874(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1875(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1876(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate729(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate730(.a(gate256inter0), .b(s_26), .O(gate256inter1));
  and2  gate731(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate732(.a(s_26), .O(gate256inter3));
  inv1  gate733(.a(s_27), .O(gate256inter4));
  nand2 gate734(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate735(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate736(.a(G715), .O(gate256inter7));
  inv1  gate737(.a(G751), .O(gate256inter8));
  nand2 gate738(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate739(.a(s_27), .b(gate256inter3), .O(gate256inter10));
  nor2  gate740(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate741(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate742(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1345(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1346(.a(gate258inter0), .b(s_114), .O(gate258inter1));
  and2  gate1347(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1348(.a(s_114), .O(gate258inter3));
  inv1  gate1349(.a(s_115), .O(gate258inter4));
  nand2 gate1350(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1351(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1352(.a(G756), .O(gate258inter7));
  inv1  gate1353(.a(G757), .O(gate258inter8));
  nand2 gate1354(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1355(.a(s_115), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1356(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1357(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1358(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate3207(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate3208(.a(gate259inter0), .b(s_380), .O(gate259inter1));
  and2  gate3209(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate3210(.a(s_380), .O(gate259inter3));
  inv1  gate3211(.a(s_381), .O(gate259inter4));
  nand2 gate3212(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate3213(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate3214(.a(G758), .O(gate259inter7));
  inv1  gate3215(.a(G759), .O(gate259inter8));
  nand2 gate3216(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate3217(.a(s_381), .b(gate259inter3), .O(gate259inter10));
  nor2  gate3218(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate3219(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate3220(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1121(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1122(.a(gate261inter0), .b(s_82), .O(gate261inter1));
  and2  gate1123(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1124(.a(s_82), .O(gate261inter3));
  inv1  gate1125(.a(s_83), .O(gate261inter4));
  nand2 gate1126(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1127(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1128(.a(G762), .O(gate261inter7));
  inv1  gate1129(.a(G763), .O(gate261inter8));
  nand2 gate1130(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1131(.a(s_83), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1132(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1133(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1134(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate3123(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate3124(.a(gate262inter0), .b(s_368), .O(gate262inter1));
  and2  gate3125(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate3126(.a(s_368), .O(gate262inter3));
  inv1  gate3127(.a(s_369), .O(gate262inter4));
  nand2 gate3128(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate3129(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate3130(.a(G764), .O(gate262inter7));
  inv1  gate3131(.a(G765), .O(gate262inter8));
  nand2 gate3132(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate3133(.a(s_369), .b(gate262inter3), .O(gate262inter10));
  nor2  gate3134(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate3135(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate3136(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2353(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2354(.a(gate263inter0), .b(s_258), .O(gate263inter1));
  and2  gate2355(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2356(.a(s_258), .O(gate263inter3));
  inv1  gate2357(.a(s_259), .O(gate263inter4));
  nand2 gate2358(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2359(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2360(.a(G766), .O(gate263inter7));
  inv1  gate2361(.a(G767), .O(gate263inter8));
  nand2 gate2362(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2363(.a(s_259), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2364(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2365(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2366(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2843(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2844(.a(gate270inter0), .b(s_328), .O(gate270inter1));
  and2  gate2845(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2846(.a(s_328), .O(gate270inter3));
  inv1  gate2847(.a(s_329), .O(gate270inter4));
  nand2 gate2848(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2849(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2850(.a(G657), .O(gate270inter7));
  inv1  gate2851(.a(G785), .O(gate270inter8));
  nand2 gate2852(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2853(.a(s_329), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2854(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2855(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2856(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate3221(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate3222(.a(gate271inter0), .b(s_382), .O(gate271inter1));
  and2  gate3223(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate3224(.a(s_382), .O(gate271inter3));
  inv1  gate3225(.a(s_383), .O(gate271inter4));
  nand2 gate3226(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate3227(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate3228(.a(G660), .O(gate271inter7));
  inv1  gate3229(.a(G788), .O(gate271inter8));
  nand2 gate3230(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate3231(.a(s_383), .b(gate271inter3), .O(gate271inter10));
  nor2  gate3232(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate3233(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate3234(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2073(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2074(.a(gate273inter0), .b(s_218), .O(gate273inter1));
  and2  gate2075(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2076(.a(s_218), .O(gate273inter3));
  inv1  gate2077(.a(s_219), .O(gate273inter4));
  nand2 gate2078(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2079(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2080(.a(G642), .O(gate273inter7));
  inv1  gate2081(.a(G794), .O(gate273inter8));
  nand2 gate2082(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2083(.a(s_219), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2084(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2085(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2086(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2479(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2480(.a(gate274inter0), .b(s_276), .O(gate274inter1));
  and2  gate2481(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2482(.a(s_276), .O(gate274inter3));
  inv1  gate2483(.a(s_277), .O(gate274inter4));
  nand2 gate2484(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2485(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2486(.a(G770), .O(gate274inter7));
  inv1  gate2487(.a(G794), .O(gate274inter8));
  nand2 gate2488(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2489(.a(s_277), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2490(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2491(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2492(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate869(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate870(.a(gate276inter0), .b(s_46), .O(gate276inter1));
  and2  gate871(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate872(.a(s_46), .O(gate276inter3));
  inv1  gate873(.a(s_47), .O(gate276inter4));
  nand2 gate874(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate875(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate876(.a(G773), .O(gate276inter7));
  inv1  gate877(.a(G797), .O(gate276inter8));
  nand2 gate878(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate879(.a(s_47), .b(gate276inter3), .O(gate276inter10));
  nor2  gate880(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate881(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate882(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate2815(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2816(.a(gate277inter0), .b(s_324), .O(gate277inter1));
  and2  gate2817(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2818(.a(s_324), .O(gate277inter3));
  inv1  gate2819(.a(s_325), .O(gate277inter4));
  nand2 gate2820(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2821(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2822(.a(G648), .O(gate277inter7));
  inv1  gate2823(.a(G800), .O(gate277inter8));
  nand2 gate2824(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2825(.a(s_325), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2826(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2827(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2828(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate2941(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2942(.a(gate278inter0), .b(s_342), .O(gate278inter1));
  and2  gate2943(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2944(.a(s_342), .O(gate278inter3));
  inv1  gate2945(.a(s_343), .O(gate278inter4));
  nand2 gate2946(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2947(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2948(.a(G776), .O(gate278inter7));
  inv1  gate2949(.a(G800), .O(gate278inter8));
  nand2 gate2950(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2951(.a(s_343), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2952(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2953(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2954(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2381(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2382(.a(gate280inter0), .b(s_262), .O(gate280inter1));
  and2  gate2383(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2384(.a(s_262), .O(gate280inter3));
  inv1  gate2385(.a(s_263), .O(gate280inter4));
  nand2 gate2386(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2387(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2388(.a(G779), .O(gate280inter7));
  inv1  gate2389(.a(G803), .O(gate280inter8));
  nand2 gate2390(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2391(.a(s_263), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2392(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2393(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2394(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate715(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate716(.a(gate282inter0), .b(s_24), .O(gate282inter1));
  and2  gate717(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate718(.a(s_24), .O(gate282inter3));
  inv1  gate719(.a(s_25), .O(gate282inter4));
  nand2 gate720(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate721(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate722(.a(G782), .O(gate282inter7));
  inv1  gate723(.a(G806), .O(gate282inter8));
  nand2 gate724(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate725(.a(s_25), .b(gate282inter3), .O(gate282inter10));
  nor2  gate726(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate727(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate728(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate3011(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate3012(.a(gate283inter0), .b(s_352), .O(gate283inter1));
  and2  gate3013(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate3014(.a(s_352), .O(gate283inter3));
  inv1  gate3015(.a(s_353), .O(gate283inter4));
  nand2 gate3016(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate3017(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate3018(.a(G657), .O(gate283inter7));
  inv1  gate3019(.a(G809), .O(gate283inter8));
  nand2 gate3020(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate3021(.a(s_353), .b(gate283inter3), .O(gate283inter10));
  nor2  gate3022(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate3023(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate3024(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1569(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1570(.a(gate287inter0), .b(s_146), .O(gate287inter1));
  and2  gate1571(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1572(.a(s_146), .O(gate287inter3));
  inv1  gate1573(.a(s_147), .O(gate287inter4));
  nand2 gate1574(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1575(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1576(.a(G663), .O(gate287inter7));
  inv1  gate1577(.a(G815), .O(gate287inter8));
  nand2 gate1578(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1579(.a(s_147), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1580(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1581(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1582(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2717(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2718(.a(gate289inter0), .b(s_310), .O(gate289inter1));
  and2  gate2719(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2720(.a(s_310), .O(gate289inter3));
  inv1  gate2721(.a(s_311), .O(gate289inter4));
  nand2 gate2722(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2723(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2724(.a(G818), .O(gate289inter7));
  inv1  gate2725(.a(G819), .O(gate289inter8));
  nand2 gate2726(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2727(.a(s_311), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2728(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2729(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2730(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate855(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate856(.a(gate291inter0), .b(s_44), .O(gate291inter1));
  and2  gate857(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate858(.a(s_44), .O(gate291inter3));
  inv1  gate859(.a(s_45), .O(gate291inter4));
  nand2 gate860(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate861(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate862(.a(G822), .O(gate291inter7));
  inv1  gate863(.a(G823), .O(gate291inter8));
  nand2 gate864(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate865(.a(s_45), .b(gate291inter3), .O(gate291inter10));
  nor2  gate866(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate867(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate868(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2045(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2046(.a(gate293inter0), .b(s_214), .O(gate293inter1));
  and2  gate2047(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2048(.a(s_214), .O(gate293inter3));
  inv1  gate2049(.a(s_215), .O(gate293inter4));
  nand2 gate2050(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2051(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2052(.a(G828), .O(gate293inter7));
  inv1  gate2053(.a(G829), .O(gate293inter8));
  nand2 gate2054(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2055(.a(s_215), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2056(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2057(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2058(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate897(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate898(.a(gate294inter0), .b(s_50), .O(gate294inter1));
  and2  gate899(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate900(.a(s_50), .O(gate294inter3));
  inv1  gate901(.a(s_51), .O(gate294inter4));
  nand2 gate902(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate903(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate904(.a(G832), .O(gate294inter7));
  inv1  gate905(.a(G833), .O(gate294inter8));
  nand2 gate906(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate907(.a(s_51), .b(gate294inter3), .O(gate294inter10));
  nor2  gate908(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate909(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate910(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1233(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1234(.a(gate295inter0), .b(s_98), .O(gate295inter1));
  and2  gate1235(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1236(.a(s_98), .O(gate295inter3));
  inv1  gate1237(.a(s_99), .O(gate295inter4));
  nand2 gate1238(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1239(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1240(.a(G830), .O(gate295inter7));
  inv1  gate1241(.a(G831), .O(gate295inter8));
  nand2 gate1242(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1243(.a(s_99), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1244(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1245(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1246(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate3053(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate3054(.a(gate296inter0), .b(s_358), .O(gate296inter1));
  and2  gate3055(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate3056(.a(s_358), .O(gate296inter3));
  inv1  gate3057(.a(s_359), .O(gate296inter4));
  nand2 gate3058(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate3059(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate3060(.a(G826), .O(gate296inter7));
  inv1  gate3061(.a(G827), .O(gate296inter8));
  nand2 gate3062(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate3063(.a(s_359), .b(gate296inter3), .O(gate296inter10));
  nor2  gate3064(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate3065(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate3066(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1219(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1220(.a(gate387inter0), .b(s_96), .O(gate387inter1));
  and2  gate1221(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1222(.a(s_96), .O(gate387inter3));
  inv1  gate1223(.a(s_97), .O(gate387inter4));
  nand2 gate1224(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1225(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1226(.a(G1), .O(gate387inter7));
  inv1  gate1227(.a(G1036), .O(gate387inter8));
  nand2 gate1228(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1229(.a(s_97), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1230(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1231(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1232(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1457(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1458(.a(gate388inter0), .b(s_130), .O(gate388inter1));
  and2  gate1459(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1460(.a(s_130), .O(gate388inter3));
  inv1  gate1461(.a(s_131), .O(gate388inter4));
  nand2 gate1462(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1463(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1464(.a(G2), .O(gate388inter7));
  inv1  gate1465(.a(G1039), .O(gate388inter8));
  nand2 gate1466(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1467(.a(s_131), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1468(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1469(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1470(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1821(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1822(.a(gate390inter0), .b(s_182), .O(gate390inter1));
  and2  gate1823(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1824(.a(s_182), .O(gate390inter3));
  inv1  gate1825(.a(s_183), .O(gate390inter4));
  nand2 gate1826(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1827(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1828(.a(G4), .O(gate390inter7));
  inv1  gate1829(.a(G1045), .O(gate390inter8));
  nand2 gate1830(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1831(.a(s_183), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1832(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1833(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1834(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1177(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1178(.a(gate391inter0), .b(s_90), .O(gate391inter1));
  and2  gate1179(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1180(.a(s_90), .O(gate391inter3));
  inv1  gate1181(.a(s_91), .O(gate391inter4));
  nand2 gate1182(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1183(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1184(.a(G5), .O(gate391inter7));
  inv1  gate1185(.a(G1048), .O(gate391inter8));
  nand2 gate1186(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1187(.a(s_91), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1188(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1189(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1190(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate911(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate912(.a(gate394inter0), .b(s_52), .O(gate394inter1));
  and2  gate913(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate914(.a(s_52), .O(gate394inter3));
  inv1  gate915(.a(s_53), .O(gate394inter4));
  nand2 gate916(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate917(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate918(.a(G8), .O(gate394inter7));
  inv1  gate919(.a(G1057), .O(gate394inter8));
  nand2 gate920(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate921(.a(s_53), .b(gate394inter3), .O(gate394inter10));
  nor2  gate922(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate923(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate924(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate2759(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2760(.a(gate395inter0), .b(s_316), .O(gate395inter1));
  and2  gate2761(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2762(.a(s_316), .O(gate395inter3));
  inv1  gate2763(.a(s_317), .O(gate395inter4));
  nand2 gate2764(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2765(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2766(.a(G9), .O(gate395inter7));
  inv1  gate2767(.a(G1060), .O(gate395inter8));
  nand2 gate2768(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2769(.a(s_317), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2770(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2771(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2772(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1093(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1094(.a(gate396inter0), .b(s_78), .O(gate396inter1));
  and2  gate1095(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1096(.a(s_78), .O(gate396inter3));
  inv1  gate1097(.a(s_79), .O(gate396inter4));
  nand2 gate1098(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1099(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1100(.a(G10), .O(gate396inter7));
  inv1  gate1101(.a(G1063), .O(gate396inter8));
  nand2 gate1102(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1103(.a(s_79), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1104(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1105(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1106(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate3165(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate3166(.a(gate398inter0), .b(s_374), .O(gate398inter1));
  and2  gate3167(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate3168(.a(s_374), .O(gate398inter3));
  inv1  gate3169(.a(s_375), .O(gate398inter4));
  nand2 gate3170(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate3171(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate3172(.a(G12), .O(gate398inter7));
  inv1  gate3173(.a(G1069), .O(gate398inter8));
  nand2 gate3174(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate3175(.a(s_375), .b(gate398inter3), .O(gate398inter10));
  nor2  gate3176(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate3177(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate3178(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1891(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1892(.a(gate400inter0), .b(s_192), .O(gate400inter1));
  and2  gate1893(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1894(.a(s_192), .O(gate400inter3));
  inv1  gate1895(.a(s_193), .O(gate400inter4));
  nand2 gate1896(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1897(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1898(.a(G14), .O(gate400inter7));
  inv1  gate1899(.a(G1075), .O(gate400inter8));
  nand2 gate1900(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1901(.a(s_193), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1902(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1903(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1904(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1373(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1374(.a(gate402inter0), .b(s_118), .O(gate402inter1));
  and2  gate1375(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1376(.a(s_118), .O(gate402inter3));
  inv1  gate1377(.a(s_119), .O(gate402inter4));
  nand2 gate1378(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1379(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1380(.a(G16), .O(gate402inter7));
  inv1  gate1381(.a(G1081), .O(gate402inter8));
  nand2 gate1382(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1383(.a(s_119), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1384(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1385(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1386(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate2157(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2158(.a(gate405inter0), .b(s_230), .O(gate405inter1));
  and2  gate2159(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2160(.a(s_230), .O(gate405inter3));
  inv1  gate2161(.a(s_231), .O(gate405inter4));
  nand2 gate2162(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2163(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2164(.a(G19), .O(gate405inter7));
  inv1  gate2165(.a(G1090), .O(gate405inter8));
  nand2 gate2166(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2167(.a(s_231), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2168(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2169(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2170(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate673(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate674(.a(gate408inter0), .b(s_18), .O(gate408inter1));
  and2  gate675(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate676(.a(s_18), .O(gate408inter3));
  inv1  gate677(.a(s_19), .O(gate408inter4));
  nand2 gate678(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate679(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate680(.a(G22), .O(gate408inter7));
  inv1  gate681(.a(G1099), .O(gate408inter8));
  nand2 gate682(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate683(.a(s_19), .b(gate408inter3), .O(gate408inter10));
  nor2  gate684(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate685(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate686(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1723(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1724(.a(gate409inter0), .b(s_168), .O(gate409inter1));
  and2  gate1725(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1726(.a(s_168), .O(gate409inter3));
  inv1  gate1727(.a(s_169), .O(gate409inter4));
  nand2 gate1728(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1729(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1730(.a(G23), .O(gate409inter7));
  inv1  gate1731(.a(G1102), .O(gate409inter8));
  nand2 gate1732(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1733(.a(s_169), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1734(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1735(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1736(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate757(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate758(.a(gate410inter0), .b(s_30), .O(gate410inter1));
  and2  gate759(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate760(.a(s_30), .O(gate410inter3));
  inv1  gate761(.a(s_31), .O(gate410inter4));
  nand2 gate762(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate763(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate764(.a(G24), .O(gate410inter7));
  inv1  gate765(.a(G1105), .O(gate410inter8));
  nand2 gate766(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate767(.a(s_31), .b(gate410inter3), .O(gate410inter10));
  nor2  gate768(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate769(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate770(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1079(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1080(.a(gate412inter0), .b(s_76), .O(gate412inter1));
  and2  gate1081(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1082(.a(s_76), .O(gate412inter3));
  inv1  gate1083(.a(s_77), .O(gate412inter4));
  nand2 gate1084(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1085(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1086(.a(G26), .O(gate412inter7));
  inv1  gate1087(.a(G1111), .O(gate412inter8));
  nand2 gate1088(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1089(.a(s_77), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1090(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1091(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1092(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate953(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate954(.a(gate413inter0), .b(s_58), .O(gate413inter1));
  and2  gate955(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate956(.a(s_58), .O(gate413inter3));
  inv1  gate957(.a(s_59), .O(gate413inter4));
  nand2 gate958(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate959(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate960(.a(G27), .O(gate413inter7));
  inv1  gate961(.a(G1114), .O(gate413inter8));
  nand2 gate962(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate963(.a(s_59), .b(gate413inter3), .O(gate413inter10));
  nor2  gate964(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate965(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate966(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2297(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2298(.a(gate414inter0), .b(s_250), .O(gate414inter1));
  and2  gate2299(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2300(.a(s_250), .O(gate414inter3));
  inv1  gate2301(.a(s_251), .O(gate414inter4));
  nand2 gate2302(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2303(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2304(.a(G28), .O(gate414inter7));
  inv1  gate2305(.a(G1117), .O(gate414inter8));
  nand2 gate2306(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2307(.a(s_251), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2308(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2309(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2310(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate701(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate702(.a(gate415inter0), .b(s_22), .O(gate415inter1));
  and2  gate703(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate704(.a(s_22), .O(gate415inter3));
  inv1  gate705(.a(s_23), .O(gate415inter4));
  nand2 gate706(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate707(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate708(.a(G29), .O(gate415inter7));
  inv1  gate709(.a(G1120), .O(gate415inter8));
  nand2 gate710(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate711(.a(s_23), .b(gate415inter3), .O(gate415inter10));
  nor2  gate712(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate713(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate714(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1611(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1612(.a(gate417inter0), .b(s_152), .O(gate417inter1));
  and2  gate1613(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1614(.a(s_152), .O(gate417inter3));
  inv1  gate1615(.a(s_153), .O(gate417inter4));
  nand2 gate1616(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1617(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1618(.a(G31), .O(gate417inter7));
  inv1  gate1619(.a(G1126), .O(gate417inter8));
  nand2 gate1620(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1621(.a(s_153), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1622(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1623(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1624(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1471(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1472(.a(gate419inter0), .b(s_132), .O(gate419inter1));
  and2  gate1473(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1474(.a(s_132), .O(gate419inter3));
  inv1  gate1475(.a(s_133), .O(gate419inter4));
  nand2 gate1476(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1477(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1478(.a(G1), .O(gate419inter7));
  inv1  gate1479(.a(G1132), .O(gate419inter8));
  nand2 gate1480(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1481(.a(s_133), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1482(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1483(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1484(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2885(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2886(.a(gate420inter0), .b(s_334), .O(gate420inter1));
  and2  gate2887(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2888(.a(s_334), .O(gate420inter3));
  inv1  gate2889(.a(s_335), .O(gate420inter4));
  nand2 gate2890(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2891(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2892(.a(G1036), .O(gate420inter7));
  inv1  gate2893(.a(G1132), .O(gate420inter8));
  nand2 gate2894(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2895(.a(s_335), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2896(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2897(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2898(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate827(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate828(.a(gate423inter0), .b(s_40), .O(gate423inter1));
  and2  gate829(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate830(.a(s_40), .O(gate423inter3));
  inv1  gate831(.a(s_41), .O(gate423inter4));
  nand2 gate832(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate833(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate834(.a(G3), .O(gate423inter7));
  inv1  gate835(.a(G1138), .O(gate423inter8));
  nand2 gate836(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate837(.a(s_41), .b(gate423inter3), .O(gate423inter10));
  nor2  gate838(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate839(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate840(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2605(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2606(.a(gate424inter0), .b(s_294), .O(gate424inter1));
  and2  gate2607(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2608(.a(s_294), .O(gate424inter3));
  inv1  gate2609(.a(s_295), .O(gate424inter4));
  nand2 gate2610(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2611(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2612(.a(G1042), .O(gate424inter7));
  inv1  gate2613(.a(G1138), .O(gate424inter8));
  nand2 gate2614(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2615(.a(s_295), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2616(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2617(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2618(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2115(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2116(.a(gate427inter0), .b(s_224), .O(gate427inter1));
  and2  gate2117(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2118(.a(s_224), .O(gate427inter3));
  inv1  gate2119(.a(s_225), .O(gate427inter4));
  nand2 gate2120(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2121(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2122(.a(G5), .O(gate427inter7));
  inv1  gate2123(.a(G1144), .O(gate427inter8));
  nand2 gate2124(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2125(.a(s_225), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2126(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2127(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2128(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate743(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate744(.a(gate428inter0), .b(s_28), .O(gate428inter1));
  and2  gate745(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate746(.a(s_28), .O(gate428inter3));
  inv1  gate747(.a(s_29), .O(gate428inter4));
  nand2 gate748(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate749(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate750(.a(G1048), .O(gate428inter7));
  inv1  gate751(.a(G1144), .O(gate428inter8));
  nand2 gate752(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate753(.a(s_29), .b(gate428inter3), .O(gate428inter10));
  nor2  gate754(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate755(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate756(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate2899(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2900(.a(gate429inter0), .b(s_336), .O(gate429inter1));
  and2  gate2901(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2902(.a(s_336), .O(gate429inter3));
  inv1  gate2903(.a(s_337), .O(gate429inter4));
  nand2 gate2904(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2905(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2906(.a(G6), .O(gate429inter7));
  inv1  gate2907(.a(G1147), .O(gate429inter8));
  nand2 gate2908(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2909(.a(s_337), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2910(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2911(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2912(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate3081(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate3082(.a(gate431inter0), .b(s_362), .O(gate431inter1));
  and2  gate3083(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate3084(.a(s_362), .O(gate431inter3));
  inv1  gate3085(.a(s_363), .O(gate431inter4));
  nand2 gate3086(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate3087(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate3088(.a(G7), .O(gate431inter7));
  inv1  gate3089(.a(G1150), .O(gate431inter8));
  nand2 gate3090(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate3091(.a(s_363), .b(gate431inter3), .O(gate431inter10));
  nor2  gate3092(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate3093(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate3094(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1583(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1584(.a(gate432inter0), .b(s_148), .O(gate432inter1));
  and2  gate1585(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1586(.a(s_148), .O(gate432inter3));
  inv1  gate1587(.a(s_149), .O(gate432inter4));
  nand2 gate1588(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1589(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1590(.a(G1054), .O(gate432inter7));
  inv1  gate1591(.a(G1150), .O(gate432inter8));
  nand2 gate1592(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1593(.a(s_149), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1594(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1595(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1596(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2969(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2970(.a(gate435inter0), .b(s_346), .O(gate435inter1));
  and2  gate2971(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2972(.a(s_346), .O(gate435inter3));
  inv1  gate2973(.a(s_347), .O(gate435inter4));
  nand2 gate2974(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2975(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2976(.a(G9), .O(gate435inter7));
  inv1  gate2977(.a(G1156), .O(gate435inter8));
  nand2 gate2978(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2979(.a(s_347), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2980(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2981(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2982(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1681(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1682(.a(gate446inter0), .b(s_162), .O(gate446inter1));
  and2  gate1683(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1684(.a(s_162), .O(gate446inter3));
  inv1  gate1685(.a(s_163), .O(gate446inter4));
  nand2 gate1686(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1687(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1688(.a(G1075), .O(gate446inter7));
  inv1  gate1689(.a(G1171), .O(gate446inter8));
  nand2 gate1690(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1691(.a(s_163), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1692(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1693(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1694(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2927(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2928(.a(gate447inter0), .b(s_340), .O(gate447inter1));
  and2  gate2929(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2930(.a(s_340), .O(gate447inter3));
  inv1  gate2931(.a(s_341), .O(gate447inter4));
  nand2 gate2932(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2933(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2934(.a(G15), .O(gate447inter7));
  inv1  gate2935(.a(G1174), .O(gate447inter8));
  nand2 gate2936(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2937(.a(s_341), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2938(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2939(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2940(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate771(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate772(.a(gate448inter0), .b(s_32), .O(gate448inter1));
  and2  gate773(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate774(.a(s_32), .O(gate448inter3));
  inv1  gate775(.a(s_33), .O(gate448inter4));
  nand2 gate776(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate777(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate778(.a(G1078), .O(gate448inter7));
  inv1  gate779(.a(G1174), .O(gate448inter8));
  nand2 gate780(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate781(.a(s_33), .b(gate448inter3), .O(gate448inter10));
  nor2  gate782(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate783(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate784(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2465(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2466(.a(gate449inter0), .b(s_274), .O(gate449inter1));
  and2  gate2467(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2468(.a(s_274), .O(gate449inter3));
  inv1  gate2469(.a(s_275), .O(gate449inter4));
  nand2 gate2470(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2471(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2472(.a(G16), .O(gate449inter7));
  inv1  gate2473(.a(G1177), .O(gate449inter8));
  nand2 gate2474(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2475(.a(s_275), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2476(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2477(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2478(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate813(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate814(.a(gate456inter0), .b(s_38), .O(gate456inter1));
  and2  gate815(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate816(.a(s_38), .O(gate456inter3));
  inv1  gate817(.a(s_39), .O(gate456inter4));
  nand2 gate818(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate819(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate820(.a(G1090), .O(gate456inter7));
  inv1  gate821(.a(G1186), .O(gate456inter8));
  nand2 gate822(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate823(.a(s_39), .b(gate456inter3), .O(gate456inter10));
  nor2  gate824(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate825(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate826(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate2647(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2648(.a(gate457inter0), .b(s_300), .O(gate457inter1));
  and2  gate2649(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2650(.a(s_300), .O(gate457inter3));
  inv1  gate2651(.a(s_301), .O(gate457inter4));
  nand2 gate2652(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2653(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2654(.a(G20), .O(gate457inter7));
  inv1  gate2655(.a(G1189), .O(gate457inter8));
  nand2 gate2656(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2657(.a(s_301), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2658(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2659(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2660(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1009(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1010(.a(gate458inter0), .b(s_66), .O(gate458inter1));
  and2  gate1011(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1012(.a(s_66), .O(gate458inter3));
  inv1  gate1013(.a(s_67), .O(gate458inter4));
  nand2 gate1014(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1015(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1016(.a(G1093), .O(gate458inter7));
  inv1  gate1017(.a(G1189), .O(gate458inter8));
  nand2 gate1018(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1019(.a(s_67), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1020(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1021(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1022(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1849(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1850(.a(gate460inter0), .b(s_186), .O(gate460inter1));
  and2  gate1851(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1852(.a(s_186), .O(gate460inter3));
  inv1  gate1853(.a(s_187), .O(gate460inter4));
  nand2 gate1854(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1855(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1856(.a(G1096), .O(gate460inter7));
  inv1  gate1857(.a(G1192), .O(gate460inter8));
  nand2 gate1858(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1859(.a(s_187), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1860(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1861(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1862(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1191(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1192(.a(gate463inter0), .b(s_92), .O(gate463inter1));
  and2  gate1193(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1194(.a(s_92), .O(gate463inter3));
  inv1  gate1195(.a(s_93), .O(gate463inter4));
  nand2 gate1196(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1197(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1198(.a(G23), .O(gate463inter7));
  inv1  gate1199(.a(G1198), .O(gate463inter8));
  nand2 gate1200(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1201(.a(s_93), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1202(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1203(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1204(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate2199(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2200(.a(gate464inter0), .b(s_236), .O(gate464inter1));
  and2  gate2201(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2202(.a(s_236), .O(gate464inter3));
  inv1  gate2203(.a(s_237), .O(gate464inter4));
  nand2 gate2204(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2205(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2206(.a(G1102), .O(gate464inter7));
  inv1  gate2207(.a(G1198), .O(gate464inter8));
  nand2 gate2208(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2209(.a(s_237), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2210(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2211(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2212(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1905(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1906(.a(gate467inter0), .b(s_194), .O(gate467inter1));
  and2  gate1907(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1908(.a(s_194), .O(gate467inter3));
  inv1  gate1909(.a(s_195), .O(gate467inter4));
  nand2 gate1910(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1911(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1912(.a(G25), .O(gate467inter7));
  inv1  gate1913(.a(G1204), .O(gate467inter8));
  nand2 gate1914(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1915(.a(s_195), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1916(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1917(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1918(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2213(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2214(.a(gate469inter0), .b(s_238), .O(gate469inter1));
  and2  gate2215(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2216(.a(s_238), .O(gate469inter3));
  inv1  gate2217(.a(s_239), .O(gate469inter4));
  nand2 gate2218(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2219(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2220(.a(G26), .O(gate469inter7));
  inv1  gate2221(.a(G1207), .O(gate469inter8));
  nand2 gate2222(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2223(.a(s_239), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2224(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2225(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2226(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate2829(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2830(.a(gate470inter0), .b(s_326), .O(gate470inter1));
  and2  gate2831(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2832(.a(s_326), .O(gate470inter3));
  inv1  gate2833(.a(s_327), .O(gate470inter4));
  nand2 gate2834(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2835(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2836(.a(G1111), .O(gate470inter7));
  inv1  gate2837(.a(G1207), .O(gate470inter8));
  nand2 gate2838(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2839(.a(s_327), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2840(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2841(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2842(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1205(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1206(.a(gate471inter0), .b(s_94), .O(gate471inter1));
  and2  gate1207(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1208(.a(s_94), .O(gate471inter3));
  inv1  gate1209(.a(s_95), .O(gate471inter4));
  nand2 gate1210(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1211(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1212(.a(G27), .O(gate471inter7));
  inv1  gate1213(.a(G1210), .O(gate471inter8));
  nand2 gate1214(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1215(.a(s_95), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1216(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1217(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1218(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1835(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1836(.a(gate476inter0), .b(s_184), .O(gate476inter1));
  and2  gate1837(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1838(.a(s_184), .O(gate476inter3));
  inv1  gate1839(.a(s_185), .O(gate476inter4));
  nand2 gate1840(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1841(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1842(.a(G1120), .O(gate476inter7));
  inv1  gate1843(.a(G1216), .O(gate476inter8));
  nand2 gate1844(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1845(.a(s_185), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1846(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1847(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1848(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1303(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1304(.a(gate480inter0), .b(s_108), .O(gate480inter1));
  and2  gate1305(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1306(.a(s_108), .O(gate480inter3));
  inv1  gate1307(.a(s_109), .O(gate480inter4));
  nand2 gate1308(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1309(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1310(.a(G1126), .O(gate480inter7));
  inv1  gate1311(.a(G1222), .O(gate480inter8));
  nand2 gate1312(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1313(.a(s_109), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1314(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1315(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1316(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2423(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2424(.a(gate482inter0), .b(s_268), .O(gate482inter1));
  and2  gate2425(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2426(.a(s_268), .O(gate482inter3));
  inv1  gate2427(.a(s_269), .O(gate482inter4));
  nand2 gate2428(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2429(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2430(.a(G1129), .O(gate482inter7));
  inv1  gate2431(.a(G1225), .O(gate482inter8));
  nand2 gate2432(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2433(.a(s_269), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2434(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2435(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2436(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1359(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1360(.a(gate487inter0), .b(s_116), .O(gate487inter1));
  and2  gate1361(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1362(.a(s_116), .O(gate487inter3));
  inv1  gate1363(.a(s_117), .O(gate487inter4));
  nand2 gate1364(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1365(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1366(.a(G1236), .O(gate487inter7));
  inv1  gate1367(.a(G1237), .O(gate487inter8));
  nand2 gate1368(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1369(.a(s_117), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1370(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1371(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1372(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1667(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1668(.a(gate490inter0), .b(s_160), .O(gate490inter1));
  and2  gate1669(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1670(.a(s_160), .O(gate490inter3));
  inv1  gate1671(.a(s_161), .O(gate490inter4));
  nand2 gate1672(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1673(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1674(.a(G1242), .O(gate490inter7));
  inv1  gate1675(.a(G1243), .O(gate490inter8));
  nand2 gate1676(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1677(.a(s_161), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1678(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1679(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1680(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1163(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1164(.a(gate501inter0), .b(s_88), .O(gate501inter1));
  and2  gate1165(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1166(.a(s_88), .O(gate501inter3));
  inv1  gate1167(.a(s_89), .O(gate501inter4));
  nand2 gate1168(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1169(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1170(.a(G1264), .O(gate501inter7));
  inv1  gate1171(.a(G1265), .O(gate501inter8));
  nand2 gate1172(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1173(.a(s_89), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1174(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1175(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1176(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1275(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1276(.a(gate502inter0), .b(s_104), .O(gate502inter1));
  and2  gate1277(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1278(.a(s_104), .O(gate502inter3));
  inv1  gate1279(.a(s_105), .O(gate502inter4));
  nand2 gate1280(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1281(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1282(.a(G1266), .O(gate502inter7));
  inv1  gate1283(.a(G1267), .O(gate502inter8));
  nand2 gate1284(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1285(.a(s_105), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1286(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1287(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1288(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1919(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1920(.a(gate504inter0), .b(s_196), .O(gate504inter1));
  and2  gate1921(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1922(.a(s_196), .O(gate504inter3));
  inv1  gate1923(.a(s_197), .O(gate504inter4));
  nand2 gate1924(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1925(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1926(.a(G1270), .O(gate504inter7));
  inv1  gate1927(.a(G1271), .O(gate504inter8));
  nand2 gate1928(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1929(.a(s_197), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1930(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1931(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1932(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2493(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2494(.a(gate508inter0), .b(s_278), .O(gate508inter1));
  and2  gate2495(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2496(.a(s_278), .O(gate508inter3));
  inv1  gate2497(.a(s_279), .O(gate508inter4));
  nand2 gate2498(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2499(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2500(.a(G1278), .O(gate508inter7));
  inv1  gate2501(.a(G1279), .O(gate508inter8));
  nand2 gate2502(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2503(.a(s_279), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2504(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2505(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2506(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2171(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2172(.a(gate509inter0), .b(s_232), .O(gate509inter1));
  and2  gate2173(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2174(.a(s_232), .O(gate509inter3));
  inv1  gate2175(.a(s_233), .O(gate509inter4));
  nand2 gate2176(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2177(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2178(.a(G1280), .O(gate509inter7));
  inv1  gate2179(.a(G1281), .O(gate509inter8));
  nand2 gate2180(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2181(.a(s_233), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2182(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2183(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2184(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate2997(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2998(.a(gate510inter0), .b(s_350), .O(gate510inter1));
  and2  gate2999(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate3000(.a(s_350), .O(gate510inter3));
  inv1  gate3001(.a(s_351), .O(gate510inter4));
  nand2 gate3002(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate3003(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate3004(.a(G1282), .O(gate510inter7));
  inv1  gate3005(.a(G1283), .O(gate510inter8));
  nand2 gate3006(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate3007(.a(s_351), .b(gate510inter3), .O(gate510inter10));
  nor2  gate3008(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate3009(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate3010(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1639(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1640(.a(gate511inter0), .b(s_156), .O(gate511inter1));
  and2  gate1641(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1642(.a(s_156), .O(gate511inter3));
  inv1  gate1643(.a(s_157), .O(gate511inter4));
  nand2 gate1644(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1645(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1646(.a(G1284), .O(gate511inter7));
  inv1  gate1647(.a(G1285), .O(gate511inter8));
  nand2 gate1648(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1649(.a(s_157), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1650(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1651(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1652(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2437(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2438(.a(gate513inter0), .b(s_270), .O(gate513inter1));
  and2  gate2439(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2440(.a(s_270), .O(gate513inter3));
  inv1  gate2441(.a(s_271), .O(gate513inter4));
  nand2 gate2442(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2443(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2444(.a(G1288), .O(gate513inter7));
  inv1  gate2445(.a(G1289), .O(gate513inter8));
  nand2 gate2446(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2447(.a(s_271), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2448(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2449(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2450(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule