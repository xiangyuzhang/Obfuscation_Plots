module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1275(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1276(.a(gate17inter0), .b(s_104), .O(gate17inter1));
  and2  gate1277(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1278(.a(s_104), .O(gate17inter3));
  inv1  gate1279(.a(s_105), .O(gate17inter4));
  nand2 gate1280(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1281(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1282(.a(G17), .O(gate17inter7));
  inv1  gate1283(.a(G18), .O(gate17inter8));
  nand2 gate1284(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1285(.a(s_105), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1286(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1287(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1288(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate575(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate576(.a(gate40inter0), .b(s_4), .O(gate40inter1));
  and2  gate577(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate578(.a(s_4), .O(gate40inter3));
  inv1  gate579(.a(s_5), .O(gate40inter4));
  nand2 gate580(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate581(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate582(.a(G28), .O(gate40inter7));
  inv1  gate583(.a(G32), .O(gate40inter8));
  nand2 gate584(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate585(.a(s_5), .b(gate40inter3), .O(gate40inter10));
  nor2  gate586(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate587(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate588(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1233(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1234(.a(gate46inter0), .b(s_98), .O(gate46inter1));
  and2  gate1235(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1236(.a(s_98), .O(gate46inter3));
  inv1  gate1237(.a(s_99), .O(gate46inter4));
  nand2 gate1238(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1239(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1240(.a(G6), .O(gate46inter7));
  inv1  gate1241(.a(G272), .O(gate46inter8));
  nand2 gate1242(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1243(.a(s_99), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1244(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1245(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1246(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate743(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate744(.a(gate47inter0), .b(s_28), .O(gate47inter1));
  and2  gate745(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate746(.a(s_28), .O(gate47inter3));
  inv1  gate747(.a(s_29), .O(gate47inter4));
  nand2 gate748(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate749(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate750(.a(G7), .O(gate47inter7));
  inv1  gate751(.a(G275), .O(gate47inter8));
  nand2 gate752(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate753(.a(s_29), .b(gate47inter3), .O(gate47inter10));
  nor2  gate754(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate755(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate756(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate547(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate548(.a(gate58inter0), .b(s_0), .O(gate58inter1));
  and2  gate549(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate550(.a(s_0), .O(gate58inter3));
  inv1  gate551(.a(s_1), .O(gate58inter4));
  nand2 gate552(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate553(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate554(.a(G18), .O(gate58inter7));
  inv1  gate555(.a(G290), .O(gate58inter8));
  nand2 gate556(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate557(.a(s_1), .b(gate58inter3), .O(gate58inter10));
  nor2  gate558(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate559(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate560(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1051(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1052(.a(gate59inter0), .b(s_72), .O(gate59inter1));
  and2  gate1053(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1054(.a(s_72), .O(gate59inter3));
  inv1  gate1055(.a(s_73), .O(gate59inter4));
  nand2 gate1056(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1057(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1058(.a(G19), .O(gate59inter7));
  inv1  gate1059(.a(G293), .O(gate59inter8));
  nand2 gate1060(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1061(.a(s_73), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1062(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1063(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1064(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate687(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate688(.a(gate61inter0), .b(s_20), .O(gate61inter1));
  and2  gate689(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate690(.a(s_20), .O(gate61inter3));
  inv1  gate691(.a(s_21), .O(gate61inter4));
  nand2 gate692(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate693(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate694(.a(G21), .O(gate61inter7));
  inv1  gate695(.a(G296), .O(gate61inter8));
  nand2 gate696(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate697(.a(s_21), .b(gate61inter3), .O(gate61inter10));
  nor2  gate698(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate699(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate700(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate701(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate702(.a(gate64inter0), .b(s_22), .O(gate64inter1));
  and2  gate703(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate704(.a(s_22), .O(gate64inter3));
  inv1  gate705(.a(s_23), .O(gate64inter4));
  nand2 gate706(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate707(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate708(.a(G24), .O(gate64inter7));
  inv1  gate709(.a(G299), .O(gate64inter8));
  nand2 gate710(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate711(.a(s_23), .b(gate64inter3), .O(gate64inter10));
  nor2  gate712(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate713(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate714(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1163(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1164(.a(gate66inter0), .b(s_88), .O(gate66inter1));
  and2  gate1165(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1166(.a(s_88), .O(gate66inter3));
  inv1  gate1167(.a(s_89), .O(gate66inter4));
  nand2 gate1168(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1169(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1170(.a(G26), .O(gate66inter7));
  inv1  gate1171(.a(G302), .O(gate66inter8));
  nand2 gate1172(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1173(.a(s_89), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1174(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1175(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1176(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate729(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate730(.a(gate70inter0), .b(s_26), .O(gate70inter1));
  and2  gate731(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate732(.a(s_26), .O(gate70inter3));
  inv1  gate733(.a(s_27), .O(gate70inter4));
  nand2 gate734(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate735(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate736(.a(G30), .O(gate70inter7));
  inv1  gate737(.a(G308), .O(gate70inter8));
  nand2 gate738(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate739(.a(s_27), .b(gate70inter3), .O(gate70inter10));
  nor2  gate740(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate741(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate742(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1121(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1122(.a(gate73inter0), .b(s_82), .O(gate73inter1));
  and2  gate1123(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1124(.a(s_82), .O(gate73inter3));
  inv1  gate1125(.a(s_83), .O(gate73inter4));
  nand2 gate1126(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1127(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1128(.a(G1), .O(gate73inter7));
  inv1  gate1129(.a(G314), .O(gate73inter8));
  nand2 gate1130(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1131(.a(s_83), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1132(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1133(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1134(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1009(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1010(.a(gate81inter0), .b(s_66), .O(gate81inter1));
  and2  gate1011(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1012(.a(s_66), .O(gate81inter3));
  inv1  gate1013(.a(s_67), .O(gate81inter4));
  nand2 gate1014(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1015(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1016(.a(G3), .O(gate81inter7));
  inv1  gate1017(.a(G326), .O(gate81inter8));
  nand2 gate1018(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1019(.a(s_67), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1020(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1021(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1022(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1261(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1262(.a(gate83inter0), .b(s_102), .O(gate83inter1));
  and2  gate1263(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1264(.a(s_102), .O(gate83inter3));
  inv1  gate1265(.a(s_103), .O(gate83inter4));
  nand2 gate1266(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1267(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1268(.a(G11), .O(gate83inter7));
  inv1  gate1269(.a(G329), .O(gate83inter8));
  nand2 gate1270(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1271(.a(s_103), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1272(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1273(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1274(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate659(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate660(.a(gate95inter0), .b(s_16), .O(gate95inter1));
  and2  gate661(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate662(.a(s_16), .O(gate95inter3));
  inv1  gate663(.a(s_17), .O(gate95inter4));
  nand2 gate664(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate665(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate666(.a(G26), .O(gate95inter7));
  inv1  gate667(.a(G347), .O(gate95inter8));
  nand2 gate668(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate669(.a(s_17), .b(gate95inter3), .O(gate95inter10));
  nor2  gate670(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate671(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate672(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate953(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate954(.a(gate99inter0), .b(s_58), .O(gate99inter1));
  and2  gate955(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate956(.a(s_58), .O(gate99inter3));
  inv1  gate957(.a(s_59), .O(gate99inter4));
  nand2 gate958(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate959(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate960(.a(G27), .O(gate99inter7));
  inv1  gate961(.a(G353), .O(gate99inter8));
  nand2 gate962(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate963(.a(s_59), .b(gate99inter3), .O(gate99inter10));
  nor2  gate964(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate965(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate966(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1135(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1136(.a(gate104inter0), .b(s_84), .O(gate104inter1));
  and2  gate1137(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1138(.a(s_84), .O(gate104inter3));
  inv1  gate1139(.a(s_85), .O(gate104inter4));
  nand2 gate1140(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1141(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1142(.a(G32), .O(gate104inter7));
  inv1  gate1143(.a(G359), .O(gate104inter8));
  nand2 gate1144(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1145(.a(s_85), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1146(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1147(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1148(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1079(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1080(.a(gate112inter0), .b(s_76), .O(gate112inter1));
  and2  gate1081(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1082(.a(s_76), .O(gate112inter3));
  inv1  gate1083(.a(s_77), .O(gate112inter4));
  nand2 gate1084(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1085(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1086(.a(G376), .O(gate112inter7));
  inv1  gate1087(.a(G377), .O(gate112inter8));
  nand2 gate1088(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1089(.a(s_77), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1090(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1091(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1092(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate911(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate912(.a(gate119inter0), .b(s_52), .O(gate119inter1));
  and2  gate913(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate914(.a(s_52), .O(gate119inter3));
  inv1  gate915(.a(s_53), .O(gate119inter4));
  nand2 gate916(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate917(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate918(.a(G390), .O(gate119inter7));
  inv1  gate919(.a(G391), .O(gate119inter8));
  nand2 gate920(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate921(.a(s_53), .b(gate119inter3), .O(gate119inter10));
  nor2  gate922(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate923(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate924(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1149(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1150(.a(gate126inter0), .b(s_86), .O(gate126inter1));
  and2  gate1151(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1152(.a(s_86), .O(gate126inter3));
  inv1  gate1153(.a(s_87), .O(gate126inter4));
  nand2 gate1154(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1155(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1156(.a(G404), .O(gate126inter7));
  inv1  gate1157(.a(G405), .O(gate126inter8));
  nand2 gate1158(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1159(.a(s_87), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1160(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1161(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1162(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1107(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1108(.a(gate142inter0), .b(s_80), .O(gate142inter1));
  and2  gate1109(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1110(.a(s_80), .O(gate142inter3));
  inv1  gate1111(.a(s_81), .O(gate142inter4));
  nand2 gate1112(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1113(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1114(.a(G456), .O(gate142inter7));
  inv1  gate1115(.a(G459), .O(gate142inter8));
  nand2 gate1116(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1117(.a(s_81), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1118(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1119(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1120(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1065(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1066(.a(gate161inter0), .b(s_74), .O(gate161inter1));
  and2  gate1067(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1068(.a(s_74), .O(gate161inter3));
  inv1  gate1069(.a(s_75), .O(gate161inter4));
  nand2 gate1070(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1071(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1072(.a(G450), .O(gate161inter7));
  inv1  gate1073(.a(G534), .O(gate161inter8));
  nand2 gate1074(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1075(.a(s_75), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1076(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1077(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1078(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate561(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate562(.a(gate164inter0), .b(s_2), .O(gate164inter1));
  and2  gate563(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate564(.a(s_2), .O(gate164inter3));
  inv1  gate565(.a(s_3), .O(gate164inter4));
  nand2 gate566(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate567(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate568(.a(G459), .O(gate164inter7));
  inv1  gate569(.a(G537), .O(gate164inter8));
  nand2 gate570(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate571(.a(s_3), .b(gate164inter3), .O(gate164inter10));
  nor2  gate572(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate573(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate574(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1191(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1192(.a(gate170inter0), .b(s_92), .O(gate170inter1));
  and2  gate1193(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1194(.a(s_92), .O(gate170inter3));
  inv1  gate1195(.a(s_93), .O(gate170inter4));
  nand2 gate1196(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1197(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1198(.a(G477), .O(gate170inter7));
  inv1  gate1199(.a(G546), .O(gate170inter8));
  nand2 gate1200(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1201(.a(s_93), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1202(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1203(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1204(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate673(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate674(.a(gate176inter0), .b(s_18), .O(gate176inter1));
  and2  gate675(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate676(.a(s_18), .O(gate176inter3));
  inv1  gate677(.a(s_19), .O(gate176inter4));
  nand2 gate678(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate679(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate680(.a(G495), .O(gate176inter7));
  inv1  gate681(.a(G555), .O(gate176inter8));
  nand2 gate682(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate683(.a(s_19), .b(gate176inter3), .O(gate176inter10));
  nor2  gate684(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate685(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate686(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1023(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1024(.a(gate180inter0), .b(s_68), .O(gate180inter1));
  and2  gate1025(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1026(.a(s_68), .O(gate180inter3));
  inv1  gate1027(.a(s_69), .O(gate180inter4));
  nand2 gate1028(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1029(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1030(.a(G507), .O(gate180inter7));
  inv1  gate1031(.a(G561), .O(gate180inter8));
  nand2 gate1032(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1033(.a(s_69), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1034(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1035(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1036(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate631(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate632(.a(gate182inter0), .b(s_12), .O(gate182inter1));
  and2  gate633(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate634(.a(s_12), .O(gate182inter3));
  inv1  gate635(.a(s_13), .O(gate182inter4));
  nand2 gate636(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate637(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate638(.a(G513), .O(gate182inter7));
  inv1  gate639(.a(G564), .O(gate182inter8));
  nand2 gate640(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate641(.a(s_13), .b(gate182inter3), .O(gate182inter10));
  nor2  gate642(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate643(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate644(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate841(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate842(.a(gate186inter0), .b(s_42), .O(gate186inter1));
  and2  gate843(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate844(.a(s_42), .O(gate186inter3));
  inv1  gate845(.a(s_43), .O(gate186inter4));
  nand2 gate846(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate847(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate848(.a(G572), .O(gate186inter7));
  inv1  gate849(.a(G573), .O(gate186inter8));
  nand2 gate850(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate851(.a(s_43), .b(gate186inter3), .O(gate186inter10));
  nor2  gate852(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate853(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate854(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate617(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate618(.a(gate190inter0), .b(s_10), .O(gate190inter1));
  and2  gate619(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate620(.a(s_10), .O(gate190inter3));
  inv1  gate621(.a(s_11), .O(gate190inter4));
  nand2 gate622(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate623(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate624(.a(G580), .O(gate190inter7));
  inv1  gate625(.a(G581), .O(gate190inter8));
  nand2 gate626(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate627(.a(s_11), .b(gate190inter3), .O(gate190inter10));
  nor2  gate628(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate629(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate630(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate799(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate800(.a(gate191inter0), .b(s_36), .O(gate191inter1));
  and2  gate801(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate802(.a(s_36), .O(gate191inter3));
  inv1  gate803(.a(s_37), .O(gate191inter4));
  nand2 gate804(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate805(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate806(.a(G582), .O(gate191inter7));
  inv1  gate807(.a(G583), .O(gate191inter8));
  nand2 gate808(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate809(.a(s_37), .b(gate191inter3), .O(gate191inter10));
  nor2  gate810(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate811(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate812(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1177(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1178(.a(gate192inter0), .b(s_90), .O(gate192inter1));
  and2  gate1179(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1180(.a(s_90), .O(gate192inter3));
  inv1  gate1181(.a(s_91), .O(gate192inter4));
  nand2 gate1182(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1183(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1184(.a(G584), .O(gate192inter7));
  inv1  gate1185(.a(G585), .O(gate192inter8));
  nand2 gate1186(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1187(.a(s_91), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1188(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1189(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1190(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1037(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1038(.a(gate198inter0), .b(s_70), .O(gate198inter1));
  and2  gate1039(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1040(.a(s_70), .O(gate198inter3));
  inv1  gate1041(.a(s_71), .O(gate198inter4));
  nand2 gate1042(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1043(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1044(.a(G596), .O(gate198inter7));
  inv1  gate1045(.a(G597), .O(gate198inter8));
  nand2 gate1046(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1047(.a(s_71), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1048(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1049(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1050(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1303(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1304(.a(gate218inter0), .b(s_108), .O(gate218inter1));
  and2  gate1305(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1306(.a(s_108), .O(gate218inter3));
  inv1  gate1307(.a(s_109), .O(gate218inter4));
  nand2 gate1308(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1309(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1310(.a(G627), .O(gate218inter7));
  inv1  gate1311(.a(G678), .O(gate218inter8));
  nand2 gate1312(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1313(.a(s_109), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1314(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1315(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1316(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate589(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate590(.a(gate235inter0), .b(s_6), .O(gate235inter1));
  and2  gate591(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate592(.a(s_6), .O(gate235inter3));
  inv1  gate593(.a(s_7), .O(gate235inter4));
  nand2 gate594(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate595(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate596(.a(G248), .O(gate235inter7));
  inv1  gate597(.a(G724), .O(gate235inter8));
  nand2 gate598(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate599(.a(s_7), .b(gate235inter3), .O(gate235inter10));
  nor2  gate600(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate601(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate602(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate603(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate604(.a(gate240inter0), .b(s_8), .O(gate240inter1));
  and2  gate605(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate606(.a(s_8), .O(gate240inter3));
  inv1  gate607(.a(s_9), .O(gate240inter4));
  nand2 gate608(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate609(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate610(.a(G263), .O(gate240inter7));
  inv1  gate611(.a(G715), .O(gate240inter8));
  nand2 gate612(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate613(.a(s_9), .b(gate240inter3), .O(gate240inter10));
  nor2  gate614(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate615(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate616(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate869(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate870(.a(gate248inter0), .b(s_46), .O(gate248inter1));
  and2  gate871(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate872(.a(s_46), .O(gate248inter3));
  inv1  gate873(.a(s_47), .O(gate248inter4));
  nand2 gate874(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate875(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate876(.a(G727), .O(gate248inter7));
  inv1  gate877(.a(G739), .O(gate248inter8));
  nand2 gate878(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate879(.a(s_47), .b(gate248inter3), .O(gate248inter10));
  nor2  gate880(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate881(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate882(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate883(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate884(.a(gate266inter0), .b(s_48), .O(gate266inter1));
  and2  gate885(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate886(.a(s_48), .O(gate266inter3));
  inv1  gate887(.a(s_49), .O(gate266inter4));
  nand2 gate888(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate889(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate890(.a(G645), .O(gate266inter7));
  inv1  gate891(.a(G773), .O(gate266inter8));
  nand2 gate892(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate893(.a(s_49), .b(gate266inter3), .O(gate266inter10));
  nor2  gate894(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate895(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate896(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate771(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate772(.a(gate283inter0), .b(s_32), .O(gate283inter1));
  and2  gate773(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate774(.a(s_32), .O(gate283inter3));
  inv1  gate775(.a(s_33), .O(gate283inter4));
  nand2 gate776(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate777(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate778(.a(G657), .O(gate283inter7));
  inv1  gate779(.a(G809), .O(gate283inter8));
  nand2 gate780(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate781(.a(s_33), .b(gate283inter3), .O(gate283inter10));
  nor2  gate782(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate783(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate784(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate939(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate940(.a(gate388inter0), .b(s_56), .O(gate388inter1));
  and2  gate941(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate942(.a(s_56), .O(gate388inter3));
  inv1  gate943(.a(s_57), .O(gate388inter4));
  nand2 gate944(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate945(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate946(.a(G2), .O(gate388inter7));
  inv1  gate947(.a(G1039), .O(gate388inter8));
  nand2 gate948(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate949(.a(s_57), .b(gate388inter3), .O(gate388inter10));
  nor2  gate950(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate951(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate952(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate813(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate814(.a(gate394inter0), .b(s_38), .O(gate394inter1));
  and2  gate815(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate816(.a(s_38), .O(gate394inter3));
  inv1  gate817(.a(s_39), .O(gate394inter4));
  nand2 gate818(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate819(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate820(.a(G8), .O(gate394inter7));
  inv1  gate821(.a(G1057), .O(gate394inter8));
  nand2 gate822(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate823(.a(s_39), .b(gate394inter3), .O(gate394inter10));
  nor2  gate824(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate825(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate826(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1219(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1220(.a(gate406inter0), .b(s_96), .O(gate406inter1));
  and2  gate1221(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1222(.a(s_96), .O(gate406inter3));
  inv1  gate1223(.a(s_97), .O(gate406inter4));
  nand2 gate1224(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1225(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1226(.a(G20), .O(gate406inter7));
  inv1  gate1227(.a(G1093), .O(gate406inter8));
  nand2 gate1228(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1229(.a(s_97), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1230(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1231(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1232(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1205(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1206(.a(gate407inter0), .b(s_94), .O(gate407inter1));
  and2  gate1207(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1208(.a(s_94), .O(gate407inter3));
  inv1  gate1209(.a(s_95), .O(gate407inter4));
  nand2 gate1210(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1211(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1212(.a(G21), .O(gate407inter7));
  inv1  gate1213(.a(G1096), .O(gate407inter8));
  nand2 gate1214(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1215(.a(s_95), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1216(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1217(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1218(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1093(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1094(.a(gate408inter0), .b(s_78), .O(gate408inter1));
  and2  gate1095(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1096(.a(s_78), .O(gate408inter3));
  inv1  gate1097(.a(s_79), .O(gate408inter4));
  nand2 gate1098(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1099(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1100(.a(G22), .O(gate408inter7));
  inv1  gate1101(.a(G1099), .O(gate408inter8));
  nand2 gate1102(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1103(.a(s_79), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1104(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1105(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1106(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate645(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate646(.a(gate411inter0), .b(s_14), .O(gate411inter1));
  and2  gate647(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate648(.a(s_14), .O(gate411inter3));
  inv1  gate649(.a(s_15), .O(gate411inter4));
  nand2 gate650(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate651(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate652(.a(G25), .O(gate411inter7));
  inv1  gate653(.a(G1108), .O(gate411inter8));
  nand2 gate654(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate655(.a(s_15), .b(gate411inter3), .O(gate411inter10));
  nor2  gate656(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate657(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate658(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate785(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate786(.a(gate414inter0), .b(s_34), .O(gate414inter1));
  and2  gate787(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate788(.a(s_34), .O(gate414inter3));
  inv1  gate789(.a(s_35), .O(gate414inter4));
  nand2 gate790(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate791(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate792(.a(G28), .O(gate414inter7));
  inv1  gate793(.a(G1117), .O(gate414inter8));
  nand2 gate794(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate795(.a(s_35), .b(gate414inter3), .O(gate414inter10));
  nor2  gate796(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate797(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate798(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1289(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1290(.a(gate418inter0), .b(s_106), .O(gate418inter1));
  and2  gate1291(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1292(.a(s_106), .O(gate418inter3));
  inv1  gate1293(.a(s_107), .O(gate418inter4));
  nand2 gate1294(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1295(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1296(.a(G32), .O(gate418inter7));
  inv1  gate1297(.a(G1129), .O(gate418inter8));
  nand2 gate1298(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1299(.a(s_107), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1300(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1301(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1302(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate967(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate968(.a(gate423inter0), .b(s_60), .O(gate423inter1));
  and2  gate969(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate970(.a(s_60), .O(gate423inter3));
  inv1  gate971(.a(s_61), .O(gate423inter4));
  nand2 gate972(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate973(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate974(.a(G3), .O(gate423inter7));
  inv1  gate975(.a(G1138), .O(gate423inter8));
  nand2 gate976(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate977(.a(s_61), .b(gate423inter3), .O(gate423inter10));
  nor2  gate978(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate979(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate980(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate827(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate828(.a(gate424inter0), .b(s_40), .O(gate424inter1));
  and2  gate829(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate830(.a(s_40), .O(gate424inter3));
  inv1  gate831(.a(s_41), .O(gate424inter4));
  nand2 gate832(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate833(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate834(.a(G1042), .O(gate424inter7));
  inv1  gate835(.a(G1138), .O(gate424inter8));
  nand2 gate836(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate837(.a(s_41), .b(gate424inter3), .O(gate424inter10));
  nor2  gate838(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate839(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate840(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate715(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate716(.a(gate435inter0), .b(s_24), .O(gate435inter1));
  and2  gate717(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate718(.a(s_24), .O(gate435inter3));
  inv1  gate719(.a(s_25), .O(gate435inter4));
  nand2 gate720(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate721(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate722(.a(G9), .O(gate435inter7));
  inv1  gate723(.a(G1156), .O(gate435inter8));
  nand2 gate724(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate725(.a(s_25), .b(gate435inter3), .O(gate435inter10));
  nor2  gate726(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate727(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate728(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1317(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1318(.a(gate443inter0), .b(s_110), .O(gate443inter1));
  and2  gate1319(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1320(.a(s_110), .O(gate443inter3));
  inv1  gate1321(.a(s_111), .O(gate443inter4));
  nand2 gate1322(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1323(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1324(.a(G13), .O(gate443inter7));
  inv1  gate1325(.a(G1168), .O(gate443inter8));
  nand2 gate1326(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1327(.a(s_111), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1328(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1329(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1330(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1247(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1248(.a(gate465inter0), .b(s_100), .O(gate465inter1));
  and2  gate1249(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1250(.a(s_100), .O(gate465inter3));
  inv1  gate1251(.a(s_101), .O(gate465inter4));
  nand2 gate1252(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1253(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1254(.a(G24), .O(gate465inter7));
  inv1  gate1255(.a(G1201), .O(gate465inter8));
  nand2 gate1256(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1257(.a(s_101), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1258(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1259(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1260(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate757(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate758(.a(gate472inter0), .b(s_30), .O(gate472inter1));
  and2  gate759(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate760(.a(s_30), .O(gate472inter3));
  inv1  gate761(.a(s_31), .O(gate472inter4));
  nand2 gate762(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate763(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate764(.a(G1114), .O(gate472inter7));
  inv1  gate765(.a(G1210), .O(gate472inter8));
  nand2 gate766(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate767(.a(s_31), .b(gate472inter3), .O(gate472inter10));
  nor2  gate768(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate769(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate770(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate925(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate926(.a(gate482inter0), .b(s_54), .O(gate482inter1));
  and2  gate927(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate928(.a(s_54), .O(gate482inter3));
  inv1  gate929(.a(s_55), .O(gate482inter4));
  nand2 gate930(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate931(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate932(.a(G1129), .O(gate482inter7));
  inv1  gate933(.a(G1225), .O(gate482inter8));
  nand2 gate934(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate935(.a(s_55), .b(gate482inter3), .O(gate482inter10));
  nor2  gate936(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate937(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate938(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate855(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate856(.a(gate483inter0), .b(s_44), .O(gate483inter1));
  and2  gate857(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate858(.a(s_44), .O(gate483inter3));
  inv1  gate859(.a(s_45), .O(gate483inter4));
  nand2 gate860(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate861(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate862(.a(G1228), .O(gate483inter7));
  inv1  gate863(.a(G1229), .O(gate483inter8));
  nand2 gate864(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate865(.a(s_45), .b(gate483inter3), .O(gate483inter10));
  nor2  gate866(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate867(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate868(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate981(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate982(.a(gate494inter0), .b(s_62), .O(gate494inter1));
  and2  gate983(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate984(.a(s_62), .O(gate494inter3));
  inv1  gate985(.a(s_63), .O(gate494inter4));
  nand2 gate986(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate987(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate988(.a(G1250), .O(gate494inter7));
  inv1  gate989(.a(G1251), .O(gate494inter8));
  nand2 gate990(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate991(.a(s_63), .b(gate494inter3), .O(gate494inter10));
  nor2  gate992(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate993(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate994(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate897(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate898(.a(gate497inter0), .b(s_50), .O(gate497inter1));
  and2  gate899(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate900(.a(s_50), .O(gate497inter3));
  inv1  gate901(.a(s_51), .O(gate497inter4));
  nand2 gate902(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate903(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate904(.a(G1256), .O(gate497inter7));
  inv1  gate905(.a(G1257), .O(gate497inter8));
  nand2 gate906(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate907(.a(s_51), .b(gate497inter3), .O(gate497inter10));
  nor2  gate908(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate909(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate910(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate995(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate996(.a(gate506inter0), .b(s_64), .O(gate506inter1));
  and2  gate997(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate998(.a(s_64), .O(gate506inter3));
  inv1  gate999(.a(s_65), .O(gate506inter4));
  nand2 gate1000(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1001(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1002(.a(G1274), .O(gate506inter7));
  inv1  gate1003(.a(G1275), .O(gate506inter8));
  nand2 gate1004(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1005(.a(s_65), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1006(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1007(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1008(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule