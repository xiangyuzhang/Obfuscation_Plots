module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate911(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate912(.a(gate11inter0), .b(s_52), .O(gate11inter1));
  and2  gate913(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate914(.a(s_52), .O(gate11inter3));
  inv1  gate915(.a(s_53), .O(gate11inter4));
  nand2 gate916(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate917(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate918(.a(G5), .O(gate11inter7));
  inv1  gate919(.a(G6), .O(gate11inter8));
  nand2 gate920(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate921(.a(s_53), .b(gate11inter3), .O(gate11inter10));
  nor2  gate922(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate923(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate924(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1415(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1416(.a(gate15inter0), .b(s_124), .O(gate15inter1));
  and2  gate1417(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1418(.a(s_124), .O(gate15inter3));
  inv1  gate1419(.a(s_125), .O(gate15inter4));
  nand2 gate1420(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1421(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1422(.a(G13), .O(gate15inter7));
  inv1  gate1423(.a(G14), .O(gate15inter8));
  nand2 gate1424(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1425(.a(s_125), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1426(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1427(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1428(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1555(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1556(.a(gate17inter0), .b(s_144), .O(gate17inter1));
  and2  gate1557(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1558(.a(s_144), .O(gate17inter3));
  inv1  gate1559(.a(s_145), .O(gate17inter4));
  nand2 gate1560(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1561(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1562(.a(G17), .O(gate17inter7));
  inv1  gate1563(.a(G18), .O(gate17inter8));
  nand2 gate1564(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1565(.a(s_145), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1566(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1567(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1568(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1121(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1122(.a(gate31inter0), .b(s_82), .O(gate31inter1));
  and2  gate1123(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1124(.a(s_82), .O(gate31inter3));
  inv1  gate1125(.a(s_83), .O(gate31inter4));
  nand2 gate1126(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1127(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1128(.a(G4), .O(gate31inter7));
  inv1  gate1129(.a(G8), .O(gate31inter8));
  nand2 gate1130(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1131(.a(s_83), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1132(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1133(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1134(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate631(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate632(.a(gate35inter0), .b(s_12), .O(gate35inter1));
  and2  gate633(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate634(.a(s_12), .O(gate35inter3));
  inv1  gate635(.a(s_13), .O(gate35inter4));
  nand2 gate636(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate637(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate638(.a(G18), .O(gate35inter7));
  inv1  gate639(.a(G22), .O(gate35inter8));
  nand2 gate640(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate641(.a(s_13), .b(gate35inter3), .O(gate35inter10));
  nor2  gate642(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate643(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate644(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1345(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1346(.a(gate36inter0), .b(s_114), .O(gate36inter1));
  and2  gate1347(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1348(.a(s_114), .O(gate36inter3));
  inv1  gate1349(.a(s_115), .O(gate36inter4));
  nand2 gate1350(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1351(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1352(.a(G26), .O(gate36inter7));
  inv1  gate1353(.a(G30), .O(gate36inter8));
  nand2 gate1354(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1355(.a(s_115), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1356(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1357(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1358(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1051(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1052(.a(gate39inter0), .b(s_72), .O(gate39inter1));
  and2  gate1053(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1054(.a(s_72), .O(gate39inter3));
  inv1  gate1055(.a(s_73), .O(gate39inter4));
  nand2 gate1056(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1057(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1058(.a(G20), .O(gate39inter7));
  inv1  gate1059(.a(G24), .O(gate39inter8));
  nand2 gate1060(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1061(.a(s_73), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1062(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1063(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1064(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate617(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate618(.a(gate40inter0), .b(s_10), .O(gate40inter1));
  and2  gate619(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate620(.a(s_10), .O(gate40inter3));
  inv1  gate621(.a(s_11), .O(gate40inter4));
  nand2 gate622(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate623(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate624(.a(G28), .O(gate40inter7));
  inv1  gate625(.a(G32), .O(gate40inter8));
  nand2 gate626(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate627(.a(s_11), .b(gate40inter3), .O(gate40inter10));
  nor2  gate628(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate629(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate630(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1471(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1472(.a(gate43inter0), .b(s_132), .O(gate43inter1));
  and2  gate1473(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1474(.a(s_132), .O(gate43inter3));
  inv1  gate1475(.a(s_133), .O(gate43inter4));
  nand2 gate1476(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1477(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1478(.a(G3), .O(gate43inter7));
  inv1  gate1479(.a(G269), .O(gate43inter8));
  nand2 gate1480(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1481(.a(s_133), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1482(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1483(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1484(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1513(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1514(.a(gate45inter0), .b(s_138), .O(gate45inter1));
  and2  gate1515(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1516(.a(s_138), .O(gate45inter3));
  inv1  gate1517(.a(s_139), .O(gate45inter4));
  nand2 gate1518(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1519(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1520(.a(G5), .O(gate45inter7));
  inv1  gate1521(.a(G272), .O(gate45inter8));
  nand2 gate1522(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1523(.a(s_139), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1524(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1525(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1526(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1037(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1038(.a(gate46inter0), .b(s_70), .O(gate46inter1));
  and2  gate1039(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1040(.a(s_70), .O(gate46inter3));
  inv1  gate1041(.a(s_71), .O(gate46inter4));
  nand2 gate1042(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1043(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1044(.a(G6), .O(gate46inter7));
  inv1  gate1045(.a(G272), .O(gate46inter8));
  nand2 gate1046(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1047(.a(s_71), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1048(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1049(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1050(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1429(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1430(.a(gate51inter0), .b(s_126), .O(gate51inter1));
  and2  gate1431(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1432(.a(s_126), .O(gate51inter3));
  inv1  gate1433(.a(s_127), .O(gate51inter4));
  nand2 gate1434(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1435(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1436(.a(G11), .O(gate51inter7));
  inv1  gate1437(.a(G281), .O(gate51inter8));
  nand2 gate1438(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1439(.a(s_127), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1440(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1441(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1442(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate659(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate660(.a(gate53inter0), .b(s_16), .O(gate53inter1));
  and2  gate661(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate662(.a(s_16), .O(gate53inter3));
  inv1  gate663(.a(s_17), .O(gate53inter4));
  nand2 gate664(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate665(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate666(.a(G13), .O(gate53inter7));
  inv1  gate667(.a(G284), .O(gate53inter8));
  nand2 gate668(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate669(.a(s_17), .b(gate53inter3), .O(gate53inter10));
  nor2  gate670(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate671(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate672(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate785(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate786(.a(gate59inter0), .b(s_34), .O(gate59inter1));
  and2  gate787(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate788(.a(s_34), .O(gate59inter3));
  inv1  gate789(.a(s_35), .O(gate59inter4));
  nand2 gate790(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate791(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate792(.a(G19), .O(gate59inter7));
  inv1  gate793(.a(G293), .O(gate59inter8));
  nand2 gate794(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate795(.a(s_35), .b(gate59inter3), .O(gate59inter10));
  nor2  gate796(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate797(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate798(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate701(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate702(.a(gate65inter0), .b(s_22), .O(gate65inter1));
  and2  gate703(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate704(.a(s_22), .O(gate65inter3));
  inv1  gate705(.a(s_23), .O(gate65inter4));
  nand2 gate706(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate707(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate708(.a(G25), .O(gate65inter7));
  inv1  gate709(.a(G302), .O(gate65inter8));
  nand2 gate710(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate711(.a(s_23), .b(gate65inter3), .O(gate65inter10));
  nor2  gate712(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate713(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate714(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1065(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1066(.a(gate66inter0), .b(s_74), .O(gate66inter1));
  and2  gate1067(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1068(.a(s_74), .O(gate66inter3));
  inv1  gate1069(.a(s_75), .O(gate66inter4));
  nand2 gate1070(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1071(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1072(.a(G26), .O(gate66inter7));
  inv1  gate1073(.a(G302), .O(gate66inter8));
  nand2 gate1074(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1075(.a(s_75), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1076(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1077(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1078(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1597(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1598(.a(gate67inter0), .b(s_150), .O(gate67inter1));
  and2  gate1599(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1600(.a(s_150), .O(gate67inter3));
  inv1  gate1601(.a(s_151), .O(gate67inter4));
  nand2 gate1602(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1603(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1604(.a(G27), .O(gate67inter7));
  inv1  gate1605(.a(G305), .O(gate67inter8));
  nand2 gate1606(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1607(.a(s_151), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1608(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1609(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1610(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1639(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1640(.a(gate68inter0), .b(s_156), .O(gate68inter1));
  and2  gate1641(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1642(.a(s_156), .O(gate68inter3));
  inv1  gate1643(.a(s_157), .O(gate68inter4));
  nand2 gate1644(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1645(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1646(.a(G28), .O(gate68inter7));
  inv1  gate1647(.a(G305), .O(gate68inter8));
  nand2 gate1648(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1649(.a(s_157), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1650(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1651(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1652(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1401(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1402(.a(gate70inter0), .b(s_122), .O(gate70inter1));
  and2  gate1403(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1404(.a(s_122), .O(gate70inter3));
  inv1  gate1405(.a(s_123), .O(gate70inter4));
  nand2 gate1406(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1407(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1408(.a(G30), .O(gate70inter7));
  inv1  gate1409(.a(G308), .O(gate70inter8));
  nand2 gate1410(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1411(.a(s_123), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1412(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1413(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1414(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1583(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1584(.a(gate75inter0), .b(s_148), .O(gate75inter1));
  and2  gate1585(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1586(.a(s_148), .O(gate75inter3));
  inv1  gate1587(.a(s_149), .O(gate75inter4));
  nand2 gate1588(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1589(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1590(.a(G9), .O(gate75inter7));
  inv1  gate1591(.a(G317), .O(gate75inter8));
  nand2 gate1592(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1593(.a(s_149), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1594(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1595(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1596(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate589(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate590(.a(gate81inter0), .b(s_6), .O(gate81inter1));
  and2  gate591(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate592(.a(s_6), .O(gate81inter3));
  inv1  gate593(.a(s_7), .O(gate81inter4));
  nand2 gate594(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate595(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate596(.a(G3), .O(gate81inter7));
  inv1  gate597(.a(G326), .O(gate81inter8));
  nand2 gate598(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate599(.a(s_7), .b(gate81inter3), .O(gate81inter10));
  nor2  gate600(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate601(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate602(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1023(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1024(.a(gate82inter0), .b(s_68), .O(gate82inter1));
  and2  gate1025(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1026(.a(s_68), .O(gate82inter3));
  inv1  gate1027(.a(s_69), .O(gate82inter4));
  nand2 gate1028(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1029(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1030(.a(G7), .O(gate82inter7));
  inv1  gate1031(.a(G326), .O(gate82inter8));
  nand2 gate1032(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1033(.a(s_69), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1034(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1035(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1036(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1303(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1304(.a(gate86inter0), .b(s_108), .O(gate86inter1));
  and2  gate1305(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1306(.a(s_108), .O(gate86inter3));
  inv1  gate1307(.a(s_109), .O(gate86inter4));
  nand2 gate1308(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1309(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1310(.a(G8), .O(gate86inter7));
  inv1  gate1311(.a(G332), .O(gate86inter8));
  nand2 gate1312(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1313(.a(s_109), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1314(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1315(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1316(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1541(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1542(.a(gate87inter0), .b(s_142), .O(gate87inter1));
  and2  gate1543(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1544(.a(s_142), .O(gate87inter3));
  inv1  gate1545(.a(s_143), .O(gate87inter4));
  nand2 gate1546(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1547(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1548(.a(G12), .O(gate87inter7));
  inv1  gate1549(.a(G335), .O(gate87inter8));
  nand2 gate1550(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1551(.a(s_143), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1552(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1553(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1554(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1611(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1612(.a(gate88inter0), .b(s_152), .O(gate88inter1));
  and2  gate1613(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1614(.a(s_152), .O(gate88inter3));
  inv1  gate1615(.a(s_153), .O(gate88inter4));
  nand2 gate1616(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1617(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1618(.a(G16), .O(gate88inter7));
  inv1  gate1619(.a(G335), .O(gate88inter8));
  nand2 gate1620(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1621(.a(s_153), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1622(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1623(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1624(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate547(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate548(.a(gate95inter0), .b(s_0), .O(gate95inter1));
  and2  gate549(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate550(.a(s_0), .O(gate95inter3));
  inv1  gate551(.a(s_1), .O(gate95inter4));
  nand2 gate552(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate553(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate554(.a(G26), .O(gate95inter7));
  inv1  gate555(.a(G347), .O(gate95inter8));
  nand2 gate556(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate557(.a(s_1), .b(gate95inter3), .O(gate95inter10));
  nor2  gate558(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate559(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate560(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1009(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1010(.a(gate100inter0), .b(s_66), .O(gate100inter1));
  and2  gate1011(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1012(.a(s_66), .O(gate100inter3));
  inv1  gate1013(.a(s_67), .O(gate100inter4));
  nand2 gate1014(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1015(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1016(.a(G31), .O(gate100inter7));
  inv1  gate1017(.a(G353), .O(gate100inter8));
  nand2 gate1018(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1019(.a(s_67), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1020(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1021(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1022(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1569(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1570(.a(gate105inter0), .b(s_146), .O(gate105inter1));
  and2  gate1571(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1572(.a(s_146), .O(gate105inter3));
  inv1  gate1573(.a(s_147), .O(gate105inter4));
  nand2 gate1574(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1575(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1576(.a(G362), .O(gate105inter7));
  inv1  gate1577(.a(G363), .O(gate105inter8));
  nand2 gate1578(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1579(.a(s_147), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1580(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1581(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1582(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1359(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1360(.a(gate123inter0), .b(s_116), .O(gate123inter1));
  and2  gate1361(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1362(.a(s_116), .O(gate123inter3));
  inv1  gate1363(.a(s_117), .O(gate123inter4));
  nand2 gate1364(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1365(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1366(.a(G398), .O(gate123inter7));
  inv1  gate1367(.a(G399), .O(gate123inter8));
  nand2 gate1368(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1369(.a(s_117), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1370(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1371(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1372(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1387(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1388(.a(gate133inter0), .b(s_120), .O(gate133inter1));
  and2  gate1389(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1390(.a(s_120), .O(gate133inter3));
  inv1  gate1391(.a(s_121), .O(gate133inter4));
  nand2 gate1392(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1393(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1394(.a(G418), .O(gate133inter7));
  inv1  gate1395(.a(G419), .O(gate133inter8));
  nand2 gate1396(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1397(.a(s_121), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1398(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1399(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1400(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1093(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1094(.a(gate136inter0), .b(s_78), .O(gate136inter1));
  and2  gate1095(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1096(.a(s_78), .O(gate136inter3));
  inv1  gate1097(.a(s_79), .O(gate136inter4));
  nand2 gate1098(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1099(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1100(.a(G424), .O(gate136inter7));
  inv1  gate1101(.a(G425), .O(gate136inter8));
  nand2 gate1102(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1103(.a(s_79), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1104(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1105(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1106(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate995(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate996(.a(gate149inter0), .b(s_64), .O(gate149inter1));
  and2  gate997(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate998(.a(s_64), .O(gate149inter3));
  inv1  gate999(.a(s_65), .O(gate149inter4));
  nand2 gate1000(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1001(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1002(.a(G498), .O(gate149inter7));
  inv1  gate1003(.a(G501), .O(gate149inter8));
  nand2 gate1004(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1005(.a(s_65), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1006(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1007(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1008(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1667(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1668(.a(gate151inter0), .b(s_160), .O(gate151inter1));
  and2  gate1669(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1670(.a(s_160), .O(gate151inter3));
  inv1  gate1671(.a(s_161), .O(gate151inter4));
  nand2 gate1672(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1673(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1674(.a(G510), .O(gate151inter7));
  inv1  gate1675(.a(G513), .O(gate151inter8));
  nand2 gate1676(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1677(.a(s_161), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1678(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1679(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1680(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate883(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate884(.a(gate155inter0), .b(s_48), .O(gate155inter1));
  and2  gate885(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate886(.a(s_48), .O(gate155inter3));
  inv1  gate887(.a(s_49), .O(gate155inter4));
  nand2 gate888(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate889(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate890(.a(G432), .O(gate155inter7));
  inv1  gate891(.a(G525), .O(gate155inter8));
  nand2 gate892(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate893(.a(s_49), .b(gate155inter3), .O(gate155inter10));
  nor2  gate894(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate895(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate896(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate981(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate982(.a(gate156inter0), .b(s_62), .O(gate156inter1));
  and2  gate983(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate984(.a(s_62), .O(gate156inter3));
  inv1  gate985(.a(s_63), .O(gate156inter4));
  nand2 gate986(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate987(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate988(.a(G435), .O(gate156inter7));
  inv1  gate989(.a(G525), .O(gate156inter8));
  nand2 gate990(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate991(.a(s_63), .b(gate156inter3), .O(gate156inter10));
  nor2  gate992(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate993(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate994(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate855(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate856(.a(gate159inter0), .b(s_44), .O(gate159inter1));
  and2  gate857(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate858(.a(s_44), .O(gate159inter3));
  inv1  gate859(.a(s_45), .O(gate159inter4));
  nand2 gate860(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate861(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate862(.a(G444), .O(gate159inter7));
  inv1  gate863(.a(G531), .O(gate159inter8));
  nand2 gate864(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate865(.a(s_45), .b(gate159inter3), .O(gate159inter10));
  nor2  gate866(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate867(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate868(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1499(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1500(.a(gate170inter0), .b(s_136), .O(gate170inter1));
  and2  gate1501(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1502(.a(s_136), .O(gate170inter3));
  inv1  gate1503(.a(s_137), .O(gate170inter4));
  nand2 gate1504(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1505(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1506(.a(G477), .O(gate170inter7));
  inv1  gate1507(.a(G546), .O(gate170inter8));
  nand2 gate1508(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1509(.a(s_137), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1510(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1511(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1512(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate743(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate744(.a(gate172inter0), .b(s_28), .O(gate172inter1));
  and2  gate745(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate746(.a(s_28), .O(gate172inter3));
  inv1  gate747(.a(s_29), .O(gate172inter4));
  nand2 gate748(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate749(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate750(.a(G483), .O(gate172inter7));
  inv1  gate751(.a(G549), .O(gate172inter8));
  nand2 gate752(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate753(.a(s_29), .b(gate172inter3), .O(gate172inter10));
  nor2  gate754(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate755(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate756(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate729(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate730(.a(gate177inter0), .b(s_26), .O(gate177inter1));
  and2  gate731(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate732(.a(s_26), .O(gate177inter3));
  inv1  gate733(.a(s_27), .O(gate177inter4));
  nand2 gate734(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate735(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate736(.a(G498), .O(gate177inter7));
  inv1  gate737(.a(G558), .O(gate177inter8));
  nand2 gate738(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate739(.a(s_27), .b(gate177inter3), .O(gate177inter10));
  nor2  gate740(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate741(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate742(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate841(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate842(.a(gate183inter0), .b(s_42), .O(gate183inter1));
  and2  gate843(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate844(.a(s_42), .O(gate183inter3));
  inv1  gate845(.a(s_43), .O(gate183inter4));
  nand2 gate846(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate847(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate848(.a(G516), .O(gate183inter7));
  inv1  gate849(.a(G567), .O(gate183inter8));
  nand2 gate850(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate851(.a(s_43), .b(gate183inter3), .O(gate183inter10));
  nor2  gate852(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate853(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate854(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1135(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1136(.a(gate186inter0), .b(s_84), .O(gate186inter1));
  and2  gate1137(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1138(.a(s_84), .O(gate186inter3));
  inv1  gate1139(.a(s_85), .O(gate186inter4));
  nand2 gate1140(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1141(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1142(.a(G572), .O(gate186inter7));
  inv1  gate1143(.a(G573), .O(gate186inter8));
  nand2 gate1144(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1145(.a(s_85), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1146(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1147(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1148(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1107(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1108(.a(gate214inter0), .b(s_80), .O(gate214inter1));
  and2  gate1109(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1110(.a(s_80), .O(gate214inter3));
  inv1  gate1111(.a(s_81), .O(gate214inter4));
  nand2 gate1112(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1113(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1114(.a(G612), .O(gate214inter7));
  inv1  gate1115(.a(G672), .O(gate214inter8));
  nand2 gate1116(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1117(.a(s_81), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1118(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1119(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1120(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate645(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate646(.a(gate225inter0), .b(s_14), .O(gate225inter1));
  and2  gate647(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate648(.a(s_14), .O(gate225inter3));
  inv1  gate649(.a(s_15), .O(gate225inter4));
  nand2 gate650(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate651(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate652(.a(G690), .O(gate225inter7));
  inv1  gate653(.a(G691), .O(gate225inter8));
  nand2 gate654(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate655(.a(s_15), .b(gate225inter3), .O(gate225inter10));
  nor2  gate656(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate657(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate658(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1191(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1192(.a(gate226inter0), .b(s_92), .O(gate226inter1));
  and2  gate1193(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1194(.a(s_92), .O(gate226inter3));
  inv1  gate1195(.a(s_93), .O(gate226inter4));
  nand2 gate1196(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1197(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1198(.a(G692), .O(gate226inter7));
  inv1  gate1199(.a(G693), .O(gate226inter8));
  nand2 gate1200(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1201(.a(s_93), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1202(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1203(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1204(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate869(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate870(.a(gate234inter0), .b(s_46), .O(gate234inter1));
  and2  gate871(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate872(.a(s_46), .O(gate234inter3));
  inv1  gate873(.a(s_47), .O(gate234inter4));
  nand2 gate874(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate875(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate876(.a(G245), .O(gate234inter7));
  inv1  gate877(.a(G721), .O(gate234inter8));
  nand2 gate878(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate879(.a(s_47), .b(gate234inter3), .O(gate234inter10));
  nor2  gate880(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate881(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate882(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate603(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate604(.a(gate235inter0), .b(s_8), .O(gate235inter1));
  and2  gate605(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate606(.a(s_8), .O(gate235inter3));
  inv1  gate607(.a(s_9), .O(gate235inter4));
  nand2 gate608(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate609(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate610(.a(G248), .O(gate235inter7));
  inv1  gate611(.a(G724), .O(gate235inter8));
  nand2 gate612(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate613(.a(s_9), .b(gate235inter3), .O(gate235inter10));
  nor2  gate614(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate615(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate616(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate953(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate954(.a(gate236inter0), .b(s_58), .O(gate236inter1));
  and2  gate955(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate956(.a(s_58), .O(gate236inter3));
  inv1  gate957(.a(s_59), .O(gate236inter4));
  nand2 gate958(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate959(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate960(.a(G251), .O(gate236inter7));
  inv1  gate961(.a(G727), .O(gate236inter8));
  nand2 gate962(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate963(.a(s_59), .b(gate236inter3), .O(gate236inter10));
  nor2  gate964(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate965(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate966(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate813(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate814(.a(gate241inter0), .b(s_38), .O(gate241inter1));
  and2  gate815(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate816(.a(s_38), .O(gate241inter3));
  inv1  gate817(.a(s_39), .O(gate241inter4));
  nand2 gate818(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate819(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate820(.a(G242), .O(gate241inter7));
  inv1  gate821(.a(G730), .O(gate241inter8));
  nand2 gate822(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate823(.a(s_39), .b(gate241inter3), .O(gate241inter10));
  nor2  gate824(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate825(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate826(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate925(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate926(.a(gate247inter0), .b(s_54), .O(gate247inter1));
  and2  gate927(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate928(.a(s_54), .O(gate247inter3));
  inv1  gate929(.a(s_55), .O(gate247inter4));
  nand2 gate930(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate931(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate932(.a(G251), .O(gate247inter7));
  inv1  gate933(.a(G739), .O(gate247inter8));
  nand2 gate934(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate935(.a(s_55), .b(gate247inter3), .O(gate247inter10));
  nor2  gate936(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate937(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate938(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate561(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate562(.a(gate253inter0), .b(s_2), .O(gate253inter1));
  and2  gate563(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate564(.a(s_2), .O(gate253inter3));
  inv1  gate565(.a(s_3), .O(gate253inter4));
  nand2 gate566(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate567(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate568(.a(G260), .O(gate253inter7));
  inv1  gate569(.a(G748), .O(gate253inter8));
  nand2 gate570(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate571(.a(s_3), .b(gate253inter3), .O(gate253inter10));
  nor2  gate572(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate573(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate574(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate757(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate758(.a(gate257inter0), .b(s_30), .O(gate257inter1));
  and2  gate759(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate760(.a(s_30), .O(gate257inter3));
  inv1  gate761(.a(s_31), .O(gate257inter4));
  nand2 gate762(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate763(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate764(.a(G754), .O(gate257inter7));
  inv1  gate765(.a(G755), .O(gate257inter8));
  nand2 gate766(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate767(.a(s_31), .b(gate257inter3), .O(gate257inter10));
  nor2  gate768(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate769(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate770(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1457(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1458(.a(gate260inter0), .b(s_130), .O(gate260inter1));
  and2  gate1459(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1460(.a(s_130), .O(gate260inter3));
  inv1  gate1461(.a(s_131), .O(gate260inter4));
  nand2 gate1462(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1463(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1464(.a(G760), .O(gate260inter7));
  inv1  gate1465(.a(G761), .O(gate260inter8));
  nand2 gate1466(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1467(.a(s_131), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1468(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1469(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1470(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate673(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate674(.a(gate261inter0), .b(s_18), .O(gate261inter1));
  and2  gate675(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate676(.a(s_18), .O(gate261inter3));
  inv1  gate677(.a(s_19), .O(gate261inter4));
  nand2 gate678(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate679(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate680(.a(G762), .O(gate261inter7));
  inv1  gate681(.a(G763), .O(gate261inter8));
  nand2 gate682(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate683(.a(s_19), .b(gate261inter3), .O(gate261inter10));
  nor2  gate684(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate685(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate686(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1527(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1528(.a(gate263inter0), .b(s_140), .O(gate263inter1));
  and2  gate1529(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1530(.a(s_140), .O(gate263inter3));
  inv1  gate1531(.a(s_141), .O(gate263inter4));
  nand2 gate1532(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1533(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1534(.a(G766), .O(gate263inter7));
  inv1  gate1535(.a(G767), .O(gate263inter8));
  nand2 gate1536(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1537(.a(s_141), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1538(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1539(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1540(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1317(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1318(.a(gate286inter0), .b(s_110), .O(gate286inter1));
  and2  gate1319(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1320(.a(s_110), .O(gate286inter3));
  inv1  gate1321(.a(s_111), .O(gate286inter4));
  nand2 gate1322(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1323(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1324(.a(G788), .O(gate286inter7));
  inv1  gate1325(.a(G812), .O(gate286inter8));
  nand2 gate1326(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1327(.a(s_111), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1328(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1329(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1330(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate575(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate576(.a(gate390inter0), .b(s_4), .O(gate390inter1));
  and2  gate577(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate578(.a(s_4), .O(gate390inter3));
  inv1  gate579(.a(s_5), .O(gate390inter4));
  nand2 gate580(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate581(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate582(.a(G4), .O(gate390inter7));
  inv1  gate583(.a(G1045), .O(gate390inter8));
  nand2 gate584(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate585(.a(s_5), .b(gate390inter3), .O(gate390inter10));
  nor2  gate586(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate587(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate588(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate897(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate898(.a(gate395inter0), .b(s_50), .O(gate395inter1));
  and2  gate899(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate900(.a(s_50), .O(gate395inter3));
  inv1  gate901(.a(s_51), .O(gate395inter4));
  nand2 gate902(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate903(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate904(.a(G9), .O(gate395inter7));
  inv1  gate905(.a(G1060), .O(gate395inter8));
  nand2 gate906(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate907(.a(s_51), .b(gate395inter3), .O(gate395inter10));
  nor2  gate908(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate909(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate910(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1079(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1080(.a(gate403inter0), .b(s_76), .O(gate403inter1));
  and2  gate1081(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1082(.a(s_76), .O(gate403inter3));
  inv1  gate1083(.a(s_77), .O(gate403inter4));
  nand2 gate1084(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1085(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1086(.a(G17), .O(gate403inter7));
  inv1  gate1087(.a(G1084), .O(gate403inter8));
  nand2 gate1088(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1089(.a(s_77), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1090(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1091(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1092(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1653(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1654(.a(gate404inter0), .b(s_158), .O(gate404inter1));
  and2  gate1655(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1656(.a(s_158), .O(gate404inter3));
  inv1  gate1657(.a(s_159), .O(gate404inter4));
  nand2 gate1658(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1659(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1660(.a(G18), .O(gate404inter7));
  inv1  gate1661(.a(G1087), .O(gate404inter8));
  nand2 gate1662(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1663(.a(s_159), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1664(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1665(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1666(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate799(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate800(.a(gate409inter0), .b(s_36), .O(gate409inter1));
  and2  gate801(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate802(.a(s_36), .O(gate409inter3));
  inv1  gate803(.a(s_37), .O(gate409inter4));
  nand2 gate804(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate805(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate806(.a(G23), .O(gate409inter7));
  inv1  gate807(.a(G1102), .O(gate409inter8));
  nand2 gate808(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate809(.a(s_37), .b(gate409inter3), .O(gate409inter10));
  nor2  gate810(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate811(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate812(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1485(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1486(.a(gate410inter0), .b(s_134), .O(gate410inter1));
  and2  gate1487(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1488(.a(s_134), .O(gate410inter3));
  inv1  gate1489(.a(s_135), .O(gate410inter4));
  nand2 gate1490(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1491(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1492(.a(G24), .O(gate410inter7));
  inv1  gate1493(.a(G1105), .O(gate410inter8));
  nand2 gate1494(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1495(.a(s_135), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1496(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1497(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1498(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1275(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1276(.a(gate414inter0), .b(s_104), .O(gate414inter1));
  and2  gate1277(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1278(.a(s_104), .O(gate414inter3));
  inv1  gate1279(.a(s_105), .O(gate414inter4));
  nand2 gate1280(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1281(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1282(.a(G28), .O(gate414inter7));
  inv1  gate1283(.a(G1117), .O(gate414inter8));
  nand2 gate1284(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1285(.a(s_105), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1286(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1287(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1288(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1443(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1444(.a(gate417inter0), .b(s_128), .O(gate417inter1));
  and2  gate1445(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1446(.a(s_128), .O(gate417inter3));
  inv1  gate1447(.a(s_129), .O(gate417inter4));
  nand2 gate1448(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1449(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1450(.a(G31), .O(gate417inter7));
  inv1  gate1451(.a(G1126), .O(gate417inter8));
  nand2 gate1452(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1453(.a(s_129), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1454(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1455(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1456(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1261(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1262(.a(gate418inter0), .b(s_102), .O(gate418inter1));
  and2  gate1263(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1264(.a(s_102), .O(gate418inter3));
  inv1  gate1265(.a(s_103), .O(gate418inter4));
  nand2 gate1266(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1267(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1268(.a(G32), .O(gate418inter7));
  inv1  gate1269(.a(G1129), .O(gate418inter8));
  nand2 gate1270(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1271(.a(s_103), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1272(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1273(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1274(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1233(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1234(.a(gate420inter0), .b(s_98), .O(gate420inter1));
  and2  gate1235(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1236(.a(s_98), .O(gate420inter3));
  inv1  gate1237(.a(s_99), .O(gate420inter4));
  nand2 gate1238(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1239(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1240(.a(G1036), .O(gate420inter7));
  inv1  gate1241(.a(G1132), .O(gate420inter8));
  nand2 gate1242(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1243(.a(s_99), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1244(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1245(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1246(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1163(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1164(.a(gate422inter0), .b(s_88), .O(gate422inter1));
  and2  gate1165(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1166(.a(s_88), .O(gate422inter3));
  inv1  gate1167(.a(s_89), .O(gate422inter4));
  nand2 gate1168(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1169(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1170(.a(G1039), .O(gate422inter7));
  inv1  gate1171(.a(G1135), .O(gate422inter8));
  nand2 gate1172(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1173(.a(s_89), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1174(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1175(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1176(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1247(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1248(.a(gate424inter0), .b(s_100), .O(gate424inter1));
  and2  gate1249(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1250(.a(s_100), .O(gate424inter3));
  inv1  gate1251(.a(s_101), .O(gate424inter4));
  nand2 gate1252(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1253(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1254(.a(G1042), .O(gate424inter7));
  inv1  gate1255(.a(G1138), .O(gate424inter8));
  nand2 gate1256(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1257(.a(s_101), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1258(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1259(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1260(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate939(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate940(.a(gate429inter0), .b(s_56), .O(gate429inter1));
  and2  gate941(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate942(.a(s_56), .O(gate429inter3));
  inv1  gate943(.a(s_57), .O(gate429inter4));
  nand2 gate944(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate945(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate946(.a(G6), .O(gate429inter7));
  inv1  gate947(.a(G1147), .O(gate429inter8));
  nand2 gate948(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate949(.a(s_57), .b(gate429inter3), .O(gate429inter10));
  nor2  gate950(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate951(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate952(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1219(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1220(.a(gate430inter0), .b(s_96), .O(gate430inter1));
  and2  gate1221(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1222(.a(s_96), .O(gate430inter3));
  inv1  gate1223(.a(s_97), .O(gate430inter4));
  nand2 gate1224(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1225(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1226(.a(G1051), .O(gate430inter7));
  inv1  gate1227(.a(G1147), .O(gate430inter8));
  nand2 gate1228(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1229(.a(s_97), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1230(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1231(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1232(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1331(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1332(.a(gate435inter0), .b(s_112), .O(gate435inter1));
  and2  gate1333(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1334(.a(s_112), .O(gate435inter3));
  inv1  gate1335(.a(s_113), .O(gate435inter4));
  nand2 gate1336(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1337(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1338(.a(G9), .O(gate435inter7));
  inv1  gate1339(.a(G1156), .O(gate435inter8));
  nand2 gate1340(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1341(.a(s_113), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1342(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1343(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1344(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate687(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate688(.a(gate449inter0), .b(s_20), .O(gate449inter1));
  and2  gate689(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate690(.a(s_20), .O(gate449inter3));
  inv1  gate691(.a(s_21), .O(gate449inter4));
  nand2 gate692(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate693(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate694(.a(G16), .O(gate449inter7));
  inv1  gate695(.a(G1177), .O(gate449inter8));
  nand2 gate696(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate697(.a(s_21), .b(gate449inter3), .O(gate449inter10));
  nor2  gate698(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate699(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate700(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1205(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1206(.a(gate455inter0), .b(s_94), .O(gate455inter1));
  and2  gate1207(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1208(.a(s_94), .O(gate455inter3));
  inv1  gate1209(.a(s_95), .O(gate455inter4));
  nand2 gate1210(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1211(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1212(.a(G19), .O(gate455inter7));
  inv1  gate1213(.a(G1186), .O(gate455inter8));
  nand2 gate1214(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1215(.a(s_95), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1216(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1217(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1218(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate715(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate716(.a(gate463inter0), .b(s_24), .O(gate463inter1));
  and2  gate717(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate718(.a(s_24), .O(gate463inter3));
  inv1  gate719(.a(s_25), .O(gate463inter4));
  nand2 gate720(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate721(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate722(.a(G23), .O(gate463inter7));
  inv1  gate723(.a(G1198), .O(gate463inter8));
  nand2 gate724(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate725(.a(s_25), .b(gate463inter3), .O(gate463inter10));
  nor2  gate726(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate727(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate728(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate771(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate772(.a(gate471inter0), .b(s_32), .O(gate471inter1));
  and2  gate773(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate774(.a(s_32), .O(gate471inter3));
  inv1  gate775(.a(s_33), .O(gate471inter4));
  nand2 gate776(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate777(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate778(.a(G27), .O(gate471inter7));
  inv1  gate779(.a(G1210), .O(gate471inter8));
  nand2 gate780(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate781(.a(s_33), .b(gate471inter3), .O(gate471inter10));
  nor2  gate782(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate783(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate784(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate967(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate968(.a(gate477inter0), .b(s_60), .O(gate477inter1));
  and2  gate969(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate970(.a(s_60), .O(gate477inter3));
  inv1  gate971(.a(s_61), .O(gate477inter4));
  nand2 gate972(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate973(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate974(.a(G30), .O(gate477inter7));
  inv1  gate975(.a(G1219), .O(gate477inter8));
  nand2 gate976(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate977(.a(s_61), .b(gate477inter3), .O(gate477inter10));
  nor2  gate978(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate979(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate980(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1177(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1178(.a(gate479inter0), .b(s_90), .O(gate479inter1));
  and2  gate1179(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1180(.a(s_90), .O(gate479inter3));
  inv1  gate1181(.a(s_91), .O(gate479inter4));
  nand2 gate1182(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1183(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1184(.a(G31), .O(gate479inter7));
  inv1  gate1185(.a(G1222), .O(gate479inter8));
  nand2 gate1186(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1187(.a(s_91), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1188(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1189(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1190(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate827(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate828(.a(gate486inter0), .b(s_40), .O(gate486inter1));
  and2  gate829(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate830(.a(s_40), .O(gate486inter3));
  inv1  gate831(.a(s_41), .O(gate486inter4));
  nand2 gate832(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate833(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate834(.a(G1234), .O(gate486inter7));
  inv1  gate835(.a(G1235), .O(gate486inter8));
  nand2 gate836(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate837(.a(s_41), .b(gate486inter3), .O(gate486inter10));
  nor2  gate838(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate839(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate840(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1625(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1626(.a(gate492inter0), .b(s_154), .O(gate492inter1));
  and2  gate1627(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1628(.a(s_154), .O(gate492inter3));
  inv1  gate1629(.a(s_155), .O(gate492inter4));
  nand2 gate1630(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1631(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1632(.a(G1246), .O(gate492inter7));
  inv1  gate1633(.a(G1247), .O(gate492inter8));
  nand2 gate1634(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1635(.a(s_155), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1636(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1637(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1638(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1149(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1150(.a(gate497inter0), .b(s_86), .O(gate497inter1));
  and2  gate1151(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1152(.a(s_86), .O(gate497inter3));
  inv1  gate1153(.a(s_87), .O(gate497inter4));
  nand2 gate1154(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1155(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1156(.a(G1256), .O(gate497inter7));
  inv1  gate1157(.a(G1257), .O(gate497inter8));
  nand2 gate1158(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1159(.a(s_87), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1160(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1161(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1162(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1289(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1290(.a(gate504inter0), .b(s_106), .O(gate504inter1));
  and2  gate1291(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1292(.a(s_106), .O(gate504inter3));
  inv1  gate1293(.a(s_107), .O(gate504inter4));
  nand2 gate1294(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1295(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1296(.a(G1270), .O(gate504inter7));
  inv1  gate1297(.a(G1271), .O(gate504inter8));
  nand2 gate1298(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1299(.a(s_107), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1300(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1301(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1302(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1373(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1374(.a(gate514inter0), .b(s_118), .O(gate514inter1));
  and2  gate1375(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1376(.a(s_118), .O(gate514inter3));
  inv1  gate1377(.a(s_119), .O(gate514inter4));
  nand2 gate1378(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1379(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1380(.a(G1290), .O(gate514inter7));
  inv1  gate1381(.a(G1291), .O(gate514inter8));
  nand2 gate1382(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1383(.a(s_119), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1384(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1385(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1386(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule