module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1191(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1192(.a(gate16inter0), .b(s_92), .O(gate16inter1));
  and2  gate1193(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1194(.a(s_92), .O(gate16inter3));
  inv1  gate1195(.a(s_93), .O(gate16inter4));
  nand2 gate1196(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1197(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1198(.a(G15), .O(gate16inter7));
  inv1  gate1199(.a(G16), .O(gate16inter8));
  nand2 gate1200(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1201(.a(s_93), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1202(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1203(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1204(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1177(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1178(.a(gate20inter0), .b(s_90), .O(gate20inter1));
  and2  gate1179(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1180(.a(s_90), .O(gate20inter3));
  inv1  gate1181(.a(s_91), .O(gate20inter4));
  nand2 gate1182(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1183(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1184(.a(G23), .O(gate20inter7));
  inv1  gate1185(.a(G24), .O(gate20inter8));
  nand2 gate1186(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1187(.a(s_91), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1188(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1189(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1190(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1149(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1150(.a(gate26inter0), .b(s_86), .O(gate26inter1));
  and2  gate1151(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1152(.a(s_86), .O(gate26inter3));
  inv1  gate1153(.a(s_87), .O(gate26inter4));
  nand2 gate1154(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1155(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1156(.a(G9), .O(gate26inter7));
  inv1  gate1157(.a(G13), .O(gate26inter8));
  nand2 gate1158(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1159(.a(s_87), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1160(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1161(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1162(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1373(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1374(.a(gate33inter0), .b(s_118), .O(gate33inter1));
  and2  gate1375(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1376(.a(s_118), .O(gate33inter3));
  inv1  gate1377(.a(s_119), .O(gate33inter4));
  nand2 gate1378(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1379(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1380(.a(G17), .O(gate33inter7));
  inv1  gate1381(.a(G21), .O(gate33inter8));
  nand2 gate1382(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1383(.a(s_119), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1384(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1385(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1386(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate827(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate828(.a(gate39inter0), .b(s_40), .O(gate39inter1));
  and2  gate829(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate830(.a(s_40), .O(gate39inter3));
  inv1  gate831(.a(s_41), .O(gate39inter4));
  nand2 gate832(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate833(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate834(.a(G20), .O(gate39inter7));
  inv1  gate835(.a(G24), .O(gate39inter8));
  nand2 gate836(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate837(.a(s_41), .b(gate39inter3), .O(gate39inter10));
  nor2  gate838(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate839(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate840(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate771(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate772(.a(gate45inter0), .b(s_32), .O(gate45inter1));
  and2  gate773(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate774(.a(s_32), .O(gate45inter3));
  inv1  gate775(.a(s_33), .O(gate45inter4));
  nand2 gate776(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate777(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate778(.a(G5), .O(gate45inter7));
  inv1  gate779(.a(G272), .O(gate45inter8));
  nand2 gate780(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate781(.a(s_33), .b(gate45inter3), .O(gate45inter10));
  nor2  gate782(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate783(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate784(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1079(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1080(.a(gate52inter0), .b(s_76), .O(gate52inter1));
  and2  gate1081(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1082(.a(s_76), .O(gate52inter3));
  inv1  gate1083(.a(s_77), .O(gate52inter4));
  nand2 gate1084(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1085(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1086(.a(G12), .O(gate52inter7));
  inv1  gate1087(.a(G281), .O(gate52inter8));
  nand2 gate1088(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1089(.a(s_77), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1090(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1091(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1092(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1289(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1290(.a(gate54inter0), .b(s_106), .O(gate54inter1));
  and2  gate1291(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1292(.a(s_106), .O(gate54inter3));
  inv1  gate1293(.a(s_107), .O(gate54inter4));
  nand2 gate1294(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1295(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1296(.a(G14), .O(gate54inter7));
  inv1  gate1297(.a(G284), .O(gate54inter8));
  nand2 gate1298(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1299(.a(s_107), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1300(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1301(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1302(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1205(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1206(.a(gate58inter0), .b(s_94), .O(gate58inter1));
  and2  gate1207(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1208(.a(s_94), .O(gate58inter3));
  inv1  gate1209(.a(s_95), .O(gate58inter4));
  nand2 gate1210(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1211(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1212(.a(G18), .O(gate58inter7));
  inv1  gate1213(.a(G290), .O(gate58inter8));
  nand2 gate1214(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1215(.a(s_95), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1216(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1217(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1218(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1443(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1444(.a(gate63inter0), .b(s_128), .O(gate63inter1));
  and2  gate1445(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1446(.a(s_128), .O(gate63inter3));
  inv1  gate1447(.a(s_129), .O(gate63inter4));
  nand2 gate1448(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1449(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1450(.a(G23), .O(gate63inter7));
  inv1  gate1451(.a(G299), .O(gate63inter8));
  nand2 gate1452(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1453(.a(s_129), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1454(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1455(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1456(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate715(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate716(.a(gate66inter0), .b(s_24), .O(gate66inter1));
  and2  gate717(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate718(.a(s_24), .O(gate66inter3));
  inv1  gate719(.a(s_25), .O(gate66inter4));
  nand2 gate720(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate721(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate722(.a(G26), .O(gate66inter7));
  inv1  gate723(.a(G302), .O(gate66inter8));
  nand2 gate724(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate725(.a(s_25), .b(gate66inter3), .O(gate66inter10));
  nor2  gate726(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate727(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate728(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1051(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1052(.a(gate90inter0), .b(s_72), .O(gate90inter1));
  and2  gate1053(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1054(.a(s_72), .O(gate90inter3));
  inv1  gate1055(.a(s_73), .O(gate90inter4));
  nand2 gate1056(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1057(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1058(.a(G21), .O(gate90inter7));
  inv1  gate1059(.a(G338), .O(gate90inter8));
  nand2 gate1060(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1061(.a(s_73), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1062(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1063(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1064(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate729(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate730(.a(gate99inter0), .b(s_26), .O(gate99inter1));
  and2  gate731(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate732(.a(s_26), .O(gate99inter3));
  inv1  gate733(.a(s_27), .O(gate99inter4));
  nand2 gate734(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate735(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate736(.a(G27), .O(gate99inter7));
  inv1  gate737(.a(G353), .O(gate99inter8));
  nand2 gate738(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate739(.a(s_27), .b(gate99inter3), .O(gate99inter10));
  nor2  gate740(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate741(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate742(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1499(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1500(.a(gate100inter0), .b(s_136), .O(gate100inter1));
  and2  gate1501(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1502(.a(s_136), .O(gate100inter3));
  inv1  gate1503(.a(s_137), .O(gate100inter4));
  nand2 gate1504(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1505(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1506(.a(G31), .O(gate100inter7));
  inv1  gate1507(.a(G353), .O(gate100inter8));
  nand2 gate1508(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1509(.a(s_137), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1510(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1511(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1512(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1387(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1388(.a(gate103inter0), .b(s_120), .O(gate103inter1));
  and2  gate1389(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1390(.a(s_120), .O(gate103inter3));
  inv1  gate1391(.a(s_121), .O(gate103inter4));
  nand2 gate1392(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1393(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1394(.a(G28), .O(gate103inter7));
  inv1  gate1395(.a(G359), .O(gate103inter8));
  nand2 gate1396(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1397(.a(s_121), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1398(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1399(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1400(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate603(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate604(.a(gate110inter0), .b(s_8), .O(gate110inter1));
  and2  gate605(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate606(.a(s_8), .O(gate110inter3));
  inv1  gate607(.a(s_9), .O(gate110inter4));
  nand2 gate608(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate609(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate610(.a(G372), .O(gate110inter7));
  inv1  gate611(.a(G373), .O(gate110inter8));
  nand2 gate612(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate613(.a(s_9), .b(gate110inter3), .O(gate110inter10));
  nor2  gate614(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate615(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate616(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1135(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1136(.a(gate117inter0), .b(s_84), .O(gate117inter1));
  and2  gate1137(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1138(.a(s_84), .O(gate117inter3));
  inv1  gate1139(.a(s_85), .O(gate117inter4));
  nand2 gate1140(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1141(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1142(.a(G386), .O(gate117inter7));
  inv1  gate1143(.a(G387), .O(gate117inter8));
  nand2 gate1144(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1145(.a(s_85), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1146(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1147(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1148(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate995(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate996(.a(gate122inter0), .b(s_64), .O(gate122inter1));
  and2  gate997(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate998(.a(s_64), .O(gate122inter3));
  inv1  gate999(.a(s_65), .O(gate122inter4));
  nand2 gate1000(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1001(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1002(.a(G396), .O(gate122inter7));
  inv1  gate1003(.a(G397), .O(gate122inter8));
  nand2 gate1004(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1005(.a(s_65), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1006(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1007(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1008(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate799(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate800(.a(gate124inter0), .b(s_36), .O(gate124inter1));
  and2  gate801(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate802(.a(s_36), .O(gate124inter3));
  inv1  gate803(.a(s_37), .O(gate124inter4));
  nand2 gate804(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate805(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate806(.a(G400), .O(gate124inter7));
  inv1  gate807(.a(G401), .O(gate124inter8));
  nand2 gate808(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate809(.a(s_37), .b(gate124inter3), .O(gate124inter10));
  nor2  gate810(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate811(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate812(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1121(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1122(.a(gate130inter0), .b(s_82), .O(gate130inter1));
  and2  gate1123(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1124(.a(s_82), .O(gate130inter3));
  inv1  gate1125(.a(s_83), .O(gate130inter4));
  nand2 gate1126(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1127(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1128(.a(G412), .O(gate130inter7));
  inv1  gate1129(.a(G413), .O(gate130inter8));
  nand2 gate1130(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1131(.a(s_83), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1132(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1133(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1134(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1163(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1164(.a(gate133inter0), .b(s_88), .O(gate133inter1));
  and2  gate1165(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1166(.a(s_88), .O(gate133inter3));
  inv1  gate1167(.a(s_89), .O(gate133inter4));
  nand2 gate1168(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1169(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1170(.a(G418), .O(gate133inter7));
  inv1  gate1171(.a(G419), .O(gate133inter8));
  nand2 gate1172(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1173(.a(s_89), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1174(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1175(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1176(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate701(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate702(.a(gate141inter0), .b(s_22), .O(gate141inter1));
  and2  gate703(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate704(.a(s_22), .O(gate141inter3));
  inv1  gate705(.a(s_23), .O(gate141inter4));
  nand2 gate706(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate707(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate708(.a(G450), .O(gate141inter7));
  inv1  gate709(.a(G453), .O(gate141inter8));
  nand2 gate710(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate711(.a(s_23), .b(gate141inter3), .O(gate141inter10));
  nor2  gate712(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate713(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate714(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate547(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate548(.a(gate148inter0), .b(s_0), .O(gate148inter1));
  and2  gate549(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate550(.a(s_0), .O(gate148inter3));
  inv1  gate551(.a(s_1), .O(gate148inter4));
  nand2 gate552(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate553(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate554(.a(G492), .O(gate148inter7));
  inv1  gate555(.a(G495), .O(gate148inter8));
  nand2 gate556(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate557(.a(s_1), .b(gate148inter3), .O(gate148inter10));
  nor2  gate558(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate559(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate560(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1219(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1220(.a(gate151inter0), .b(s_96), .O(gate151inter1));
  and2  gate1221(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1222(.a(s_96), .O(gate151inter3));
  inv1  gate1223(.a(s_97), .O(gate151inter4));
  nand2 gate1224(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1225(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1226(.a(G510), .O(gate151inter7));
  inv1  gate1227(.a(G513), .O(gate151inter8));
  nand2 gate1228(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1229(.a(s_97), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1230(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1231(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1232(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1401(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1402(.a(gate155inter0), .b(s_122), .O(gate155inter1));
  and2  gate1403(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1404(.a(s_122), .O(gate155inter3));
  inv1  gate1405(.a(s_123), .O(gate155inter4));
  nand2 gate1406(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1407(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1408(.a(G432), .O(gate155inter7));
  inv1  gate1409(.a(G525), .O(gate155inter8));
  nand2 gate1410(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1411(.a(s_123), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1412(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1413(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1414(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate617(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate618(.a(gate158inter0), .b(s_10), .O(gate158inter1));
  and2  gate619(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate620(.a(s_10), .O(gate158inter3));
  inv1  gate621(.a(s_11), .O(gate158inter4));
  nand2 gate622(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate623(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate624(.a(G441), .O(gate158inter7));
  inv1  gate625(.a(G528), .O(gate158inter8));
  nand2 gate626(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate627(.a(s_11), .b(gate158inter3), .O(gate158inter10));
  nor2  gate628(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate629(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate630(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1485(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1486(.a(gate168inter0), .b(s_134), .O(gate168inter1));
  and2  gate1487(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1488(.a(s_134), .O(gate168inter3));
  inv1  gate1489(.a(s_135), .O(gate168inter4));
  nand2 gate1490(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1491(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1492(.a(G471), .O(gate168inter7));
  inv1  gate1493(.a(G543), .O(gate168inter8));
  nand2 gate1494(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1495(.a(s_135), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1496(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1497(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1498(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate897(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate898(.a(gate185inter0), .b(s_50), .O(gate185inter1));
  and2  gate899(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate900(.a(s_50), .O(gate185inter3));
  inv1  gate901(.a(s_51), .O(gate185inter4));
  nand2 gate902(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate903(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate904(.a(G570), .O(gate185inter7));
  inv1  gate905(.a(G571), .O(gate185inter8));
  nand2 gate906(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate907(.a(s_51), .b(gate185inter3), .O(gate185inter10));
  nor2  gate908(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate909(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate910(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1303(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1304(.a(gate190inter0), .b(s_108), .O(gate190inter1));
  and2  gate1305(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1306(.a(s_108), .O(gate190inter3));
  inv1  gate1307(.a(s_109), .O(gate190inter4));
  nand2 gate1308(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1309(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1310(.a(G580), .O(gate190inter7));
  inv1  gate1311(.a(G581), .O(gate190inter8));
  nand2 gate1312(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1313(.a(s_109), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1314(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1315(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1316(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate561(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate562(.a(gate198inter0), .b(s_2), .O(gate198inter1));
  and2  gate563(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate564(.a(s_2), .O(gate198inter3));
  inv1  gate565(.a(s_3), .O(gate198inter4));
  nand2 gate566(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate567(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate568(.a(G596), .O(gate198inter7));
  inv1  gate569(.a(G597), .O(gate198inter8));
  nand2 gate570(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate571(.a(s_3), .b(gate198inter3), .O(gate198inter10));
  nor2  gate572(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate573(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate574(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1345(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1346(.a(gate199inter0), .b(s_114), .O(gate199inter1));
  and2  gate1347(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1348(.a(s_114), .O(gate199inter3));
  inv1  gate1349(.a(s_115), .O(gate199inter4));
  nand2 gate1350(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1351(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1352(.a(G598), .O(gate199inter7));
  inv1  gate1353(.a(G599), .O(gate199inter8));
  nand2 gate1354(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1355(.a(s_115), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1356(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1357(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1358(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate575(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate576(.a(gate201inter0), .b(s_4), .O(gate201inter1));
  and2  gate577(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate578(.a(s_4), .O(gate201inter3));
  inv1  gate579(.a(s_5), .O(gate201inter4));
  nand2 gate580(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate581(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate582(.a(G602), .O(gate201inter7));
  inv1  gate583(.a(G607), .O(gate201inter8));
  nand2 gate584(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate585(.a(s_5), .b(gate201inter3), .O(gate201inter10));
  nor2  gate586(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate587(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate588(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1513(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1514(.a(gate208inter0), .b(s_138), .O(gate208inter1));
  and2  gate1515(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1516(.a(s_138), .O(gate208inter3));
  inv1  gate1517(.a(s_139), .O(gate208inter4));
  nand2 gate1518(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1519(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1520(.a(G627), .O(gate208inter7));
  inv1  gate1521(.a(G637), .O(gate208inter8));
  nand2 gate1522(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1523(.a(s_139), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1524(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1525(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1526(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate869(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate870(.a(gate228inter0), .b(s_46), .O(gate228inter1));
  and2  gate871(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate872(.a(s_46), .O(gate228inter3));
  inv1  gate873(.a(s_47), .O(gate228inter4));
  nand2 gate874(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate875(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate876(.a(G696), .O(gate228inter7));
  inv1  gate877(.a(G697), .O(gate228inter8));
  nand2 gate878(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate879(.a(s_47), .b(gate228inter3), .O(gate228inter10));
  nor2  gate880(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate881(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate882(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate673(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate674(.a(gate231inter0), .b(s_18), .O(gate231inter1));
  and2  gate675(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate676(.a(s_18), .O(gate231inter3));
  inv1  gate677(.a(s_19), .O(gate231inter4));
  nand2 gate678(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate679(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate680(.a(G702), .O(gate231inter7));
  inv1  gate681(.a(G703), .O(gate231inter8));
  nand2 gate682(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate683(.a(s_19), .b(gate231inter3), .O(gate231inter10));
  nor2  gate684(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate685(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate686(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1093(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1094(.a(gate236inter0), .b(s_78), .O(gate236inter1));
  and2  gate1095(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1096(.a(s_78), .O(gate236inter3));
  inv1  gate1097(.a(s_79), .O(gate236inter4));
  nand2 gate1098(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1099(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1100(.a(G251), .O(gate236inter7));
  inv1  gate1101(.a(G727), .O(gate236inter8));
  nand2 gate1102(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1103(.a(s_79), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1104(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1105(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1106(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate981(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate982(.a(gate247inter0), .b(s_62), .O(gate247inter1));
  and2  gate983(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate984(.a(s_62), .O(gate247inter3));
  inv1  gate985(.a(s_63), .O(gate247inter4));
  nand2 gate986(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate987(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate988(.a(G251), .O(gate247inter7));
  inv1  gate989(.a(G739), .O(gate247inter8));
  nand2 gate990(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate991(.a(s_63), .b(gate247inter3), .O(gate247inter10));
  nor2  gate992(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate993(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate994(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate883(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate884(.a(gate252inter0), .b(s_48), .O(gate252inter1));
  and2  gate885(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate886(.a(s_48), .O(gate252inter3));
  inv1  gate887(.a(s_49), .O(gate252inter4));
  nand2 gate888(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate889(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate890(.a(G709), .O(gate252inter7));
  inv1  gate891(.a(G745), .O(gate252inter8));
  nand2 gate892(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate893(.a(s_49), .b(gate252inter3), .O(gate252inter10));
  nor2  gate894(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate895(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate896(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate631(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate632(.a(gate255inter0), .b(s_12), .O(gate255inter1));
  and2  gate633(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate634(.a(s_12), .O(gate255inter3));
  inv1  gate635(.a(s_13), .O(gate255inter4));
  nand2 gate636(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate637(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate638(.a(G263), .O(gate255inter7));
  inv1  gate639(.a(G751), .O(gate255inter8));
  nand2 gate640(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate641(.a(s_13), .b(gate255inter3), .O(gate255inter10));
  nor2  gate642(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate643(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate644(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate785(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate786(.a(gate263inter0), .b(s_34), .O(gate263inter1));
  and2  gate787(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate788(.a(s_34), .O(gate263inter3));
  inv1  gate789(.a(s_35), .O(gate263inter4));
  nand2 gate790(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate791(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate792(.a(G766), .O(gate263inter7));
  inv1  gate793(.a(G767), .O(gate263inter8));
  nand2 gate794(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate795(.a(s_35), .b(gate263inter3), .O(gate263inter10));
  nor2  gate796(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate797(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate798(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1317(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1318(.a(gate267inter0), .b(s_110), .O(gate267inter1));
  and2  gate1319(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1320(.a(s_110), .O(gate267inter3));
  inv1  gate1321(.a(s_111), .O(gate267inter4));
  nand2 gate1322(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1323(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1324(.a(G648), .O(gate267inter7));
  inv1  gate1325(.a(G776), .O(gate267inter8));
  nand2 gate1326(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1327(.a(s_111), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1328(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1329(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1330(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1359(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1360(.a(gate269inter0), .b(s_116), .O(gate269inter1));
  and2  gate1361(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1362(.a(s_116), .O(gate269inter3));
  inv1  gate1363(.a(s_117), .O(gate269inter4));
  nand2 gate1364(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1365(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1366(.a(G654), .O(gate269inter7));
  inv1  gate1367(.a(G782), .O(gate269inter8));
  nand2 gate1368(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1369(.a(s_117), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1370(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1371(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1372(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate813(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate814(.a(gate270inter0), .b(s_38), .O(gate270inter1));
  and2  gate815(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate816(.a(s_38), .O(gate270inter3));
  inv1  gate817(.a(s_39), .O(gate270inter4));
  nand2 gate818(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate819(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate820(.a(G657), .O(gate270inter7));
  inv1  gate821(.a(G785), .O(gate270inter8));
  nand2 gate822(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate823(.a(s_39), .b(gate270inter3), .O(gate270inter10));
  nor2  gate824(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate825(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate826(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1247(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1248(.a(gate290inter0), .b(s_100), .O(gate290inter1));
  and2  gate1249(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1250(.a(s_100), .O(gate290inter3));
  inv1  gate1251(.a(s_101), .O(gate290inter4));
  nand2 gate1252(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1253(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1254(.a(G820), .O(gate290inter7));
  inv1  gate1255(.a(G821), .O(gate290inter8));
  nand2 gate1256(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1257(.a(s_101), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1258(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1259(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1260(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate855(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate856(.a(gate292inter0), .b(s_44), .O(gate292inter1));
  and2  gate857(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate858(.a(s_44), .O(gate292inter3));
  inv1  gate859(.a(s_45), .O(gate292inter4));
  nand2 gate860(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate861(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate862(.a(G824), .O(gate292inter7));
  inv1  gate863(.a(G825), .O(gate292inter8));
  nand2 gate864(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate865(.a(s_45), .b(gate292inter3), .O(gate292inter10));
  nor2  gate866(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate867(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate868(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate939(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate940(.a(gate293inter0), .b(s_56), .O(gate293inter1));
  and2  gate941(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate942(.a(s_56), .O(gate293inter3));
  inv1  gate943(.a(s_57), .O(gate293inter4));
  nand2 gate944(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate945(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate946(.a(G828), .O(gate293inter7));
  inv1  gate947(.a(G829), .O(gate293inter8));
  nand2 gate948(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate949(.a(s_57), .b(gate293inter3), .O(gate293inter10));
  nor2  gate950(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate951(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate952(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1037(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1038(.a(gate294inter0), .b(s_70), .O(gate294inter1));
  and2  gate1039(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1040(.a(s_70), .O(gate294inter3));
  inv1  gate1041(.a(s_71), .O(gate294inter4));
  nand2 gate1042(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1043(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1044(.a(G832), .O(gate294inter7));
  inv1  gate1045(.a(G833), .O(gate294inter8));
  nand2 gate1046(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1047(.a(s_71), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1048(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1049(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1050(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate743(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate744(.a(gate393inter0), .b(s_28), .O(gate393inter1));
  and2  gate745(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate746(.a(s_28), .O(gate393inter3));
  inv1  gate747(.a(s_29), .O(gate393inter4));
  nand2 gate748(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate749(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate750(.a(G7), .O(gate393inter7));
  inv1  gate751(.a(G1054), .O(gate393inter8));
  nand2 gate752(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate753(.a(s_29), .b(gate393inter3), .O(gate393inter10));
  nor2  gate754(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate755(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate756(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1009(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1010(.a(gate398inter0), .b(s_66), .O(gate398inter1));
  and2  gate1011(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1012(.a(s_66), .O(gate398inter3));
  inv1  gate1013(.a(s_67), .O(gate398inter4));
  nand2 gate1014(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1015(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1016(.a(G12), .O(gate398inter7));
  inv1  gate1017(.a(G1069), .O(gate398inter8));
  nand2 gate1018(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1019(.a(s_67), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1020(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1021(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1022(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1415(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1416(.a(gate399inter0), .b(s_124), .O(gate399inter1));
  and2  gate1417(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1418(.a(s_124), .O(gate399inter3));
  inv1  gate1419(.a(s_125), .O(gate399inter4));
  nand2 gate1420(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1421(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1422(.a(G13), .O(gate399inter7));
  inv1  gate1423(.a(G1072), .O(gate399inter8));
  nand2 gate1424(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1425(.a(s_125), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1426(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1427(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1428(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1233(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1234(.a(gate419inter0), .b(s_98), .O(gate419inter1));
  and2  gate1235(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1236(.a(s_98), .O(gate419inter3));
  inv1  gate1237(.a(s_99), .O(gate419inter4));
  nand2 gate1238(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1239(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1240(.a(G1), .O(gate419inter7));
  inv1  gate1241(.a(G1132), .O(gate419inter8));
  nand2 gate1242(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1243(.a(s_99), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1244(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1245(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1246(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate757(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate758(.a(gate422inter0), .b(s_30), .O(gate422inter1));
  and2  gate759(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate760(.a(s_30), .O(gate422inter3));
  inv1  gate761(.a(s_31), .O(gate422inter4));
  nand2 gate762(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate763(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate764(.a(G1039), .O(gate422inter7));
  inv1  gate765(.a(G1135), .O(gate422inter8));
  nand2 gate766(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate767(.a(s_31), .b(gate422inter3), .O(gate422inter10));
  nor2  gate768(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate769(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate770(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1331(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1332(.a(gate433inter0), .b(s_112), .O(gate433inter1));
  and2  gate1333(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1334(.a(s_112), .O(gate433inter3));
  inv1  gate1335(.a(s_113), .O(gate433inter4));
  nand2 gate1336(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1337(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1338(.a(G8), .O(gate433inter7));
  inv1  gate1339(.a(G1153), .O(gate433inter8));
  nand2 gate1340(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1341(.a(s_113), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1342(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1343(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1344(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1023(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1024(.a(gate438inter0), .b(s_68), .O(gate438inter1));
  and2  gate1025(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1026(.a(s_68), .O(gate438inter3));
  inv1  gate1027(.a(s_69), .O(gate438inter4));
  nand2 gate1028(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1029(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1030(.a(G1063), .O(gate438inter7));
  inv1  gate1031(.a(G1159), .O(gate438inter8));
  nand2 gate1032(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1033(.a(s_69), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1034(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1035(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1036(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate911(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate912(.a(gate447inter0), .b(s_52), .O(gate447inter1));
  and2  gate913(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate914(.a(s_52), .O(gate447inter3));
  inv1  gate915(.a(s_53), .O(gate447inter4));
  nand2 gate916(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate917(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate918(.a(G15), .O(gate447inter7));
  inv1  gate919(.a(G1174), .O(gate447inter8));
  nand2 gate920(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate921(.a(s_53), .b(gate447inter3), .O(gate447inter10));
  nor2  gate922(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate923(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate924(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1065(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1066(.a(gate459inter0), .b(s_74), .O(gate459inter1));
  and2  gate1067(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1068(.a(s_74), .O(gate459inter3));
  inv1  gate1069(.a(s_75), .O(gate459inter4));
  nand2 gate1070(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1071(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1072(.a(G21), .O(gate459inter7));
  inv1  gate1073(.a(G1192), .O(gate459inter8));
  nand2 gate1074(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1075(.a(s_75), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1076(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1077(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1078(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1275(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1276(.a(gate465inter0), .b(s_104), .O(gate465inter1));
  and2  gate1277(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1278(.a(s_104), .O(gate465inter3));
  inv1  gate1279(.a(s_105), .O(gate465inter4));
  nand2 gate1280(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1281(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1282(.a(G24), .O(gate465inter7));
  inv1  gate1283(.a(G1201), .O(gate465inter8));
  nand2 gate1284(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1285(.a(s_105), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1286(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1287(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1288(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1527(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1528(.a(gate467inter0), .b(s_140), .O(gate467inter1));
  and2  gate1529(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1530(.a(s_140), .O(gate467inter3));
  inv1  gate1531(.a(s_141), .O(gate467inter4));
  nand2 gate1532(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1533(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1534(.a(G25), .O(gate467inter7));
  inv1  gate1535(.a(G1204), .O(gate467inter8));
  nand2 gate1536(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1537(.a(s_141), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1538(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1539(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1540(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate841(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate842(.a(gate470inter0), .b(s_42), .O(gate470inter1));
  and2  gate843(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate844(.a(s_42), .O(gate470inter3));
  inv1  gate845(.a(s_43), .O(gate470inter4));
  nand2 gate846(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate847(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate848(.a(G1111), .O(gate470inter7));
  inv1  gate849(.a(G1207), .O(gate470inter8));
  nand2 gate850(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate851(.a(s_43), .b(gate470inter3), .O(gate470inter10));
  nor2  gate852(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate853(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate854(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1457(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1458(.a(gate472inter0), .b(s_130), .O(gate472inter1));
  and2  gate1459(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1460(.a(s_130), .O(gate472inter3));
  inv1  gate1461(.a(s_131), .O(gate472inter4));
  nand2 gate1462(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1463(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1464(.a(G1114), .O(gate472inter7));
  inv1  gate1465(.a(G1210), .O(gate472inter8));
  nand2 gate1466(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1467(.a(s_131), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1468(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1469(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1470(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate953(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate954(.a(gate473inter0), .b(s_58), .O(gate473inter1));
  and2  gate955(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate956(.a(s_58), .O(gate473inter3));
  inv1  gate957(.a(s_59), .O(gate473inter4));
  nand2 gate958(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate959(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate960(.a(G28), .O(gate473inter7));
  inv1  gate961(.a(G1213), .O(gate473inter8));
  nand2 gate962(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate963(.a(s_59), .b(gate473inter3), .O(gate473inter10));
  nor2  gate964(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate965(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate966(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate589(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate590(.a(gate475inter0), .b(s_6), .O(gate475inter1));
  and2  gate591(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate592(.a(s_6), .O(gate475inter3));
  inv1  gate593(.a(s_7), .O(gate475inter4));
  nand2 gate594(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate595(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate596(.a(G29), .O(gate475inter7));
  inv1  gate597(.a(G1216), .O(gate475inter8));
  nand2 gate598(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate599(.a(s_7), .b(gate475inter3), .O(gate475inter10));
  nor2  gate600(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate601(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate602(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate687(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate688(.a(gate485inter0), .b(s_20), .O(gate485inter1));
  and2  gate689(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate690(.a(s_20), .O(gate485inter3));
  inv1  gate691(.a(s_21), .O(gate485inter4));
  nand2 gate692(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate693(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate694(.a(G1232), .O(gate485inter7));
  inv1  gate695(.a(G1233), .O(gate485inter8));
  nand2 gate696(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate697(.a(s_21), .b(gate485inter3), .O(gate485inter10));
  nor2  gate698(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate699(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate700(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1429(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1430(.a(gate489inter0), .b(s_126), .O(gate489inter1));
  and2  gate1431(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1432(.a(s_126), .O(gate489inter3));
  inv1  gate1433(.a(s_127), .O(gate489inter4));
  nand2 gate1434(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1435(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1436(.a(G1240), .O(gate489inter7));
  inv1  gate1437(.a(G1241), .O(gate489inter8));
  nand2 gate1438(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1439(.a(s_127), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1440(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1441(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1442(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1261(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1262(.a(gate491inter0), .b(s_102), .O(gate491inter1));
  and2  gate1263(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1264(.a(s_102), .O(gate491inter3));
  inv1  gate1265(.a(s_103), .O(gate491inter4));
  nand2 gate1266(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1267(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1268(.a(G1244), .O(gate491inter7));
  inv1  gate1269(.a(G1245), .O(gate491inter8));
  nand2 gate1270(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1271(.a(s_103), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1272(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1273(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1274(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate645(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate646(.a(gate492inter0), .b(s_14), .O(gate492inter1));
  and2  gate647(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate648(.a(s_14), .O(gate492inter3));
  inv1  gate649(.a(s_15), .O(gate492inter4));
  nand2 gate650(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate651(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate652(.a(G1246), .O(gate492inter7));
  inv1  gate653(.a(G1247), .O(gate492inter8));
  nand2 gate654(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate655(.a(s_15), .b(gate492inter3), .O(gate492inter10));
  nor2  gate656(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate657(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate658(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1471(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1472(.a(gate493inter0), .b(s_132), .O(gate493inter1));
  and2  gate1473(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1474(.a(s_132), .O(gate493inter3));
  inv1  gate1475(.a(s_133), .O(gate493inter4));
  nand2 gate1476(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1477(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1478(.a(G1248), .O(gate493inter7));
  inv1  gate1479(.a(G1249), .O(gate493inter8));
  nand2 gate1480(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1481(.a(s_133), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1482(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1483(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1484(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate967(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate968(.a(gate500inter0), .b(s_60), .O(gate500inter1));
  and2  gate969(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate970(.a(s_60), .O(gate500inter3));
  inv1  gate971(.a(s_61), .O(gate500inter4));
  nand2 gate972(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate973(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate974(.a(G1262), .O(gate500inter7));
  inv1  gate975(.a(G1263), .O(gate500inter8));
  nand2 gate976(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate977(.a(s_61), .b(gate500inter3), .O(gate500inter10));
  nor2  gate978(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate979(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate980(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate925(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate926(.a(gate502inter0), .b(s_54), .O(gate502inter1));
  and2  gate927(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate928(.a(s_54), .O(gate502inter3));
  inv1  gate929(.a(s_55), .O(gate502inter4));
  nand2 gate930(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate931(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate932(.a(G1266), .O(gate502inter7));
  inv1  gate933(.a(G1267), .O(gate502inter8));
  nand2 gate934(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate935(.a(s_55), .b(gate502inter3), .O(gate502inter10));
  nor2  gate936(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate937(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate938(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1107(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1108(.a(gate509inter0), .b(s_80), .O(gate509inter1));
  and2  gate1109(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1110(.a(s_80), .O(gate509inter3));
  inv1  gate1111(.a(s_81), .O(gate509inter4));
  nand2 gate1112(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1113(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1114(.a(G1280), .O(gate509inter7));
  inv1  gate1115(.a(G1281), .O(gate509inter8));
  nand2 gate1116(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1117(.a(s_81), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1118(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1119(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1120(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate659(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate660(.a(gate511inter0), .b(s_16), .O(gate511inter1));
  and2  gate661(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate662(.a(s_16), .O(gate511inter3));
  inv1  gate663(.a(s_17), .O(gate511inter4));
  nand2 gate664(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate665(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate666(.a(G1284), .O(gate511inter7));
  inv1  gate667(.a(G1285), .O(gate511inter8));
  nand2 gate668(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate669(.a(s_17), .b(gate511inter3), .O(gate511inter10));
  nor2  gate670(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate671(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate672(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule