module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2479(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2480(.a(gate10inter0), .b(s_276), .O(gate10inter1));
  and2  gate2481(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2482(.a(s_276), .O(gate10inter3));
  inv1  gate2483(.a(s_277), .O(gate10inter4));
  nand2 gate2484(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2485(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2486(.a(G3), .O(gate10inter7));
  inv1  gate2487(.a(G4), .O(gate10inter8));
  nand2 gate2488(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2489(.a(s_277), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2490(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2491(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2492(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate659(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate660(.a(gate12inter0), .b(s_16), .O(gate12inter1));
  and2  gate661(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate662(.a(s_16), .O(gate12inter3));
  inv1  gate663(.a(s_17), .O(gate12inter4));
  nand2 gate664(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate665(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate666(.a(G7), .O(gate12inter7));
  inv1  gate667(.a(G8), .O(gate12inter8));
  nand2 gate668(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate669(.a(s_17), .b(gate12inter3), .O(gate12inter10));
  nor2  gate670(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate671(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate672(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2703(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2704(.a(gate13inter0), .b(s_308), .O(gate13inter1));
  and2  gate2705(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2706(.a(s_308), .O(gate13inter3));
  inv1  gate2707(.a(s_309), .O(gate13inter4));
  nand2 gate2708(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2709(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2710(.a(G9), .O(gate13inter7));
  inv1  gate2711(.a(G10), .O(gate13inter8));
  nand2 gate2712(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2713(.a(s_309), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2714(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2715(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2716(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1891(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1892(.a(gate15inter0), .b(s_192), .O(gate15inter1));
  and2  gate1893(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1894(.a(s_192), .O(gate15inter3));
  inv1  gate1895(.a(s_193), .O(gate15inter4));
  nand2 gate1896(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1897(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1898(.a(G13), .O(gate15inter7));
  inv1  gate1899(.a(G14), .O(gate15inter8));
  nand2 gate1900(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1901(.a(s_193), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1902(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1903(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1904(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1401(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1402(.a(gate16inter0), .b(s_122), .O(gate16inter1));
  and2  gate1403(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1404(.a(s_122), .O(gate16inter3));
  inv1  gate1405(.a(s_123), .O(gate16inter4));
  nand2 gate1406(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1407(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1408(.a(G15), .O(gate16inter7));
  inv1  gate1409(.a(G16), .O(gate16inter8));
  nand2 gate1410(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1411(.a(s_123), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1412(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1413(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1414(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1191(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1192(.a(gate23inter0), .b(s_92), .O(gate23inter1));
  and2  gate1193(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1194(.a(s_92), .O(gate23inter3));
  inv1  gate1195(.a(s_93), .O(gate23inter4));
  nand2 gate1196(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1197(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1198(.a(G29), .O(gate23inter7));
  inv1  gate1199(.a(G30), .O(gate23inter8));
  nand2 gate1200(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1201(.a(s_93), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1202(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1203(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1204(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1093(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1094(.a(gate26inter0), .b(s_78), .O(gate26inter1));
  and2  gate1095(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1096(.a(s_78), .O(gate26inter3));
  inv1  gate1097(.a(s_79), .O(gate26inter4));
  nand2 gate1098(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1099(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1100(.a(G9), .O(gate26inter7));
  inv1  gate1101(.a(G13), .O(gate26inter8));
  nand2 gate1102(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1103(.a(s_79), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1104(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1105(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1106(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1849(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1850(.a(gate29inter0), .b(s_186), .O(gate29inter1));
  and2  gate1851(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1852(.a(s_186), .O(gate29inter3));
  inv1  gate1853(.a(s_187), .O(gate29inter4));
  nand2 gate1854(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1855(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1856(.a(G3), .O(gate29inter7));
  inv1  gate1857(.a(G7), .O(gate29inter8));
  nand2 gate1858(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1859(.a(s_187), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1860(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1861(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1862(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2395(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2396(.a(gate33inter0), .b(s_264), .O(gate33inter1));
  and2  gate2397(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2398(.a(s_264), .O(gate33inter3));
  inv1  gate2399(.a(s_265), .O(gate33inter4));
  nand2 gate2400(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2401(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2402(.a(G17), .O(gate33inter7));
  inv1  gate2403(.a(G21), .O(gate33inter8));
  nand2 gate2404(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2405(.a(s_265), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2406(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2407(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2408(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2661(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2662(.a(gate34inter0), .b(s_302), .O(gate34inter1));
  and2  gate2663(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2664(.a(s_302), .O(gate34inter3));
  inv1  gate2665(.a(s_303), .O(gate34inter4));
  nand2 gate2666(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2667(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2668(.a(G25), .O(gate34inter7));
  inv1  gate2669(.a(G29), .O(gate34inter8));
  nand2 gate2670(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2671(.a(s_303), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2672(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2673(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2674(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1597(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1598(.a(gate36inter0), .b(s_150), .O(gate36inter1));
  and2  gate1599(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1600(.a(s_150), .O(gate36inter3));
  inv1  gate1601(.a(s_151), .O(gate36inter4));
  nand2 gate1602(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1603(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1604(.a(G26), .O(gate36inter7));
  inv1  gate1605(.a(G30), .O(gate36inter8));
  nand2 gate1606(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1607(.a(s_151), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1608(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1609(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1610(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1289(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1290(.a(gate38inter0), .b(s_106), .O(gate38inter1));
  and2  gate1291(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1292(.a(s_106), .O(gate38inter3));
  inv1  gate1293(.a(s_107), .O(gate38inter4));
  nand2 gate1294(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1295(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1296(.a(G27), .O(gate38inter7));
  inv1  gate1297(.a(G31), .O(gate38inter8));
  nand2 gate1298(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1299(.a(s_107), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1300(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1301(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1302(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1527(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1528(.a(gate39inter0), .b(s_140), .O(gate39inter1));
  and2  gate1529(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1530(.a(s_140), .O(gate39inter3));
  inv1  gate1531(.a(s_141), .O(gate39inter4));
  nand2 gate1532(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1533(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1534(.a(G20), .O(gate39inter7));
  inv1  gate1535(.a(G24), .O(gate39inter8));
  nand2 gate1536(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1537(.a(s_141), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1538(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1539(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1540(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1303(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1304(.a(gate41inter0), .b(s_108), .O(gate41inter1));
  and2  gate1305(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1306(.a(s_108), .O(gate41inter3));
  inv1  gate1307(.a(s_109), .O(gate41inter4));
  nand2 gate1308(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1309(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1310(.a(G1), .O(gate41inter7));
  inv1  gate1311(.a(G266), .O(gate41inter8));
  nand2 gate1312(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1313(.a(s_109), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1314(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1315(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1316(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate631(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate632(.a(gate45inter0), .b(s_12), .O(gate45inter1));
  and2  gate633(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate634(.a(s_12), .O(gate45inter3));
  inv1  gate635(.a(s_13), .O(gate45inter4));
  nand2 gate636(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate637(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate638(.a(G5), .O(gate45inter7));
  inv1  gate639(.a(G272), .O(gate45inter8));
  nand2 gate640(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate641(.a(s_13), .b(gate45inter3), .O(gate45inter10));
  nor2  gate642(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate643(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate644(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2619(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2620(.a(gate47inter0), .b(s_296), .O(gate47inter1));
  and2  gate2621(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2622(.a(s_296), .O(gate47inter3));
  inv1  gate2623(.a(s_297), .O(gate47inter4));
  nand2 gate2624(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2625(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2626(.a(G7), .O(gate47inter7));
  inv1  gate2627(.a(G275), .O(gate47inter8));
  nand2 gate2628(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2629(.a(s_297), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2630(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2631(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2632(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2185(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2186(.a(gate51inter0), .b(s_234), .O(gate51inter1));
  and2  gate2187(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2188(.a(s_234), .O(gate51inter3));
  inv1  gate2189(.a(s_235), .O(gate51inter4));
  nand2 gate2190(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2191(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2192(.a(G11), .O(gate51inter7));
  inv1  gate2193(.a(G281), .O(gate51inter8));
  nand2 gate2194(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2195(.a(s_235), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2196(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2197(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2198(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate2213(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2214(.a(gate52inter0), .b(s_238), .O(gate52inter1));
  and2  gate2215(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2216(.a(s_238), .O(gate52inter3));
  inv1  gate2217(.a(s_239), .O(gate52inter4));
  nand2 gate2218(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2219(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2220(.a(G12), .O(gate52inter7));
  inv1  gate2221(.a(G281), .O(gate52inter8));
  nand2 gate2222(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2223(.a(s_239), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2224(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2225(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2226(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2115(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2116(.a(gate54inter0), .b(s_224), .O(gate54inter1));
  and2  gate2117(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2118(.a(s_224), .O(gate54inter3));
  inv1  gate2119(.a(s_225), .O(gate54inter4));
  nand2 gate2120(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2121(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2122(.a(G14), .O(gate54inter7));
  inv1  gate2123(.a(G284), .O(gate54inter8));
  nand2 gate2124(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2125(.a(s_225), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2126(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2127(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2128(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1695(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1696(.a(gate56inter0), .b(s_164), .O(gate56inter1));
  and2  gate1697(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1698(.a(s_164), .O(gate56inter3));
  inv1  gate1699(.a(s_165), .O(gate56inter4));
  nand2 gate1700(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1701(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1702(.a(G16), .O(gate56inter7));
  inv1  gate1703(.a(G287), .O(gate56inter8));
  nand2 gate1704(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1705(.a(s_165), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1706(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1707(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1708(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate855(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate856(.a(gate59inter0), .b(s_44), .O(gate59inter1));
  and2  gate857(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate858(.a(s_44), .O(gate59inter3));
  inv1  gate859(.a(s_45), .O(gate59inter4));
  nand2 gate860(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate861(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate862(.a(G19), .O(gate59inter7));
  inv1  gate863(.a(G293), .O(gate59inter8));
  nand2 gate864(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate865(.a(s_45), .b(gate59inter3), .O(gate59inter10));
  nor2  gate866(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate867(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate868(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1051(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1052(.a(gate60inter0), .b(s_72), .O(gate60inter1));
  and2  gate1053(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1054(.a(s_72), .O(gate60inter3));
  inv1  gate1055(.a(s_73), .O(gate60inter4));
  nand2 gate1056(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1057(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1058(.a(G20), .O(gate60inter7));
  inv1  gate1059(.a(G293), .O(gate60inter8));
  nand2 gate1060(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1061(.a(s_73), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1062(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1063(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1064(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1107(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1108(.a(gate63inter0), .b(s_80), .O(gate63inter1));
  and2  gate1109(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1110(.a(s_80), .O(gate63inter3));
  inv1  gate1111(.a(s_81), .O(gate63inter4));
  nand2 gate1112(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1113(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1114(.a(G23), .O(gate63inter7));
  inv1  gate1115(.a(G299), .O(gate63inter8));
  nand2 gate1116(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1117(.a(s_81), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1118(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1119(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1120(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate953(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate954(.a(gate66inter0), .b(s_58), .O(gate66inter1));
  and2  gate955(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate956(.a(s_58), .O(gate66inter3));
  inv1  gate957(.a(s_59), .O(gate66inter4));
  nand2 gate958(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate959(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate960(.a(G26), .O(gate66inter7));
  inv1  gate961(.a(G302), .O(gate66inter8));
  nand2 gate962(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate963(.a(s_59), .b(gate66inter3), .O(gate66inter10));
  nor2  gate964(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate965(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate966(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1275(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1276(.a(gate67inter0), .b(s_104), .O(gate67inter1));
  and2  gate1277(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1278(.a(s_104), .O(gate67inter3));
  inv1  gate1279(.a(s_105), .O(gate67inter4));
  nand2 gate1280(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1281(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1282(.a(G27), .O(gate67inter7));
  inv1  gate1283(.a(G305), .O(gate67inter8));
  nand2 gate1284(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1285(.a(s_105), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1286(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1287(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1288(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1653(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1654(.a(gate71inter0), .b(s_158), .O(gate71inter1));
  and2  gate1655(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1656(.a(s_158), .O(gate71inter3));
  inv1  gate1657(.a(s_159), .O(gate71inter4));
  nand2 gate1658(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1659(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1660(.a(G31), .O(gate71inter7));
  inv1  gate1661(.a(G311), .O(gate71inter8));
  nand2 gate1662(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1663(.a(s_159), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1664(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1665(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1666(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate2465(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2466(.a(gate73inter0), .b(s_274), .O(gate73inter1));
  and2  gate2467(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2468(.a(s_274), .O(gate73inter3));
  inv1  gate2469(.a(s_275), .O(gate73inter4));
  nand2 gate2470(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2471(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2472(.a(G1), .O(gate73inter7));
  inv1  gate2473(.a(G314), .O(gate73inter8));
  nand2 gate2474(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2475(.a(s_275), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2476(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2477(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2478(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1457(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1458(.a(gate74inter0), .b(s_130), .O(gate74inter1));
  and2  gate1459(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1460(.a(s_130), .O(gate74inter3));
  inv1  gate1461(.a(s_131), .O(gate74inter4));
  nand2 gate1462(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1463(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1464(.a(G5), .O(gate74inter7));
  inv1  gate1465(.a(G314), .O(gate74inter8));
  nand2 gate1466(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1467(.a(s_131), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1468(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1469(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1470(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1205(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1206(.a(gate80inter0), .b(s_94), .O(gate80inter1));
  and2  gate1207(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1208(.a(s_94), .O(gate80inter3));
  inv1  gate1209(.a(s_95), .O(gate80inter4));
  nand2 gate1210(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1211(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1212(.a(G14), .O(gate80inter7));
  inv1  gate1213(.a(G323), .O(gate80inter8));
  nand2 gate1214(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1215(.a(s_95), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1216(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1217(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1218(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2577(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2578(.a(gate81inter0), .b(s_290), .O(gate81inter1));
  and2  gate2579(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2580(.a(s_290), .O(gate81inter3));
  inv1  gate2581(.a(s_291), .O(gate81inter4));
  nand2 gate2582(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2583(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2584(.a(G3), .O(gate81inter7));
  inv1  gate2585(.a(G326), .O(gate81inter8));
  nand2 gate2586(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2587(.a(s_291), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2588(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2589(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2590(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2367(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2368(.a(gate84inter0), .b(s_260), .O(gate84inter1));
  and2  gate2369(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2370(.a(s_260), .O(gate84inter3));
  inv1  gate2371(.a(s_261), .O(gate84inter4));
  nand2 gate2372(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2373(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2374(.a(G15), .O(gate84inter7));
  inv1  gate2375(.a(G329), .O(gate84inter8));
  nand2 gate2376(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2377(.a(s_261), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2378(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2379(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2380(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2227(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2228(.a(gate86inter0), .b(s_240), .O(gate86inter1));
  and2  gate2229(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2230(.a(s_240), .O(gate86inter3));
  inv1  gate2231(.a(s_241), .O(gate86inter4));
  nand2 gate2232(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2233(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2234(.a(G8), .O(gate86inter7));
  inv1  gate2235(.a(G332), .O(gate86inter8));
  nand2 gate2236(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2237(.a(s_241), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2238(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2239(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2240(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1933(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1934(.a(gate90inter0), .b(s_198), .O(gate90inter1));
  and2  gate1935(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1936(.a(s_198), .O(gate90inter3));
  inv1  gate1937(.a(s_199), .O(gate90inter4));
  nand2 gate1938(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1939(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1940(.a(G21), .O(gate90inter7));
  inv1  gate1941(.a(G338), .O(gate90inter8));
  nand2 gate1942(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1943(.a(s_199), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1944(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1945(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1946(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1723(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1724(.a(gate91inter0), .b(s_168), .O(gate91inter1));
  and2  gate1725(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1726(.a(s_168), .O(gate91inter3));
  inv1  gate1727(.a(s_169), .O(gate91inter4));
  nand2 gate1728(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1729(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1730(.a(G25), .O(gate91inter7));
  inv1  gate1731(.a(G341), .O(gate91inter8));
  nand2 gate1732(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1733(.a(s_169), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1734(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1735(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1736(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2647(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2648(.a(gate94inter0), .b(s_300), .O(gate94inter1));
  and2  gate2649(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2650(.a(s_300), .O(gate94inter3));
  inv1  gate2651(.a(s_301), .O(gate94inter4));
  nand2 gate2652(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2653(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2654(.a(G22), .O(gate94inter7));
  inv1  gate2655(.a(G344), .O(gate94inter8));
  nand2 gate2656(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2657(.a(s_301), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2658(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2659(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2660(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1485(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1486(.a(gate96inter0), .b(s_134), .O(gate96inter1));
  and2  gate1487(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1488(.a(s_134), .O(gate96inter3));
  inv1  gate1489(.a(s_135), .O(gate96inter4));
  nand2 gate1490(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1491(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1492(.a(G30), .O(gate96inter7));
  inv1  gate1493(.a(G347), .O(gate96inter8));
  nand2 gate1494(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1495(.a(s_135), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1496(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1497(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1498(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate701(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate702(.a(gate99inter0), .b(s_22), .O(gate99inter1));
  and2  gate703(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate704(.a(s_22), .O(gate99inter3));
  inv1  gate705(.a(s_23), .O(gate99inter4));
  nand2 gate706(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate707(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate708(.a(G27), .O(gate99inter7));
  inv1  gate709(.a(G353), .O(gate99inter8));
  nand2 gate710(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate711(.a(s_23), .b(gate99inter3), .O(gate99inter10));
  nor2  gate712(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate713(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate714(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2353(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2354(.a(gate107inter0), .b(s_258), .O(gate107inter1));
  and2  gate2355(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2356(.a(s_258), .O(gate107inter3));
  inv1  gate2357(.a(s_259), .O(gate107inter4));
  nand2 gate2358(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2359(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2360(.a(G366), .O(gate107inter7));
  inv1  gate2361(.a(G367), .O(gate107inter8));
  nand2 gate2362(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2363(.a(s_259), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2364(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2365(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2366(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1219(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1220(.a(gate108inter0), .b(s_96), .O(gate108inter1));
  and2  gate1221(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1222(.a(s_96), .O(gate108inter3));
  inv1  gate1223(.a(s_97), .O(gate108inter4));
  nand2 gate1224(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1225(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1226(.a(G368), .O(gate108inter7));
  inv1  gate1227(.a(G369), .O(gate108inter8));
  nand2 gate1228(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1229(.a(s_97), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1230(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1231(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1232(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1331(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1332(.a(gate114inter0), .b(s_112), .O(gate114inter1));
  and2  gate1333(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1334(.a(s_112), .O(gate114inter3));
  inv1  gate1335(.a(s_113), .O(gate114inter4));
  nand2 gate1336(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1337(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1338(.a(G380), .O(gate114inter7));
  inv1  gate1339(.a(G381), .O(gate114inter8));
  nand2 gate1340(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1341(.a(s_113), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1342(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1343(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1344(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1233(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1234(.a(gate115inter0), .b(s_98), .O(gate115inter1));
  and2  gate1235(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1236(.a(s_98), .O(gate115inter3));
  inv1  gate1237(.a(s_99), .O(gate115inter4));
  nand2 gate1238(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1239(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1240(.a(G382), .O(gate115inter7));
  inv1  gate1241(.a(G383), .O(gate115inter8));
  nand2 gate1242(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1243(.a(s_99), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1244(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1245(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1246(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate2605(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2606(.a(gate116inter0), .b(s_294), .O(gate116inter1));
  and2  gate2607(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2608(.a(s_294), .O(gate116inter3));
  inv1  gate2609(.a(s_295), .O(gate116inter4));
  nand2 gate2610(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2611(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2612(.a(G384), .O(gate116inter7));
  inv1  gate2613(.a(G385), .O(gate116inter8));
  nand2 gate2614(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2615(.a(s_295), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2616(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2617(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2618(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate785(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate786(.a(gate117inter0), .b(s_34), .O(gate117inter1));
  and2  gate787(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate788(.a(s_34), .O(gate117inter3));
  inv1  gate789(.a(s_35), .O(gate117inter4));
  nand2 gate790(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate791(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate792(.a(G386), .O(gate117inter7));
  inv1  gate793(.a(G387), .O(gate117inter8));
  nand2 gate794(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate795(.a(s_35), .b(gate117inter3), .O(gate117inter10));
  nor2  gate796(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate797(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate798(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate981(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate982(.a(gate119inter0), .b(s_62), .O(gate119inter1));
  and2  gate983(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate984(.a(s_62), .O(gate119inter3));
  inv1  gate985(.a(s_63), .O(gate119inter4));
  nand2 gate986(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate987(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate988(.a(G390), .O(gate119inter7));
  inv1  gate989(.a(G391), .O(gate119inter8));
  nand2 gate990(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate991(.a(s_63), .b(gate119inter3), .O(gate119inter10));
  nor2  gate992(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate993(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate994(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate2717(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate2718(.a(gate123inter0), .b(s_310), .O(gate123inter1));
  and2  gate2719(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate2720(.a(s_310), .O(gate123inter3));
  inv1  gate2721(.a(s_311), .O(gate123inter4));
  nand2 gate2722(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate2723(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate2724(.a(G398), .O(gate123inter7));
  inv1  gate2725(.a(G399), .O(gate123inter8));
  nand2 gate2726(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate2727(.a(s_311), .b(gate123inter3), .O(gate123inter10));
  nor2  gate2728(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate2729(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate2730(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1429(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1430(.a(gate124inter0), .b(s_126), .O(gate124inter1));
  and2  gate1431(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1432(.a(s_126), .O(gate124inter3));
  inv1  gate1433(.a(s_127), .O(gate124inter4));
  nand2 gate1434(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1435(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1436(.a(G400), .O(gate124inter7));
  inv1  gate1437(.a(G401), .O(gate124inter8));
  nand2 gate1438(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1439(.a(s_127), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1440(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1441(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1442(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1975(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1976(.a(gate125inter0), .b(s_204), .O(gate125inter1));
  and2  gate1977(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1978(.a(s_204), .O(gate125inter3));
  inv1  gate1979(.a(s_205), .O(gate125inter4));
  nand2 gate1980(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1981(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1982(.a(G402), .O(gate125inter7));
  inv1  gate1983(.a(G403), .O(gate125inter8));
  nand2 gate1984(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1985(.a(s_205), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1986(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1987(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1988(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1471(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1472(.a(gate132inter0), .b(s_132), .O(gate132inter1));
  and2  gate1473(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1474(.a(s_132), .O(gate132inter3));
  inv1  gate1475(.a(s_133), .O(gate132inter4));
  nand2 gate1476(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1477(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1478(.a(G416), .O(gate132inter7));
  inv1  gate1479(.a(G417), .O(gate132inter8));
  nand2 gate1480(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1481(.a(s_133), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1482(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1483(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1484(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate617(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate618(.a(gate135inter0), .b(s_10), .O(gate135inter1));
  and2  gate619(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate620(.a(s_10), .O(gate135inter3));
  inv1  gate621(.a(s_11), .O(gate135inter4));
  nand2 gate622(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate623(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate624(.a(G422), .O(gate135inter7));
  inv1  gate625(.a(G423), .O(gate135inter8));
  nand2 gate626(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate627(.a(s_11), .b(gate135inter3), .O(gate135inter10));
  nor2  gate628(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate629(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate630(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1569(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1570(.a(gate137inter0), .b(s_146), .O(gate137inter1));
  and2  gate1571(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1572(.a(s_146), .O(gate137inter3));
  inv1  gate1573(.a(s_147), .O(gate137inter4));
  nand2 gate1574(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1575(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1576(.a(G426), .O(gate137inter7));
  inv1  gate1577(.a(G429), .O(gate137inter8));
  nand2 gate1578(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1579(.a(s_147), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1580(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1581(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1582(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate673(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate674(.a(gate144inter0), .b(s_18), .O(gate144inter1));
  and2  gate675(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate676(.a(s_18), .O(gate144inter3));
  inv1  gate677(.a(s_19), .O(gate144inter4));
  nand2 gate678(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate679(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate680(.a(G468), .O(gate144inter7));
  inv1  gate681(.a(G471), .O(gate144inter8));
  nand2 gate682(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate683(.a(s_19), .b(gate144inter3), .O(gate144inter10));
  nor2  gate684(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate685(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate686(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate589(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate590(.a(gate145inter0), .b(s_6), .O(gate145inter1));
  and2  gate591(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate592(.a(s_6), .O(gate145inter3));
  inv1  gate593(.a(s_7), .O(gate145inter4));
  nand2 gate594(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate595(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate596(.a(G474), .O(gate145inter7));
  inv1  gate597(.a(G477), .O(gate145inter8));
  nand2 gate598(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate599(.a(s_7), .b(gate145inter3), .O(gate145inter10));
  nor2  gate600(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate601(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate602(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1499(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1500(.a(gate149inter0), .b(s_136), .O(gate149inter1));
  and2  gate1501(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1502(.a(s_136), .O(gate149inter3));
  inv1  gate1503(.a(s_137), .O(gate149inter4));
  nand2 gate1504(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1505(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1506(.a(G498), .O(gate149inter7));
  inv1  gate1507(.a(G501), .O(gate149inter8));
  nand2 gate1508(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1509(.a(s_137), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1510(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1511(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1512(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate827(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate828(.a(gate152inter0), .b(s_40), .O(gate152inter1));
  and2  gate829(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate830(.a(s_40), .O(gate152inter3));
  inv1  gate831(.a(s_41), .O(gate152inter4));
  nand2 gate832(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate833(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate834(.a(G516), .O(gate152inter7));
  inv1  gate835(.a(G519), .O(gate152inter8));
  nand2 gate836(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate837(.a(s_41), .b(gate152inter3), .O(gate152inter10));
  nor2  gate838(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate839(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate840(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2311(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2312(.a(gate154inter0), .b(s_252), .O(gate154inter1));
  and2  gate2313(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2314(.a(s_252), .O(gate154inter3));
  inv1  gate2315(.a(s_253), .O(gate154inter4));
  nand2 gate2316(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2317(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2318(.a(G429), .O(gate154inter7));
  inv1  gate2319(.a(G522), .O(gate154inter8));
  nand2 gate2320(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2321(.a(s_253), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2322(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2323(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2324(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2451(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2452(.a(gate155inter0), .b(s_272), .O(gate155inter1));
  and2  gate2453(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2454(.a(s_272), .O(gate155inter3));
  inv1  gate2455(.a(s_273), .O(gate155inter4));
  nand2 gate2456(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2457(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2458(.a(G432), .O(gate155inter7));
  inv1  gate2459(.a(G525), .O(gate155inter8));
  nand2 gate2460(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2461(.a(s_273), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2462(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2463(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2464(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate799(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate800(.a(gate159inter0), .b(s_36), .O(gate159inter1));
  and2  gate801(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate802(.a(s_36), .O(gate159inter3));
  inv1  gate803(.a(s_37), .O(gate159inter4));
  nand2 gate804(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate805(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate806(.a(G444), .O(gate159inter7));
  inv1  gate807(.a(G531), .O(gate159inter8));
  nand2 gate808(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate809(.a(s_37), .b(gate159inter3), .O(gate159inter10));
  nor2  gate810(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate811(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate812(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2563(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2564(.a(gate161inter0), .b(s_288), .O(gate161inter1));
  and2  gate2565(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2566(.a(s_288), .O(gate161inter3));
  inv1  gate2567(.a(s_289), .O(gate161inter4));
  nand2 gate2568(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2569(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2570(.a(G450), .O(gate161inter7));
  inv1  gate2571(.a(G534), .O(gate161inter8));
  nand2 gate2572(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2573(.a(s_289), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2574(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2575(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2576(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1177(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1178(.a(gate162inter0), .b(s_90), .O(gate162inter1));
  and2  gate1179(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1180(.a(s_90), .O(gate162inter3));
  inv1  gate1181(.a(s_91), .O(gate162inter4));
  nand2 gate1182(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1183(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1184(.a(G453), .O(gate162inter7));
  inv1  gate1185(.a(G534), .O(gate162inter8));
  nand2 gate1186(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1187(.a(s_91), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1188(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1189(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1190(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate1779(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1780(.a(gate163inter0), .b(s_176), .O(gate163inter1));
  and2  gate1781(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1782(.a(s_176), .O(gate163inter3));
  inv1  gate1783(.a(s_177), .O(gate163inter4));
  nand2 gate1784(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1785(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1786(.a(G456), .O(gate163inter7));
  inv1  gate1787(.a(G537), .O(gate163inter8));
  nand2 gate1788(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1789(.a(s_177), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1790(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1791(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1792(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1163(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1164(.a(gate169inter0), .b(s_88), .O(gate169inter1));
  and2  gate1165(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1166(.a(s_88), .O(gate169inter3));
  inv1  gate1167(.a(s_89), .O(gate169inter4));
  nand2 gate1168(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1169(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1170(.a(G474), .O(gate169inter7));
  inv1  gate1171(.a(G546), .O(gate169inter8));
  nand2 gate1172(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1173(.a(s_89), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1174(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1175(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1176(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1821(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1822(.a(gate171inter0), .b(s_182), .O(gate171inter1));
  and2  gate1823(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1824(.a(s_182), .O(gate171inter3));
  inv1  gate1825(.a(s_183), .O(gate171inter4));
  nand2 gate1826(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1827(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1828(.a(G480), .O(gate171inter7));
  inv1  gate1829(.a(G549), .O(gate171inter8));
  nand2 gate1830(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1831(.a(s_183), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1832(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1833(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1834(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate729(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate730(.a(gate172inter0), .b(s_26), .O(gate172inter1));
  and2  gate731(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate732(.a(s_26), .O(gate172inter3));
  inv1  gate733(.a(s_27), .O(gate172inter4));
  nand2 gate734(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate735(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate736(.a(G483), .O(gate172inter7));
  inv1  gate737(.a(G549), .O(gate172inter8));
  nand2 gate738(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate739(.a(s_27), .b(gate172inter3), .O(gate172inter10));
  nor2  gate740(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate741(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate742(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1877(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1878(.a(gate175inter0), .b(s_190), .O(gate175inter1));
  and2  gate1879(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1880(.a(s_190), .O(gate175inter3));
  inv1  gate1881(.a(s_191), .O(gate175inter4));
  nand2 gate1882(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1883(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1884(.a(G492), .O(gate175inter7));
  inv1  gate1885(.a(G555), .O(gate175inter8));
  nand2 gate1886(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1887(.a(s_191), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1888(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1889(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1890(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1583(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1584(.a(gate181inter0), .b(s_148), .O(gate181inter1));
  and2  gate1585(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1586(.a(s_148), .O(gate181inter3));
  inv1  gate1587(.a(s_149), .O(gate181inter4));
  nand2 gate1588(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1589(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1590(.a(G510), .O(gate181inter7));
  inv1  gate1591(.a(G564), .O(gate181inter8));
  nand2 gate1592(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1593(.a(s_149), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1594(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1595(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1596(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1737(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1738(.a(gate183inter0), .b(s_170), .O(gate183inter1));
  and2  gate1739(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1740(.a(s_170), .O(gate183inter3));
  inv1  gate1741(.a(s_171), .O(gate183inter4));
  nand2 gate1742(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1743(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1744(.a(G516), .O(gate183inter7));
  inv1  gate1745(.a(G567), .O(gate183inter8));
  nand2 gate1746(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1747(.a(s_171), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1748(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1749(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1750(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2101(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2102(.a(gate185inter0), .b(s_222), .O(gate185inter1));
  and2  gate2103(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2104(.a(s_222), .O(gate185inter3));
  inv1  gate2105(.a(s_223), .O(gate185inter4));
  nand2 gate2106(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2107(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2108(.a(G570), .O(gate185inter7));
  inv1  gate2109(.a(G571), .O(gate185inter8));
  nand2 gate2110(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2111(.a(s_223), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2112(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2113(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2114(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1919(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1920(.a(gate186inter0), .b(s_196), .O(gate186inter1));
  and2  gate1921(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1922(.a(s_196), .O(gate186inter3));
  inv1  gate1923(.a(s_197), .O(gate186inter4));
  nand2 gate1924(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1925(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1926(.a(G572), .O(gate186inter7));
  inv1  gate1927(.a(G573), .O(gate186inter8));
  nand2 gate1928(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1929(.a(s_197), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1930(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1931(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1932(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate939(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate940(.a(gate187inter0), .b(s_56), .O(gate187inter1));
  and2  gate941(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate942(.a(s_56), .O(gate187inter3));
  inv1  gate943(.a(s_57), .O(gate187inter4));
  nand2 gate944(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate945(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate946(.a(G574), .O(gate187inter7));
  inv1  gate947(.a(G575), .O(gate187inter8));
  nand2 gate948(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate949(.a(s_57), .b(gate187inter3), .O(gate187inter10));
  nor2  gate950(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate951(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate952(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1793(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1794(.a(gate191inter0), .b(s_178), .O(gate191inter1));
  and2  gate1795(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1796(.a(s_178), .O(gate191inter3));
  inv1  gate1797(.a(s_179), .O(gate191inter4));
  nand2 gate1798(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1799(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1800(.a(G582), .O(gate191inter7));
  inv1  gate1801(.a(G583), .O(gate191inter8));
  nand2 gate1802(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1803(.a(s_179), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1804(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1805(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1806(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate869(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate870(.a(gate199inter0), .b(s_46), .O(gate199inter1));
  and2  gate871(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate872(.a(s_46), .O(gate199inter3));
  inv1  gate873(.a(s_47), .O(gate199inter4));
  nand2 gate874(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate875(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate876(.a(G598), .O(gate199inter7));
  inv1  gate877(.a(G599), .O(gate199inter8));
  nand2 gate878(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate879(.a(s_47), .b(gate199inter3), .O(gate199inter10));
  nor2  gate880(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate881(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate882(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2017(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2018(.a(gate201inter0), .b(s_210), .O(gate201inter1));
  and2  gate2019(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2020(.a(s_210), .O(gate201inter3));
  inv1  gate2021(.a(s_211), .O(gate201inter4));
  nand2 gate2022(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2023(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2024(.a(G602), .O(gate201inter7));
  inv1  gate2025(.a(G607), .O(gate201inter8));
  nand2 gate2026(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2027(.a(s_211), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2028(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2029(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2030(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1121(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1122(.a(gate203inter0), .b(s_82), .O(gate203inter1));
  and2  gate1123(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1124(.a(s_82), .O(gate203inter3));
  inv1  gate1125(.a(s_83), .O(gate203inter4));
  nand2 gate1126(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1127(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1128(.a(G602), .O(gate203inter7));
  inv1  gate1129(.a(G612), .O(gate203inter8));
  nand2 gate1130(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1131(.a(s_83), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1132(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1133(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1134(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1709(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1710(.a(gate205inter0), .b(s_166), .O(gate205inter1));
  and2  gate1711(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1712(.a(s_166), .O(gate205inter3));
  inv1  gate1713(.a(s_167), .O(gate205inter4));
  nand2 gate1714(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1715(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1716(.a(G622), .O(gate205inter7));
  inv1  gate1717(.a(G627), .O(gate205inter8));
  nand2 gate1718(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1719(.a(s_167), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1720(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1721(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1722(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1751(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1752(.a(gate206inter0), .b(s_172), .O(gate206inter1));
  and2  gate1753(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1754(.a(s_172), .O(gate206inter3));
  inv1  gate1755(.a(s_173), .O(gate206inter4));
  nand2 gate1756(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1757(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1758(.a(G632), .O(gate206inter7));
  inv1  gate1759(.a(G637), .O(gate206inter8));
  nand2 gate1760(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1761(.a(s_173), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1762(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1763(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1764(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1443(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1444(.a(gate207inter0), .b(s_128), .O(gate207inter1));
  and2  gate1445(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1446(.a(s_128), .O(gate207inter3));
  inv1  gate1447(.a(s_129), .O(gate207inter4));
  nand2 gate1448(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1449(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1450(.a(G622), .O(gate207inter7));
  inv1  gate1451(.a(G632), .O(gate207inter8));
  nand2 gate1452(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1453(.a(s_129), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1454(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1455(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1456(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate883(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate884(.a(gate211inter0), .b(s_48), .O(gate211inter1));
  and2  gate885(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate886(.a(s_48), .O(gate211inter3));
  inv1  gate887(.a(s_49), .O(gate211inter4));
  nand2 gate888(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate889(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate890(.a(G612), .O(gate211inter7));
  inv1  gate891(.a(G669), .O(gate211inter8));
  nand2 gate892(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate893(.a(s_49), .b(gate211inter3), .O(gate211inter10));
  nor2  gate894(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate895(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate896(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1947(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1948(.a(gate216inter0), .b(s_200), .O(gate216inter1));
  and2  gate1949(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1950(.a(s_200), .O(gate216inter3));
  inv1  gate1951(.a(s_201), .O(gate216inter4));
  nand2 gate1952(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1953(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1954(.a(G617), .O(gate216inter7));
  inv1  gate1955(.a(G675), .O(gate216inter8));
  nand2 gate1956(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1957(.a(s_201), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1958(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1959(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1960(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1079(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1080(.a(gate218inter0), .b(s_76), .O(gate218inter1));
  and2  gate1081(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1082(.a(s_76), .O(gate218inter3));
  inv1  gate1083(.a(s_77), .O(gate218inter4));
  nand2 gate1084(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1085(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1086(.a(G627), .O(gate218inter7));
  inv1  gate1087(.a(G678), .O(gate218inter8));
  nand2 gate1088(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1089(.a(s_77), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1090(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1091(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1092(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1961(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1962(.a(gate221inter0), .b(s_202), .O(gate221inter1));
  and2  gate1963(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1964(.a(s_202), .O(gate221inter3));
  inv1  gate1965(.a(s_203), .O(gate221inter4));
  nand2 gate1966(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1967(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1968(.a(G622), .O(gate221inter7));
  inv1  gate1969(.a(G684), .O(gate221inter8));
  nand2 gate1970(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1971(.a(s_203), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1972(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1973(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1974(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2255(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2256(.a(gate224inter0), .b(s_244), .O(gate224inter1));
  and2  gate2257(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2258(.a(s_244), .O(gate224inter3));
  inv1  gate2259(.a(s_245), .O(gate224inter4));
  nand2 gate2260(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2261(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2262(.a(G637), .O(gate224inter7));
  inv1  gate2263(.a(G687), .O(gate224inter8));
  nand2 gate2264(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2265(.a(s_245), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2266(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2267(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2268(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2059(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2060(.a(gate227inter0), .b(s_216), .O(gate227inter1));
  and2  gate2061(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2062(.a(s_216), .O(gate227inter3));
  inv1  gate2063(.a(s_217), .O(gate227inter4));
  nand2 gate2064(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2065(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2066(.a(G694), .O(gate227inter7));
  inv1  gate2067(.a(G695), .O(gate227inter8));
  nand2 gate2068(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2069(.a(s_217), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2070(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2071(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2072(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2689(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2690(.a(gate229inter0), .b(s_306), .O(gate229inter1));
  and2  gate2691(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2692(.a(s_306), .O(gate229inter3));
  inv1  gate2693(.a(s_307), .O(gate229inter4));
  nand2 gate2694(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2695(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2696(.a(G698), .O(gate229inter7));
  inv1  gate2697(.a(G699), .O(gate229inter8));
  nand2 gate2698(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2699(.a(s_307), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2700(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2701(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2702(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate2437(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2438(.a(gate230inter0), .b(s_270), .O(gate230inter1));
  and2  gate2439(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2440(.a(s_270), .O(gate230inter3));
  inv1  gate2441(.a(s_271), .O(gate230inter4));
  nand2 gate2442(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2443(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2444(.a(G700), .O(gate230inter7));
  inv1  gate2445(.a(G701), .O(gate230inter8));
  nand2 gate2446(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2447(.a(s_271), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2448(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2449(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2450(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1345(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1346(.a(gate232inter0), .b(s_114), .O(gate232inter1));
  and2  gate1347(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1348(.a(s_114), .O(gate232inter3));
  inv1  gate1349(.a(s_115), .O(gate232inter4));
  nand2 gate1350(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1351(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1352(.a(G704), .O(gate232inter7));
  inv1  gate1353(.a(G705), .O(gate232inter8));
  nand2 gate1354(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1355(.a(s_115), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1356(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1357(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1358(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate2143(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2144(.a(gate235inter0), .b(s_228), .O(gate235inter1));
  and2  gate2145(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2146(.a(s_228), .O(gate235inter3));
  inv1  gate2147(.a(s_229), .O(gate235inter4));
  nand2 gate2148(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2149(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2150(.a(G248), .O(gate235inter7));
  inv1  gate2151(.a(G724), .O(gate235inter8));
  nand2 gate2152(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2153(.a(s_229), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2154(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2155(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2156(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate645(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate646(.a(gate241inter0), .b(s_14), .O(gate241inter1));
  and2  gate647(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate648(.a(s_14), .O(gate241inter3));
  inv1  gate649(.a(s_15), .O(gate241inter4));
  nand2 gate650(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate651(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate652(.a(G242), .O(gate241inter7));
  inv1  gate653(.a(G730), .O(gate241inter8));
  nand2 gate654(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate655(.a(s_15), .b(gate241inter3), .O(gate241inter10));
  nor2  gate656(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate657(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate658(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate547(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate548(.a(gate242inter0), .b(s_0), .O(gate242inter1));
  and2  gate549(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate550(.a(s_0), .O(gate242inter3));
  inv1  gate551(.a(s_1), .O(gate242inter4));
  nand2 gate552(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate553(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate554(.a(G718), .O(gate242inter7));
  inv1  gate555(.a(G730), .O(gate242inter8));
  nand2 gate556(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate557(.a(s_1), .b(gate242inter3), .O(gate242inter10));
  nor2  gate558(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate559(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate560(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1863(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1864(.a(gate243inter0), .b(s_188), .O(gate243inter1));
  and2  gate1865(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1866(.a(s_188), .O(gate243inter3));
  inv1  gate1867(.a(s_189), .O(gate243inter4));
  nand2 gate1868(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1869(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1870(.a(G245), .O(gate243inter7));
  inv1  gate1871(.a(G733), .O(gate243inter8));
  nand2 gate1872(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1873(.a(s_189), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1874(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1875(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1876(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2591(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2592(.a(gate245inter0), .b(s_292), .O(gate245inter1));
  and2  gate2593(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2594(.a(s_292), .O(gate245inter3));
  inv1  gate2595(.a(s_293), .O(gate245inter4));
  nand2 gate2596(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2597(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2598(.a(G248), .O(gate245inter7));
  inv1  gate2599(.a(G736), .O(gate245inter8));
  nand2 gate2600(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2601(.a(s_293), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2602(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2603(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2604(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1149(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1150(.a(gate246inter0), .b(s_86), .O(gate246inter1));
  and2  gate1151(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1152(.a(s_86), .O(gate246inter3));
  inv1  gate1153(.a(s_87), .O(gate246inter4));
  nand2 gate1154(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1155(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1156(.a(G724), .O(gate246inter7));
  inv1  gate1157(.a(G736), .O(gate246inter8));
  nand2 gate1158(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1159(.a(s_87), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1160(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1161(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1162(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1905(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1906(.a(gate252inter0), .b(s_194), .O(gate252inter1));
  and2  gate1907(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1908(.a(s_194), .O(gate252inter3));
  inv1  gate1909(.a(s_195), .O(gate252inter4));
  nand2 gate1910(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1911(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1912(.a(G709), .O(gate252inter7));
  inv1  gate1913(.a(G745), .O(gate252inter8));
  nand2 gate1914(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1915(.a(s_195), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1916(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1917(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1918(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1415(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1416(.a(gate260inter0), .b(s_124), .O(gate260inter1));
  and2  gate1417(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1418(.a(s_124), .O(gate260inter3));
  inv1  gate1419(.a(s_125), .O(gate260inter4));
  nand2 gate1420(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1421(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1422(.a(G760), .O(gate260inter7));
  inv1  gate1423(.a(G761), .O(gate260inter8));
  nand2 gate1424(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1425(.a(s_125), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1426(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1427(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1428(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate995(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate996(.a(gate267inter0), .b(s_64), .O(gate267inter1));
  and2  gate997(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate998(.a(s_64), .O(gate267inter3));
  inv1  gate999(.a(s_65), .O(gate267inter4));
  nand2 gate1000(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1001(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1002(.a(G648), .O(gate267inter7));
  inv1  gate1003(.a(G776), .O(gate267inter8));
  nand2 gate1004(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1005(.a(s_65), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1006(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1007(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1008(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1359(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1360(.a(gate270inter0), .b(s_116), .O(gate270inter1));
  and2  gate1361(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1362(.a(s_116), .O(gate270inter3));
  inv1  gate1363(.a(s_117), .O(gate270inter4));
  nand2 gate1364(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1365(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1366(.a(G657), .O(gate270inter7));
  inv1  gate1367(.a(G785), .O(gate270inter8));
  nand2 gate1368(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1369(.a(s_117), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1370(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1371(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1372(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2073(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2074(.a(gate271inter0), .b(s_218), .O(gate271inter1));
  and2  gate2075(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2076(.a(s_218), .O(gate271inter3));
  inv1  gate2077(.a(s_219), .O(gate271inter4));
  nand2 gate2078(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2079(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2080(.a(G660), .O(gate271inter7));
  inv1  gate2081(.a(G788), .O(gate271inter8));
  nand2 gate2082(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2083(.a(s_219), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2084(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2085(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2086(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2381(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2382(.a(gate272inter0), .b(s_262), .O(gate272inter1));
  and2  gate2383(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2384(.a(s_262), .O(gate272inter3));
  inv1  gate2385(.a(s_263), .O(gate272inter4));
  nand2 gate2386(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2387(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2388(.a(G663), .O(gate272inter7));
  inv1  gate2389(.a(G791), .O(gate272inter8));
  nand2 gate2390(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2391(.a(s_263), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2392(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2393(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2394(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate561(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate562(.a(gate273inter0), .b(s_2), .O(gate273inter1));
  and2  gate563(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate564(.a(s_2), .O(gate273inter3));
  inv1  gate565(.a(s_3), .O(gate273inter4));
  nand2 gate566(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate567(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate568(.a(G642), .O(gate273inter7));
  inv1  gate569(.a(G794), .O(gate273inter8));
  nand2 gate570(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate571(.a(s_3), .b(gate273inter3), .O(gate273inter10));
  nor2  gate572(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate573(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate574(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1135(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1136(.a(gate275inter0), .b(s_84), .O(gate275inter1));
  and2  gate1137(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1138(.a(s_84), .O(gate275inter3));
  inv1  gate1139(.a(s_85), .O(gate275inter4));
  nand2 gate1140(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1141(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1142(.a(G645), .O(gate275inter7));
  inv1  gate1143(.a(G797), .O(gate275inter8));
  nand2 gate1144(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1145(.a(s_85), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1146(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1147(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1148(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate2675(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2676(.a(gate276inter0), .b(s_304), .O(gate276inter1));
  and2  gate2677(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2678(.a(s_304), .O(gate276inter3));
  inv1  gate2679(.a(s_305), .O(gate276inter4));
  nand2 gate2680(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2681(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2682(.a(G773), .O(gate276inter7));
  inv1  gate2683(.a(G797), .O(gate276inter8));
  nand2 gate2684(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2685(.a(s_305), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2686(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2687(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2688(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate757(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate758(.a(gate279inter0), .b(s_30), .O(gate279inter1));
  and2  gate759(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate760(.a(s_30), .O(gate279inter3));
  inv1  gate761(.a(s_31), .O(gate279inter4));
  nand2 gate762(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate763(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate764(.a(G651), .O(gate279inter7));
  inv1  gate765(.a(G803), .O(gate279inter8));
  nand2 gate766(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate767(.a(s_31), .b(gate279inter3), .O(gate279inter10));
  nor2  gate768(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate769(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate770(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2339(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2340(.a(gate289inter0), .b(s_256), .O(gate289inter1));
  and2  gate2341(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2342(.a(s_256), .O(gate289inter3));
  inv1  gate2343(.a(s_257), .O(gate289inter4));
  nand2 gate2344(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2345(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2346(.a(G818), .O(gate289inter7));
  inv1  gate2347(.a(G819), .O(gate289inter8));
  nand2 gate2348(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2349(.a(s_257), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2350(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2351(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2352(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2087(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2088(.a(gate291inter0), .b(s_220), .O(gate291inter1));
  and2  gate2089(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2090(.a(s_220), .O(gate291inter3));
  inv1  gate2091(.a(s_221), .O(gate291inter4));
  nand2 gate2092(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2093(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2094(.a(G822), .O(gate291inter7));
  inv1  gate2095(.a(G823), .O(gate291inter8));
  nand2 gate2096(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2097(.a(s_221), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2098(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2099(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2100(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2171(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2172(.a(gate296inter0), .b(s_232), .O(gate296inter1));
  and2  gate2173(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2174(.a(s_232), .O(gate296inter3));
  inv1  gate2175(.a(s_233), .O(gate296inter4));
  nand2 gate2176(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2177(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2178(.a(G826), .O(gate296inter7));
  inv1  gate2179(.a(G827), .O(gate296inter8));
  nand2 gate2180(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2181(.a(s_233), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2182(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2183(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2184(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1989(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1990(.a(gate393inter0), .b(s_206), .O(gate393inter1));
  and2  gate1991(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1992(.a(s_206), .O(gate393inter3));
  inv1  gate1993(.a(s_207), .O(gate393inter4));
  nand2 gate1994(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1995(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1996(.a(G7), .O(gate393inter7));
  inv1  gate1997(.a(G1054), .O(gate393inter8));
  nand2 gate1998(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1999(.a(s_207), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2000(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2001(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2002(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2283(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2284(.a(gate394inter0), .b(s_248), .O(gate394inter1));
  and2  gate2285(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2286(.a(s_248), .O(gate394inter3));
  inv1  gate2287(.a(s_249), .O(gate394inter4));
  nand2 gate2288(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2289(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2290(.a(G8), .O(gate394inter7));
  inv1  gate2291(.a(G1057), .O(gate394inter8));
  nand2 gate2292(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2293(.a(s_249), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2294(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2295(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2296(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2535(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2536(.a(gate397inter0), .b(s_284), .O(gate397inter1));
  and2  gate2537(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2538(.a(s_284), .O(gate397inter3));
  inv1  gate2539(.a(s_285), .O(gate397inter4));
  nand2 gate2540(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2541(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2542(.a(G11), .O(gate397inter7));
  inv1  gate2543(.a(G1066), .O(gate397inter8));
  nand2 gate2544(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2545(.a(s_285), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2546(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2547(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2548(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1037(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1038(.a(gate398inter0), .b(s_70), .O(gate398inter1));
  and2  gate1039(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1040(.a(s_70), .O(gate398inter3));
  inv1  gate1041(.a(s_71), .O(gate398inter4));
  nand2 gate1042(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1043(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1044(.a(G12), .O(gate398inter7));
  inv1  gate1045(.a(G1069), .O(gate398inter8));
  nand2 gate1046(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1047(.a(s_71), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1048(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1049(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1050(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1835(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1836(.a(gate400inter0), .b(s_184), .O(gate400inter1));
  and2  gate1837(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1838(.a(s_184), .O(gate400inter3));
  inv1  gate1839(.a(s_185), .O(gate400inter4));
  nand2 gate1840(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1841(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1842(.a(G14), .O(gate400inter7));
  inv1  gate1843(.a(G1075), .O(gate400inter8));
  nand2 gate1844(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1845(.a(s_185), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1846(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1847(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1848(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2423(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2424(.a(gate401inter0), .b(s_268), .O(gate401inter1));
  and2  gate2425(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2426(.a(s_268), .O(gate401inter3));
  inv1  gate2427(.a(s_269), .O(gate401inter4));
  nand2 gate2428(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2429(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2430(.a(G15), .O(gate401inter7));
  inv1  gate2431(.a(G1078), .O(gate401inter8));
  nand2 gate2432(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2433(.a(s_269), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2434(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2435(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2436(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1625(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1626(.a(gate403inter0), .b(s_154), .O(gate403inter1));
  and2  gate1627(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1628(.a(s_154), .O(gate403inter3));
  inv1  gate1629(.a(s_155), .O(gate403inter4));
  nand2 gate1630(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1631(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1632(.a(G17), .O(gate403inter7));
  inv1  gate1633(.a(G1084), .O(gate403inter8));
  nand2 gate1634(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1635(.a(s_155), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1636(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1637(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1638(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate575(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate576(.a(gate404inter0), .b(s_4), .O(gate404inter1));
  and2  gate577(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate578(.a(s_4), .O(gate404inter3));
  inv1  gate579(.a(s_5), .O(gate404inter4));
  nand2 gate580(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate581(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate582(.a(G18), .O(gate404inter7));
  inv1  gate583(.a(G1087), .O(gate404inter8));
  nand2 gate584(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate585(.a(s_5), .b(gate404inter3), .O(gate404inter10));
  nor2  gate586(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate587(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate588(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1009(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1010(.a(gate405inter0), .b(s_66), .O(gate405inter1));
  and2  gate1011(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1012(.a(s_66), .O(gate405inter3));
  inv1  gate1013(.a(s_67), .O(gate405inter4));
  nand2 gate1014(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1015(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1016(.a(G19), .O(gate405inter7));
  inv1  gate1017(.a(G1090), .O(gate405inter8));
  nand2 gate1018(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1019(.a(s_67), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1020(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1021(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1022(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate2549(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2550(.a(gate409inter0), .b(s_286), .O(gate409inter1));
  and2  gate2551(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2552(.a(s_286), .O(gate409inter3));
  inv1  gate2553(.a(s_287), .O(gate409inter4));
  nand2 gate2554(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2555(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2556(.a(G23), .O(gate409inter7));
  inv1  gate2557(.a(G1102), .O(gate409inter8));
  nand2 gate2558(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2559(.a(s_287), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2560(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2561(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2562(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate967(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate968(.a(gate410inter0), .b(s_60), .O(gate410inter1));
  and2  gate969(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate970(.a(s_60), .O(gate410inter3));
  inv1  gate971(.a(s_61), .O(gate410inter4));
  nand2 gate972(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate973(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate974(.a(G24), .O(gate410inter7));
  inv1  gate975(.a(G1105), .O(gate410inter8));
  nand2 gate976(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate977(.a(s_61), .b(gate410inter3), .O(gate410inter10));
  nor2  gate978(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate979(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate980(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate2003(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2004(.a(gate414inter0), .b(s_208), .O(gate414inter1));
  and2  gate2005(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2006(.a(s_208), .O(gate414inter3));
  inv1  gate2007(.a(s_209), .O(gate414inter4));
  nand2 gate2008(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2009(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2010(.a(G28), .O(gate414inter7));
  inv1  gate2011(.a(G1117), .O(gate414inter8));
  nand2 gate2012(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2013(.a(s_209), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2014(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2015(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2016(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate813(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate814(.a(gate418inter0), .b(s_38), .O(gate418inter1));
  and2  gate815(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate816(.a(s_38), .O(gate418inter3));
  inv1  gate817(.a(s_39), .O(gate418inter4));
  nand2 gate818(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate819(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate820(.a(G32), .O(gate418inter7));
  inv1  gate821(.a(G1129), .O(gate418inter8));
  nand2 gate822(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate823(.a(s_39), .b(gate418inter3), .O(gate418inter10));
  nor2  gate824(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate825(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate826(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2157(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2158(.a(gate419inter0), .b(s_230), .O(gate419inter1));
  and2  gate2159(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2160(.a(s_230), .O(gate419inter3));
  inv1  gate2161(.a(s_231), .O(gate419inter4));
  nand2 gate2162(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2163(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2164(.a(G1), .O(gate419inter7));
  inv1  gate2165(.a(G1132), .O(gate419inter8));
  nand2 gate2166(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2167(.a(s_231), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2168(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2169(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2170(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1023(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1024(.a(gate421inter0), .b(s_68), .O(gate421inter1));
  and2  gate1025(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1026(.a(s_68), .O(gate421inter3));
  inv1  gate1027(.a(s_69), .O(gate421inter4));
  nand2 gate1028(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1029(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1030(.a(G2), .O(gate421inter7));
  inv1  gate1031(.a(G1135), .O(gate421inter8));
  nand2 gate1032(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1033(.a(s_69), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1034(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1035(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1036(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2325(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2326(.a(gate422inter0), .b(s_254), .O(gate422inter1));
  and2  gate2327(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2328(.a(s_254), .O(gate422inter3));
  inv1  gate2329(.a(s_255), .O(gate422inter4));
  nand2 gate2330(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2331(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2332(.a(G1039), .O(gate422inter7));
  inv1  gate2333(.a(G1135), .O(gate422inter8));
  nand2 gate2334(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2335(.a(s_255), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2336(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2337(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2338(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1261(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1262(.a(gate425inter0), .b(s_102), .O(gate425inter1));
  and2  gate1263(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1264(.a(s_102), .O(gate425inter3));
  inv1  gate1265(.a(s_103), .O(gate425inter4));
  nand2 gate1266(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1267(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1268(.a(G4), .O(gate425inter7));
  inv1  gate1269(.a(G1141), .O(gate425inter8));
  nand2 gate1270(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1271(.a(s_103), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1272(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1273(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1274(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1387(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1388(.a(gate426inter0), .b(s_120), .O(gate426inter1));
  and2  gate1389(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1390(.a(s_120), .O(gate426inter3));
  inv1  gate1391(.a(s_121), .O(gate426inter4));
  nand2 gate1392(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1393(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1394(.a(G1045), .O(gate426inter7));
  inv1  gate1395(.a(G1141), .O(gate426inter8));
  nand2 gate1396(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1397(.a(s_121), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1398(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1399(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1400(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1317(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1318(.a(gate428inter0), .b(s_110), .O(gate428inter1));
  and2  gate1319(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1320(.a(s_110), .O(gate428inter3));
  inv1  gate1321(.a(s_111), .O(gate428inter4));
  nand2 gate1322(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1323(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1324(.a(G1048), .O(gate428inter7));
  inv1  gate1325(.a(G1144), .O(gate428inter8));
  nand2 gate1326(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1327(.a(s_111), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1328(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1329(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1330(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1681(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1682(.a(gate432inter0), .b(s_162), .O(gate432inter1));
  and2  gate1683(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1684(.a(s_162), .O(gate432inter3));
  inv1  gate1685(.a(s_163), .O(gate432inter4));
  nand2 gate1686(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1687(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1688(.a(G1054), .O(gate432inter7));
  inv1  gate1689(.a(G1150), .O(gate432inter8));
  nand2 gate1690(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1691(.a(s_163), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1692(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1693(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1694(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2269(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2270(.a(gate433inter0), .b(s_246), .O(gate433inter1));
  and2  gate2271(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2272(.a(s_246), .O(gate433inter3));
  inv1  gate2273(.a(s_247), .O(gate433inter4));
  nand2 gate2274(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2275(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2276(.a(G8), .O(gate433inter7));
  inv1  gate2277(.a(G1153), .O(gate433inter8));
  nand2 gate2278(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2279(.a(s_247), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2280(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2281(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2282(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1765(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1766(.a(gate436inter0), .b(s_174), .O(gate436inter1));
  and2  gate1767(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1768(.a(s_174), .O(gate436inter3));
  inv1  gate1769(.a(s_175), .O(gate436inter4));
  nand2 gate1770(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1771(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1772(.a(G1060), .O(gate436inter7));
  inv1  gate1773(.a(G1156), .O(gate436inter8));
  nand2 gate1774(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1775(.a(s_175), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1776(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1777(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1778(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1513(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1514(.a(gate439inter0), .b(s_138), .O(gate439inter1));
  and2  gate1515(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1516(.a(s_138), .O(gate439inter3));
  inv1  gate1517(.a(s_139), .O(gate439inter4));
  nand2 gate1518(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1519(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1520(.a(G11), .O(gate439inter7));
  inv1  gate1521(.a(G1162), .O(gate439inter8));
  nand2 gate1522(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1523(.a(s_139), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1524(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1525(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1526(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1611(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1612(.a(gate440inter0), .b(s_152), .O(gate440inter1));
  and2  gate1613(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1614(.a(s_152), .O(gate440inter3));
  inv1  gate1615(.a(s_153), .O(gate440inter4));
  nand2 gate1616(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1617(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1618(.a(G1066), .O(gate440inter7));
  inv1  gate1619(.a(G1162), .O(gate440inter8));
  nand2 gate1620(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1621(.a(s_153), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1622(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1623(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1624(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1247(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1248(.a(gate441inter0), .b(s_100), .O(gate441inter1));
  and2  gate1249(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1250(.a(s_100), .O(gate441inter3));
  inv1  gate1251(.a(s_101), .O(gate441inter4));
  nand2 gate1252(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1253(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1254(.a(G12), .O(gate441inter7));
  inv1  gate1255(.a(G1165), .O(gate441inter8));
  nand2 gate1256(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1257(.a(s_101), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1258(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1259(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1260(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2521(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2522(.a(gate444inter0), .b(s_282), .O(gate444inter1));
  and2  gate2523(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2524(.a(s_282), .O(gate444inter3));
  inv1  gate2525(.a(s_283), .O(gate444inter4));
  nand2 gate2526(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2527(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2528(.a(G1072), .O(gate444inter7));
  inv1  gate2529(.a(G1168), .O(gate444inter8));
  nand2 gate2530(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2531(.a(s_283), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2532(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2533(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2534(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate2241(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2242(.a(gate445inter0), .b(s_242), .O(gate445inter1));
  and2  gate2243(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2244(.a(s_242), .O(gate445inter3));
  inv1  gate2245(.a(s_243), .O(gate445inter4));
  nand2 gate2246(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2247(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2248(.a(G14), .O(gate445inter7));
  inv1  gate2249(.a(G1171), .O(gate445inter8));
  nand2 gate2250(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2251(.a(s_243), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2252(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2253(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2254(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate2045(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2046(.a(gate446inter0), .b(s_214), .O(gate446inter1));
  and2  gate2047(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2048(.a(s_214), .O(gate446inter3));
  inv1  gate2049(.a(s_215), .O(gate446inter4));
  nand2 gate2050(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2051(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2052(.a(G1075), .O(gate446inter7));
  inv1  gate2053(.a(G1171), .O(gate446inter8));
  nand2 gate2054(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2055(.a(s_215), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2056(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2057(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2058(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1639(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1640(.a(gate447inter0), .b(s_156), .O(gate447inter1));
  and2  gate1641(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1642(.a(s_156), .O(gate447inter3));
  inv1  gate1643(.a(s_157), .O(gate447inter4));
  nand2 gate1644(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1645(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1646(.a(G15), .O(gate447inter7));
  inv1  gate1647(.a(G1174), .O(gate447inter8));
  nand2 gate1648(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1649(.a(s_157), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1650(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1651(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1652(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate897(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate898(.a(gate448inter0), .b(s_50), .O(gate448inter1));
  and2  gate899(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate900(.a(s_50), .O(gate448inter3));
  inv1  gate901(.a(s_51), .O(gate448inter4));
  nand2 gate902(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate903(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate904(.a(G1078), .O(gate448inter7));
  inv1  gate905(.a(G1174), .O(gate448inter8));
  nand2 gate906(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate907(.a(s_51), .b(gate448inter3), .O(gate448inter10));
  nor2  gate908(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate909(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate910(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1065(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1066(.a(gate449inter0), .b(s_74), .O(gate449inter1));
  and2  gate1067(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1068(.a(s_74), .O(gate449inter3));
  inv1  gate1069(.a(s_75), .O(gate449inter4));
  nand2 gate1070(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1071(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1072(.a(G16), .O(gate449inter7));
  inv1  gate1073(.a(G1177), .O(gate449inter8));
  nand2 gate1074(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1075(.a(s_75), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1076(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1077(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1078(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate911(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate912(.a(gate453inter0), .b(s_52), .O(gate453inter1));
  and2  gate913(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate914(.a(s_52), .O(gate453inter3));
  inv1  gate915(.a(s_53), .O(gate453inter4));
  nand2 gate916(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate917(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate918(.a(G18), .O(gate453inter7));
  inv1  gate919(.a(G1183), .O(gate453inter8));
  nand2 gate920(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate921(.a(s_53), .b(gate453inter3), .O(gate453inter10));
  nor2  gate922(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate923(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate924(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2493(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2494(.a(gate455inter0), .b(s_278), .O(gate455inter1));
  and2  gate2495(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2496(.a(s_278), .O(gate455inter3));
  inv1  gate2497(.a(s_279), .O(gate455inter4));
  nand2 gate2498(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2499(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2500(.a(G19), .O(gate455inter7));
  inv1  gate2501(.a(G1186), .O(gate455inter8));
  nand2 gate2502(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2503(.a(s_279), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2504(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2505(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2506(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2199(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2200(.a(gate457inter0), .b(s_236), .O(gate457inter1));
  and2  gate2201(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2202(.a(s_236), .O(gate457inter3));
  inv1  gate2203(.a(s_237), .O(gate457inter4));
  nand2 gate2204(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2205(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2206(.a(G20), .O(gate457inter7));
  inv1  gate2207(.a(G1189), .O(gate457inter8));
  nand2 gate2208(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2209(.a(s_237), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2210(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2211(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2212(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2409(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2410(.a(gate459inter0), .b(s_266), .O(gate459inter1));
  and2  gate2411(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2412(.a(s_266), .O(gate459inter3));
  inv1  gate2413(.a(s_267), .O(gate459inter4));
  nand2 gate2414(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2415(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2416(.a(G21), .O(gate459inter7));
  inv1  gate2417(.a(G1192), .O(gate459inter8));
  nand2 gate2418(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2419(.a(s_267), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2420(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2421(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2422(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2129(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2130(.a(gate461inter0), .b(s_226), .O(gate461inter1));
  and2  gate2131(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2132(.a(s_226), .O(gate461inter3));
  inv1  gate2133(.a(s_227), .O(gate461inter4));
  nand2 gate2134(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2135(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2136(.a(G22), .O(gate461inter7));
  inv1  gate2137(.a(G1195), .O(gate461inter8));
  nand2 gate2138(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2139(.a(s_227), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2140(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2141(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2142(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate743(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate744(.a(gate462inter0), .b(s_28), .O(gate462inter1));
  and2  gate745(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate746(.a(s_28), .O(gate462inter3));
  inv1  gate747(.a(s_29), .O(gate462inter4));
  nand2 gate748(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate749(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate750(.a(G1099), .O(gate462inter7));
  inv1  gate751(.a(G1195), .O(gate462inter8));
  nand2 gate752(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate753(.a(s_29), .b(gate462inter3), .O(gate462inter10));
  nor2  gate754(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate755(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate756(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2507(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2508(.a(gate466inter0), .b(s_280), .O(gate466inter1));
  and2  gate2509(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2510(.a(s_280), .O(gate466inter3));
  inv1  gate2511(.a(s_281), .O(gate466inter4));
  nand2 gate2512(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2513(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2514(.a(G1105), .O(gate466inter7));
  inv1  gate2515(.a(G1201), .O(gate466inter8));
  nand2 gate2516(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2517(.a(s_281), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2518(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2519(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2520(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate771(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate772(.a(gate467inter0), .b(s_32), .O(gate467inter1));
  and2  gate773(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate774(.a(s_32), .O(gate467inter3));
  inv1  gate775(.a(s_33), .O(gate467inter4));
  nand2 gate776(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate777(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate778(.a(G25), .O(gate467inter7));
  inv1  gate779(.a(G1204), .O(gate467inter8));
  nand2 gate780(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate781(.a(s_33), .b(gate467inter3), .O(gate467inter10));
  nor2  gate782(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate783(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate784(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate687(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate688(.a(gate468inter0), .b(s_20), .O(gate468inter1));
  and2  gate689(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate690(.a(s_20), .O(gate468inter3));
  inv1  gate691(.a(s_21), .O(gate468inter4));
  nand2 gate692(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate693(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate694(.a(G1108), .O(gate468inter7));
  inv1  gate695(.a(G1204), .O(gate468inter8));
  nand2 gate696(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate697(.a(s_21), .b(gate468inter3), .O(gate468inter10));
  nor2  gate698(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate699(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate700(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate715(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate716(.a(gate471inter0), .b(s_24), .O(gate471inter1));
  and2  gate717(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate718(.a(s_24), .O(gate471inter3));
  inv1  gate719(.a(s_25), .O(gate471inter4));
  nand2 gate720(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate721(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate722(.a(G27), .O(gate471inter7));
  inv1  gate723(.a(G1210), .O(gate471inter8));
  nand2 gate724(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate725(.a(s_25), .b(gate471inter3), .O(gate471inter10));
  nor2  gate726(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate727(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate728(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2031(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2032(.a(gate475inter0), .b(s_212), .O(gate475inter1));
  and2  gate2033(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2034(.a(s_212), .O(gate475inter3));
  inv1  gate2035(.a(s_213), .O(gate475inter4));
  nand2 gate2036(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2037(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2038(.a(G29), .O(gate475inter7));
  inv1  gate2039(.a(G1216), .O(gate475inter8));
  nand2 gate2040(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2041(.a(s_213), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2042(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2043(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2044(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate925(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate926(.a(gate476inter0), .b(s_54), .O(gate476inter1));
  and2  gate927(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate928(.a(s_54), .O(gate476inter3));
  inv1  gate929(.a(s_55), .O(gate476inter4));
  nand2 gate930(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate931(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate932(.a(G1120), .O(gate476inter7));
  inv1  gate933(.a(G1216), .O(gate476inter8));
  nand2 gate934(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate935(.a(s_55), .b(gate476inter3), .O(gate476inter10));
  nor2  gate936(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate937(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate938(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1667(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1668(.a(gate486inter0), .b(s_160), .O(gate486inter1));
  and2  gate1669(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1670(.a(s_160), .O(gate486inter3));
  inv1  gate1671(.a(s_161), .O(gate486inter4));
  nand2 gate1672(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1673(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1674(.a(G1234), .O(gate486inter7));
  inv1  gate1675(.a(G1235), .O(gate486inter8));
  nand2 gate1676(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1677(.a(s_161), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1678(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1679(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1680(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2297(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2298(.a(gate489inter0), .b(s_250), .O(gate489inter1));
  and2  gate2299(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2300(.a(s_250), .O(gate489inter3));
  inv1  gate2301(.a(s_251), .O(gate489inter4));
  nand2 gate2302(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2303(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2304(.a(G1240), .O(gate489inter7));
  inv1  gate2305(.a(G1241), .O(gate489inter8));
  nand2 gate2306(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2307(.a(s_251), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2308(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2309(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2310(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1807(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1808(.a(gate492inter0), .b(s_180), .O(gate492inter1));
  and2  gate1809(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1810(.a(s_180), .O(gate492inter3));
  inv1  gate1811(.a(s_181), .O(gate492inter4));
  nand2 gate1812(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1813(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1814(.a(G1246), .O(gate492inter7));
  inv1  gate1815(.a(G1247), .O(gate492inter8));
  nand2 gate1816(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1817(.a(s_181), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1818(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1819(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1820(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1373(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1374(.a(gate497inter0), .b(s_118), .O(gate497inter1));
  and2  gate1375(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1376(.a(s_118), .O(gate497inter3));
  inv1  gate1377(.a(s_119), .O(gate497inter4));
  nand2 gate1378(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1379(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1380(.a(G1256), .O(gate497inter7));
  inv1  gate1381(.a(G1257), .O(gate497inter8));
  nand2 gate1382(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1383(.a(s_119), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1384(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1385(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1386(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1541(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1542(.a(gate499inter0), .b(s_142), .O(gate499inter1));
  and2  gate1543(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1544(.a(s_142), .O(gate499inter3));
  inv1  gate1545(.a(s_143), .O(gate499inter4));
  nand2 gate1546(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1547(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1548(.a(G1260), .O(gate499inter7));
  inv1  gate1549(.a(G1261), .O(gate499inter8));
  nand2 gate1550(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1551(.a(s_143), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1552(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1553(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1554(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2633(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2634(.a(gate508inter0), .b(s_298), .O(gate508inter1));
  and2  gate2635(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2636(.a(s_298), .O(gate508inter3));
  inv1  gate2637(.a(s_299), .O(gate508inter4));
  nand2 gate2638(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2639(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2640(.a(G1278), .O(gate508inter7));
  inv1  gate2641(.a(G1279), .O(gate508inter8));
  nand2 gate2642(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2643(.a(s_299), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2644(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2645(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2646(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate841(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate842(.a(gate510inter0), .b(s_42), .O(gate510inter1));
  and2  gate843(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate844(.a(s_42), .O(gate510inter3));
  inv1  gate845(.a(s_43), .O(gate510inter4));
  nand2 gate846(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate847(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate848(.a(G1282), .O(gate510inter7));
  inv1  gate849(.a(G1283), .O(gate510inter8));
  nand2 gate850(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate851(.a(s_43), .b(gate510inter3), .O(gate510inter10));
  nor2  gate852(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate853(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate854(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate603(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate604(.a(gate511inter0), .b(s_8), .O(gate511inter1));
  and2  gate605(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate606(.a(s_8), .O(gate511inter3));
  inv1  gate607(.a(s_9), .O(gate511inter4));
  nand2 gate608(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate609(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate610(.a(G1284), .O(gate511inter7));
  inv1  gate611(.a(G1285), .O(gate511inter8));
  nand2 gate612(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate613(.a(s_9), .b(gate511inter3), .O(gate511inter10));
  nor2  gate614(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate615(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate616(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1555(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1556(.a(gate514inter0), .b(s_144), .O(gate514inter1));
  and2  gate1557(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1558(.a(s_144), .O(gate514inter3));
  inv1  gate1559(.a(s_145), .O(gate514inter4));
  nand2 gate1560(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1561(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1562(.a(G1290), .O(gate514inter7));
  inv1  gate1563(.a(G1291), .O(gate514inter8));
  nand2 gate1564(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1565(.a(s_145), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1566(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1567(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1568(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule