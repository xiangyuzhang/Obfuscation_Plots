module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1695(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1696(.a(gate10inter0), .b(s_164), .O(gate10inter1));
  and2  gate1697(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1698(.a(s_164), .O(gate10inter3));
  inv1  gate1699(.a(s_165), .O(gate10inter4));
  nand2 gate1700(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1701(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1702(.a(G3), .O(gate10inter7));
  inv1  gate1703(.a(G4), .O(gate10inter8));
  nand2 gate1704(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1705(.a(s_165), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1706(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1707(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1708(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate2605(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2606(.a(gate21inter0), .b(s_294), .O(gate21inter1));
  and2  gate2607(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2608(.a(s_294), .O(gate21inter3));
  inv1  gate2609(.a(s_295), .O(gate21inter4));
  nand2 gate2610(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2611(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2612(.a(G25), .O(gate21inter7));
  inv1  gate2613(.a(G26), .O(gate21inter8));
  nand2 gate2614(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2615(.a(s_295), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2616(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2617(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2618(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2003(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2004(.a(gate22inter0), .b(s_208), .O(gate22inter1));
  and2  gate2005(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2006(.a(s_208), .O(gate22inter3));
  inv1  gate2007(.a(s_209), .O(gate22inter4));
  nand2 gate2008(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2009(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2010(.a(G27), .O(gate22inter7));
  inv1  gate2011(.a(G28), .O(gate22inter8));
  nand2 gate2012(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2013(.a(s_209), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2014(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2015(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2016(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1975(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1976(.a(gate23inter0), .b(s_204), .O(gate23inter1));
  and2  gate1977(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1978(.a(s_204), .O(gate23inter3));
  inv1  gate1979(.a(s_205), .O(gate23inter4));
  nand2 gate1980(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1981(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1982(.a(G29), .O(gate23inter7));
  inv1  gate1983(.a(G30), .O(gate23inter8));
  nand2 gate1984(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1985(.a(s_205), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1986(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1987(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1988(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1541(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1542(.a(gate28inter0), .b(s_142), .O(gate28inter1));
  and2  gate1543(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1544(.a(s_142), .O(gate28inter3));
  inv1  gate1545(.a(s_143), .O(gate28inter4));
  nand2 gate1546(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1547(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1548(.a(G10), .O(gate28inter7));
  inv1  gate1549(.a(G14), .O(gate28inter8));
  nand2 gate1550(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1551(.a(s_143), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1552(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1553(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1554(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1149(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1150(.a(gate31inter0), .b(s_86), .O(gate31inter1));
  and2  gate1151(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1152(.a(s_86), .O(gate31inter3));
  inv1  gate1153(.a(s_87), .O(gate31inter4));
  nand2 gate1154(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1155(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1156(.a(G4), .O(gate31inter7));
  inv1  gate1157(.a(G8), .O(gate31inter8));
  nand2 gate1158(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1159(.a(s_87), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1160(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1161(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1162(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2213(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2214(.a(gate38inter0), .b(s_238), .O(gate38inter1));
  and2  gate2215(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2216(.a(s_238), .O(gate38inter3));
  inv1  gate2217(.a(s_239), .O(gate38inter4));
  nand2 gate2218(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2219(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2220(.a(G27), .O(gate38inter7));
  inv1  gate2221(.a(G31), .O(gate38inter8));
  nand2 gate2222(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2223(.a(s_239), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2224(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2225(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2226(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2129(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2130(.a(gate40inter0), .b(s_226), .O(gate40inter1));
  and2  gate2131(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2132(.a(s_226), .O(gate40inter3));
  inv1  gate2133(.a(s_227), .O(gate40inter4));
  nand2 gate2134(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2135(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2136(.a(G28), .O(gate40inter7));
  inv1  gate2137(.a(G32), .O(gate40inter8));
  nand2 gate2138(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2139(.a(s_227), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2140(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2141(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2142(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate953(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate954(.a(gate45inter0), .b(s_58), .O(gate45inter1));
  and2  gate955(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate956(.a(s_58), .O(gate45inter3));
  inv1  gate957(.a(s_59), .O(gate45inter4));
  nand2 gate958(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate959(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate960(.a(G5), .O(gate45inter7));
  inv1  gate961(.a(G272), .O(gate45inter8));
  nand2 gate962(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate963(.a(s_59), .b(gate45inter3), .O(gate45inter10));
  nor2  gate964(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate965(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate966(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1107(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1108(.a(gate46inter0), .b(s_80), .O(gate46inter1));
  and2  gate1109(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1110(.a(s_80), .O(gate46inter3));
  inv1  gate1111(.a(s_81), .O(gate46inter4));
  nand2 gate1112(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1113(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1114(.a(G6), .O(gate46inter7));
  inv1  gate1115(.a(G272), .O(gate46inter8));
  nand2 gate1116(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1117(.a(s_81), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1118(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1119(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1120(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1863(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1864(.a(gate50inter0), .b(s_188), .O(gate50inter1));
  and2  gate1865(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1866(.a(s_188), .O(gate50inter3));
  inv1  gate1867(.a(s_189), .O(gate50inter4));
  nand2 gate1868(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1869(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1870(.a(G10), .O(gate50inter7));
  inv1  gate1871(.a(G278), .O(gate50inter8));
  nand2 gate1872(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1873(.a(s_189), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1874(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1875(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1876(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2269(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2270(.a(gate51inter0), .b(s_246), .O(gate51inter1));
  and2  gate2271(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2272(.a(s_246), .O(gate51inter3));
  inv1  gate2273(.a(s_247), .O(gate51inter4));
  nand2 gate2274(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2275(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2276(.a(G11), .O(gate51inter7));
  inv1  gate2277(.a(G281), .O(gate51inter8));
  nand2 gate2278(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2279(.a(s_247), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2280(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2281(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2282(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1499(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1500(.a(gate52inter0), .b(s_136), .O(gate52inter1));
  and2  gate1501(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1502(.a(s_136), .O(gate52inter3));
  inv1  gate1503(.a(s_137), .O(gate52inter4));
  nand2 gate1504(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1505(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1506(.a(G12), .O(gate52inter7));
  inv1  gate1507(.a(G281), .O(gate52inter8));
  nand2 gate1508(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1509(.a(s_137), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1510(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1511(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1512(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2759(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2760(.a(gate56inter0), .b(s_316), .O(gate56inter1));
  and2  gate2761(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2762(.a(s_316), .O(gate56inter3));
  inv1  gate2763(.a(s_317), .O(gate56inter4));
  nand2 gate2764(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2765(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2766(.a(G16), .O(gate56inter7));
  inv1  gate2767(.a(G287), .O(gate56inter8));
  nand2 gate2768(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2769(.a(s_317), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2770(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2771(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2772(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate841(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate842(.a(gate58inter0), .b(s_42), .O(gate58inter1));
  and2  gate843(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate844(.a(s_42), .O(gate58inter3));
  inv1  gate845(.a(s_43), .O(gate58inter4));
  nand2 gate846(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate847(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate848(.a(G18), .O(gate58inter7));
  inv1  gate849(.a(G290), .O(gate58inter8));
  nand2 gate850(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate851(.a(s_43), .b(gate58inter3), .O(gate58inter10));
  nor2  gate852(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate853(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate854(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1247(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1248(.a(gate59inter0), .b(s_100), .O(gate59inter1));
  and2  gate1249(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1250(.a(s_100), .O(gate59inter3));
  inv1  gate1251(.a(s_101), .O(gate59inter4));
  nand2 gate1252(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1253(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1254(.a(G19), .O(gate59inter7));
  inv1  gate1255(.a(G293), .O(gate59inter8));
  nand2 gate1256(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1257(.a(s_101), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1258(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1259(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1260(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1723(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1724(.a(gate60inter0), .b(s_168), .O(gate60inter1));
  and2  gate1725(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1726(.a(s_168), .O(gate60inter3));
  inv1  gate1727(.a(s_169), .O(gate60inter4));
  nand2 gate1728(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1729(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1730(.a(G20), .O(gate60inter7));
  inv1  gate1731(.a(G293), .O(gate60inter8));
  nand2 gate1732(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1733(.a(s_169), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1734(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1735(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1736(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate2857(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2858(.a(gate63inter0), .b(s_330), .O(gate63inter1));
  and2  gate2859(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2860(.a(s_330), .O(gate63inter3));
  inv1  gate2861(.a(s_331), .O(gate63inter4));
  nand2 gate2862(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2863(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2864(.a(G23), .O(gate63inter7));
  inv1  gate2865(.a(G299), .O(gate63inter8));
  nand2 gate2866(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2867(.a(s_331), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2868(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2869(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2870(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1877(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1878(.a(gate64inter0), .b(s_190), .O(gate64inter1));
  and2  gate1879(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1880(.a(s_190), .O(gate64inter3));
  inv1  gate1881(.a(s_191), .O(gate64inter4));
  nand2 gate1882(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1883(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1884(.a(G24), .O(gate64inter7));
  inv1  gate1885(.a(G299), .O(gate64inter8));
  nand2 gate1886(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1887(.a(s_191), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1888(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1889(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1890(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate939(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate940(.a(gate66inter0), .b(s_56), .O(gate66inter1));
  and2  gate941(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate942(.a(s_56), .O(gate66inter3));
  inv1  gate943(.a(s_57), .O(gate66inter4));
  nand2 gate944(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate945(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate946(.a(G26), .O(gate66inter7));
  inv1  gate947(.a(G302), .O(gate66inter8));
  nand2 gate948(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate949(.a(s_57), .b(gate66inter3), .O(gate66inter10));
  nor2  gate950(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate951(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate952(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1807(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1808(.a(gate72inter0), .b(s_180), .O(gate72inter1));
  and2  gate1809(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1810(.a(s_180), .O(gate72inter3));
  inv1  gate1811(.a(s_181), .O(gate72inter4));
  nand2 gate1812(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1813(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1814(.a(G32), .O(gate72inter7));
  inv1  gate1815(.a(G311), .O(gate72inter8));
  nand2 gate1816(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1817(.a(s_181), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1818(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1819(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1820(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate589(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate590(.a(gate73inter0), .b(s_6), .O(gate73inter1));
  and2  gate591(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate592(.a(s_6), .O(gate73inter3));
  inv1  gate593(.a(s_7), .O(gate73inter4));
  nand2 gate594(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate595(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate596(.a(G1), .O(gate73inter7));
  inv1  gate597(.a(G314), .O(gate73inter8));
  nand2 gate598(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate599(.a(s_7), .b(gate73inter3), .O(gate73inter10));
  nor2  gate600(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate601(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate602(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate967(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate968(.a(gate74inter0), .b(s_60), .O(gate74inter1));
  and2  gate969(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate970(.a(s_60), .O(gate74inter3));
  inv1  gate971(.a(s_61), .O(gate74inter4));
  nand2 gate972(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate973(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate974(.a(G5), .O(gate74inter7));
  inv1  gate975(.a(G314), .O(gate74inter8));
  nand2 gate976(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate977(.a(s_61), .b(gate74inter3), .O(gate74inter10));
  nor2  gate978(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate979(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate980(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate2087(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2088(.a(gate75inter0), .b(s_220), .O(gate75inter1));
  and2  gate2089(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2090(.a(s_220), .O(gate75inter3));
  inv1  gate2091(.a(s_221), .O(gate75inter4));
  nand2 gate2092(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2093(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2094(.a(G9), .O(gate75inter7));
  inv1  gate2095(.a(G317), .O(gate75inter8));
  nand2 gate2096(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2097(.a(s_221), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2098(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2099(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2100(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1891(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1892(.a(gate76inter0), .b(s_192), .O(gate76inter1));
  and2  gate1893(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1894(.a(s_192), .O(gate76inter3));
  inv1  gate1895(.a(s_193), .O(gate76inter4));
  nand2 gate1896(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1897(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1898(.a(G13), .O(gate76inter7));
  inv1  gate1899(.a(G317), .O(gate76inter8));
  nand2 gate1900(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1901(.a(s_193), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1902(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1903(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1904(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1989(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1990(.a(gate77inter0), .b(s_206), .O(gate77inter1));
  and2  gate1991(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1992(.a(s_206), .O(gate77inter3));
  inv1  gate1993(.a(s_207), .O(gate77inter4));
  nand2 gate1994(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1995(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1996(.a(G2), .O(gate77inter7));
  inv1  gate1997(.a(G320), .O(gate77inter8));
  nand2 gate1998(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1999(.a(s_207), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2000(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2001(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2002(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1065(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1066(.a(gate78inter0), .b(s_74), .O(gate78inter1));
  and2  gate1067(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1068(.a(s_74), .O(gate78inter3));
  inv1  gate1069(.a(s_75), .O(gate78inter4));
  nand2 gate1070(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1071(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1072(.a(G6), .O(gate78inter7));
  inv1  gate1073(.a(G320), .O(gate78inter8));
  nand2 gate1074(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1075(.a(s_75), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1076(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1077(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1078(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1597(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1598(.a(gate79inter0), .b(s_150), .O(gate79inter1));
  and2  gate1599(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1600(.a(s_150), .O(gate79inter3));
  inv1  gate1601(.a(s_151), .O(gate79inter4));
  nand2 gate1602(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1603(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1604(.a(G10), .O(gate79inter7));
  inv1  gate1605(.a(G323), .O(gate79inter8));
  nand2 gate1606(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1607(.a(s_151), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1608(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1609(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1610(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1093(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1094(.a(gate81inter0), .b(s_78), .O(gate81inter1));
  and2  gate1095(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1096(.a(s_78), .O(gate81inter3));
  inv1  gate1097(.a(s_79), .O(gate81inter4));
  nand2 gate1098(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1099(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1100(.a(G3), .O(gate81inter7));
  inv1  gate1101(.a(G326), .O(gate81inter8));
  nand2 gate1102(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1103(.a(s_79), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1104(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1105(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1106(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2073(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2074(.a(gate88inter0), .b(s_218), .O(gate88inter1));
  and2  gate2075(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2076(.a(s_218), .O(gate88inter3));
  inv1  gate2077(.a(s_219), .O(gate88inter4));
  nand2 gate2078(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2079(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2080(.a(G16), .O(gate88inter7));
  inv1  gate2081(.a(G335), .O(gate88inter8));
  nand2 gate2082(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2083(.a(s_219), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2084(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2085(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2086(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2507(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2508(.a(gate89inter0), .b(s_280), .O(gate89inter1));
  and2  gate2509(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2510(.a(s_280), .O(gate89inter3));
  inv1  gate2511(.a(s_281), .O(gate89inter4));
  nand2 gate2512(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2513(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2514(.a(G17), .O(gate89inter7));
  inv1  gate2515(.a(G338), .O(gate89inter8));
  nand2 gate2516(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2517(.a(s_281), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2518(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2519(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2520(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate687(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate688(.a(gate91inter0), .b(s_20), .O(gate91inter1));
  and2  gate689(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate690(.a(s_20), .O(gate91inter3));
  inv1  gate691(.a(s_21), .O(gate91inter4));
  nand2 gate692(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate693(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate694(.a(G25), .O(gate91inter7));
  inv1  gate695(.a(G341), .O(gate91inter8));
  nand2 gate696(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate697(.a(s_21), .b(gate91inter3), .O(gate91inter10));
  nor2  gate698(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate699(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate700(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate631(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate632(.a(gate92inter0), .b(s_12), .O(gate92inter1));
  and2  gate633(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate634(.a(s_12), .O(gate92inter3));
  inv1  gate635(.a(s_13), .O(gate92inter4));
  nand2 gate636(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate637(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate638(.a(G29), .O(gate92inter7));
  inv1  gate639(.a(G341), .O(gate92inter8));
  nand2 gate640(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate641(.a(s_13), .b(gate92inter3), .O(gate92inter10));
  nor2  gate642(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate643(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate644(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1387(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1388(.a(gate93inter0), .b(s_120), .O(gate93inter1));
  and2  gate1389(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1390(.a(s_120), .O(gate93inter3));
  inv1  gate1391(.a(s_121), .O(gate93inter4));
  nand2 gate1392(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1393(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1394(.a(G18), .O(gate93inter7));
  inv1  gate1395(.a(G344), .O(gate93inter8));
  nand2 gate1396(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1397(.a(s_121), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1398(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1399(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1400(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate575(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate576(.a(gate94inter0), .b(s_4), .O(gate94inter1));
  and2  gate577(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate578(.a(s_4), .O(gate94inter3));
  inv1  gate579(.a(s_5), .O(gate94inter4));
  nand2 gate580(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate581(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate582(.a(G22), .O(gate94inter7));
  inv1  gate583(.a(G344), .O(gate94inter8));
  nand2 gate584(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate585(.a(s_5), .b(gate94inter3), .O(gate94inter10));
  nor2  gate586(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate587(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate588(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2675(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2676(.a(gate97inter0), .b(s_304), .O(gate97inter1));
  and2  gate2677(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2678(.a(s_304), .O(gate97inter3));
  inv1  gate2679(.a(s_305), .O(gate97inter4));
  nand2 gate2680(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2681(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2682(.a(G19), .O(gate97inter7));
  inv1  gate2683(.a(G350), .O(gate97inter8));
  nand2 gate2684(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2685(.a(s_305), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2686(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2687(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2688(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1457(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1458(.a(gate98inter0), .b(s_130), .O(gate98inter1));
  and2  gate1459(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1460(.a(s_130), .O(gate98inter3));
  inv1  gate1461(.a(s_131), .O(gate98inter4));
  nand2 gate1462(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1463(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1464(.a(G23), .O(gate98inter7));
  inv1  gate1465(.a(G350), .O(gate98inter8));
  nand2 gate1466(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1467(.a(s_131), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1468(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1469(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1470(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1947(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1948(.a(gate99inter0), .b(s_200), .O(gate99inter1));
  and2  gate1949(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1950(.a(s_200), .O(gate99inter3));
  inv1  gate1951(.a(s_201), .O(gate99inter4));
  nand2 gate1952(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1953(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1954(.a(G27), .O(gate99inter7));
  inv1  gate1955(.a(G353), .O(gate99inter8));
  nand2 gate1956(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1957(.a(s_201), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1958(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1959(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1960(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate659(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate660(.a(gate107inter0), .b(s_16), .O(gate107inter1));
  and2  gate661(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate662(.a(s_16), .O(gate107inter3));
  inv1  gate663(.a(s_17), .O(gate107inter4));
  nand2 gate664(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate665(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate666(.a(G366), .O(gate107inter7));
  inv1  gate667(.a(G367), .O(gate107inter8));
  nand2 gate668(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate669(.a(s_17), .b(gate107inter3), .O(gate107inter10));
  nor2  gate670(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate671(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate672(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2829(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2830(.a(gate111inter0), .b(s_326), .O(gate111inter1));
  and2  gate2831(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2832(.a(s_326), .O(gate111inter3));
  inv1  gate2833(.a(s_327), .O(gate111inter4));
  nand2 gate2834(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2835(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2836(.a(G374), .O(gate111inter7));
  inv1  gate2837(.a(G375), .O(gate111inter8));
  nand2 gate2838(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2839(.a(s_327), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2840(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2841(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2842(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2339(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2340(.a(gate112inter0), .b(s_256), .O(gate112inter1));
  and2  gate2341(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2342(.a(s_256), .O(gate112inter3));
  inv1  gate2343(.a(s_257), .O(gate112inter4));
  nand2 gate2344(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2345(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2346(.a(G376), .O(gate112inter7));
  inv1  gate2347(.a(G377), .O(gate112inter8));
  nand2 gate2348(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2349(.a(s_257), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2350(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2351(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2352(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2059(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2060(.a(gate121inter0), .b(s_216), .O(gate121inter1));
  and2  gate2061(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2062(.a(s_216), .O(gate121inter3));
  inv1  gate2063(.a(s_217), .O(gate121inter4));
  nand2 gate2064(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2065(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2066(.a(G394), .O(gate121inter7));
  inv1  gate2067(.a(G395), .O(gate121inter8));
  nand2 gate2068(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2069(.a(s_217), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2070(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2071(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2072(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate729(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate730(.a(gate123inter0), .b(s_26), .O(gate123inter1));
  and2  gate731(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate732(.a(s_26), .O(gate123inter3));
  inv1  gate733(.a(s_27), .O(gate123inter4));
  nand2 gate734(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate735(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate736(.a(G398), .O(gate123inter7));
  inv1  gate737(.a(G399), .O(gate123inter8));
  nand2 gate738(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate739(.a(s_27), .b(gate123inter3), .O(gate123inter10));
  nor2  gate740(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate741(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate742(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1079(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1080(.a(gate124inter0), .b(s_76), .O(gate124inter1));
  and2  gate1081(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1082(.a(s_76), .O(gate124inter3));
  inv1  gate1083(.a(s_77), .O(gate124inter4));
  nand2 gate1084(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1085(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1086(.a(G400), .O(gate124inter7));
  inv1  gate1087(.a(G401), .O(gate124inter8));
  nand2 gate1088(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1089(.a(s_77), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1090(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1091(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1092(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2689(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2690(.a(gate131inter0), .b(s_306), .O(gate131inter1));
  and2  gate2691(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2692(.a(s_306), .O(gate131inter3));
  inv1  gate2693(.a(s_307), .O(gate131inter4));
  nand2 gate2694(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2695(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2696(.a(G414), .O(gate131inter7));
  inv1  gate2697(.a(G415), .O(gate131inter8));
  nand2 gate2698(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2699(.a(s_307), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2700(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2701(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2702(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate603(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate604(.a(gate135inter0), .b(s_8), .O(gate135inter1));
  and2  gate605(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate606(.a(s_8), .O(gate135inter3));
  inv1  gate607(.a(s_9), .O(gate135inter4));
  nand2 gate608(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate609(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate610(.a(G422), .O(gate135inter7));
  inv1  gate611(.a(G423), .O(gate135inter8));
  nand2 gate612(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate613(.a(s_9), .b(gate135inter3), .O(gate135inter10));
  nor2  gate614(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate615(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate616(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate785(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate786(.a(gate139inter0), .b(s_34), .O(gate139inter1));
  and2  gate787(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate788(.a(s_34), .O(gate139inter3));
  inv1  gate789(.a(s_35), .O(gate139inter4));
  nand2 gate790(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate791(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate792(.a(G438), .O(gate139inter7));
  inv1  gate793(.a(G441), .O(gate139inter8));
  nand2 gate794(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate795(.a(s_35), .b(gate139inter3), .O(gate139inter10));
  nor2  gate796(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate797(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate798(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate771(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate772(.a(gate140inter0), .b(s_32), .O(gate140inter1));
  and2  gate773(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate774(.a(s_32), .O(gate140inter3));
  inv1  gate775(.a(s_33), .O(gate140inter4));
  nand2 gate776(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate777(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate778(.a(G444), .O(gate140inter7));
  inv1  gate779(.a(G447), .O(gate140inter8));
  nand2 gate780(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate781(.a(s_33), .b(gate140inter3), .O(gate140inter10));
  nor2  gate782(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate783(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate784(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2745(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2746(.a(gate144inter0), .b(s_314), .O(gate144inter1));
  and2  gate2747(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2748(.a(s_314), .O(gate144inter3));
  inv1  gate2749(.a(s_315), .O(gate144inter4));
  nand2 gate2750(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2751(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2752(.a(G468), .O(gate144inter7));
  inv1  gate2753(.a(G471), .O(gate144inter8));
  nand2 gate2754(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2755(.a(s_315), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2756(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2757(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2758(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2591(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2592(.a(gate145inter0), .b(s_292), .O(gate145inter1));
  and2  gate2593(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2594(.a(s_292), .O(gate145inter3));
  inv1  gate2595(.a(s_293), .O(gate145inter4));
  nand2 gate2596(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2597(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2598(.a(G474), .O(gate145inter7));
  inv1  gate2599(.a(G477), .O(gate145inter8));
  nand2 gate2600(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2601(.a(s_293), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2602(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2603(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2604(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1289(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1290(.a(gate150inter0), .b(s_106), .O(gate150inter1));
  and2  gate1291(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1292(.a(s_106), .O(gate150inter3));
  inv1  gate1293(.a(s_107), .O(gate150inter4));
  nand2 gate1294(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1295(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1296(.a(G504), .O(gate150inter7));
  inv1  gate1297(.a(G507), .O(gate150inter8));
  nand2 gate1298(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1299(.a(s_107), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1300(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1301(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1302(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate855(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate856(.a(gate153inter0), .b(s_44), .O(gate153inter1));
  and2  gate857(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate858(.a(s_44), .O(gate153inter3));
  inv1  gate859(.a(s_45), .O(gate153inter4));
  nand2 gate860(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate861(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate862(.a(G426), .O(gate153inter7));
  inv1  gate863(.a(G522), .O(gate153inter8));
  nand2 gate864(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate865(.a(s_45), .b(gate153inter3), .O(gate153inter10));
  nor2  gate866(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate867(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate868(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate813(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate814(.a(gate154inter0), .b(s_38), .O(gate154inter1));
  and2  gate815(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate816(.a(s_38), .O(gate154inter3));
  inv1  gate817(.a(s_39), .O(gate154inter4));
  nand2 gate818(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate819(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate820(.a(G429), .O(gate154inter7));
  inv1  gate821(.a(G522), .O(gate154inter8));
  nand2 gate822(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate823(.a(s_39), .b(gate154inter3), .O(gate154inter10));
  nor2  gate824(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate825(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate826(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1933(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1934(.a(gate159inter0), .b(s_198), .O(gate159inter1));
  and2  gate1935(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1936(.a(s_198), .O(gate159inter3));
  inv1  gate1937(.a(s_199), .O(gate159inter4));
  nand2 gate1938(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1939(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1940(.a(G444), .O(gate159inter7));
  inv1  gate1941(.a(G531), .O(gate159inter8));
  nand2 gate1942(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1943(.a(s_199), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1944(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1945(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1946(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1121(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1122(.a(gate160inter0), .b(s_82), .O(gate160inter1));
  and2  gate1123(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1124(.a(s_82), .O(gate160inter3));
  inv1  gate1125(.a(s_83), .O(gate160inter4));
  nand2 gate1126(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1127(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1128(.a(G447), .O(gate160inter7));
  inv1  gate1129(.a(G531), .O(gate160inter8));
  nand2 gate1130(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1131(.a(s_83), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1132(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1133(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1134(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1331(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1332(.a(gate161inter0), .b(s_112), .O(gate161inter1));
  and2  gate1333(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1334(.a(s_112), .O(gate161inter3));
  inv1  gate1335(.a(s_113), .O(gate161inter4));
  nand2 gate1336(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1337(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1338(.a(G450), .O(gate161inter7));
  inv1  gate1339(.a(G534), .O(gate161inter8));
  nand2 gate1340(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1341(.a(s_113), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1342(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1343(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1344(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1737(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1738(.a(gate165inter0), .b(s_170), .O(gate165inter1));
  and2  gate1739(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1740(.a(s_170), .O(gate165inter3));
  inv1  gate1741(.a(s_171), .O(gate165inter4));
  nand2 gate1742(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1743(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1744(.a(G462), .O(gate165inter7));
  inv1  gate1745(.a(G540), .O(gate165inter8));
  nand2 gate1746(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1747(.a(s_171), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1748(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1749(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1750(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate743(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate744(.a(gate166inter0), .b(s_28), .O(gate166inter1));
  and2  gate745(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate746(.a(s_28), .O(gate166inter3));
  inv1  gate747(.a(s_29), .O(gate166inter4));
  nand2 gate748(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate749(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate750(.a(G465), .O(gate166inter7));
  inv1  gate751(.a(G540), .O(gate166inter8));
  nand2 gate752(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate753(.a(s_29), .b(gate166inter3), .O(gate166inter10));
  nor2  gate754(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate755(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate756(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1681(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1682(.a(gate167inter0), .b(s_162), .O(gate167inter1));
  and2  gate1683(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1684(.a(s_162), .O(gate167inter3));
  inv1  gate1685(.a(s_163), .O(gate167inter4));
  nand2 gate1686(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1687(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1688(.a(G468), .O(gate167inter7));
  inv1  gate1689(.a(G543), .O(gate167inter8));
  nand2 gate1690(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1691(.a(s_163), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1692(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1693(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1694(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1611(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1612(.a(gate169inter0), .b(s_152), .O(gate169inter1));
  and2  gate1613(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1614(.a(s_152), .O(gate169inter3));
  inv1  gate1615(.a(s_153), .O(gate169inter4));
  nand2 gate1616(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1617(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1618(.a(G474), .O(gate169inter7));
  inv1  gate1619(.a(G546), .O(gate169inter8));
  nand2 gate1620(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1621(.a(s_153), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1622(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1623(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1624(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1849(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1850(.a(gate173inter0), .b(s_186), .O(gate173inter1));
  and2  gate1851(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1852(.a(s_186), .O(gate173inter3));
  inv1  gate1853(.a(s_187), .O(gate173inter4));
  nand2 gate1854(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1855(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1856(.a(G486), .O(gate173inter7));
  inv1  gate1857(.a(G552), .O(gate173inter8));
  nand2 gate1858(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1859(.a(s_187), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1860(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1861(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1862(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2255(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2256(.a(gate175inter0), .b(s_244), .O(gate175inter1));
  and2  gate2257(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2258(.a(s_244), .O(gate175inter3));
  inv1  gate2259(.a(s_245), .O(gate175inter4));
  nand2 gate2260(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2261(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2262(.a(G492), .O(gate175inter7));
  inv1  gate2263(.a(G555), .O(gate175inter8));
  nand2 gate2264(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2265(.a(s_245), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2266(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2267(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2268(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1555(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1556(.a(gate176inter0), .b(s_144), .O(gate176inter1));
  and2  gate1557(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1558(.a(s_144), .O(gate176inter3));
  inv1  gate1559(.a(s_145), .O(gate176inter4));
  nand2 gate1560(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1561(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1562(.a(G495), .O(gate176inter7));
  inv1  gate1563(.a(G555), .O(gate176inter8));
  nand2 gate1564(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1565(.a(s_145), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1566(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1567(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1568(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate897(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate898(.a(gate177inter0), .b(s_50), .O(gate177inter1));
  and2  gate899(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate900(.a(s_50), .O(gate177inter3));
  inv1  gate901(.a(s_51), .O(gate177inter4));
  nand2 gate902(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate903(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate904(.a(G498), .O(gate177inter7));
  inv1  gate905(.a(G558), .O(gate177inter8));
  nand2 gate906(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate907(.a(s_51), .b(gate177inter3), .O(gate177inter10));
  nor2  gate908(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate909(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate910(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate799(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate800(.a(gate179inter0), .b(s_36), .O(gate179inter1));
  and2  gate801(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate802(.a(s_36), .O(gate179inter3));
  inv1  gate803(.a(s_37), .O(gate179inter4));
  nand2 gate804(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate805(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate806(.a(G504), .O(gate179inter7));
  inv1  gate807(.a(G561), .O(gate179inter8));
  nand2 gate808(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate809(.a(s_37), .b(gate179inter3), .O(gate179inter10));
  nor2  gate810(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate811(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate812(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1009(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1010(.a(gate181inter0), .b(s_66), .O(gate181inter1));
  and2  gate1011(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1012(.a(s_66), .O(gate181inter3));
  inv1  gate1013(.a(s_67), .O(gate181inter4));
  nand2 gate1014(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1015(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1016(.a(G510), .O(gate181inter7));
  inv1  gate1017(.a(G564), .O(gate181inter8));
  nand2 gate1018(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1019(.a(s_67), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1020(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1021(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1022(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2185(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2186(.a(gate182inter0), .b(s_234), .O(gate182inter1));
  and2  gate2187(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2188(.a(s_234), .O(gate182inter3));
  inv1  gate2189(.a(s_235), .O(gate182inter4));
  nand2 gate2190(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2191(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2192(.a(G513), .O(gate182inter7));
  inv1  gate2193(.a(G564), .O(gate182inter8));
  nand2 gate2194(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2195(.a(s_235), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2196(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2197(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2198(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate883(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate884(.a(gate183inter0), .b(s_48), .O(gate183inter1));
  and2  gate885(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate886(.a(s_48), .O(gate183inter3));
  inv1  gate887(.a(s_49), .O(gate183inter4));
  nand2 gate888(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate889(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate890(.a(G516), .O(gate183inter7));
  inv1  gate891(.a(G567), .O(gate183inter8));
  nand2 gate892(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate893(.a(s_49), .b(gate183inter3), .O(gate183inter10));
  nor2  gate894(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate895(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate896(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate2381(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2382(.a(gate186inter0), .b(s_262), .O(gate186inter1));
  and2  gate2383(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2384(.a(s_262), .O(gate186inter3));
  inv1  gate2385(.a(s_263), .O(gate186inter4));
  nand2 gate2386(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2387(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2388(.a(G572), .O(gate186inter7));
  inv1  gate2389(.a(G573), .O(gate186inter8));
  nand2 gate2390(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2391(.a(s_263), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2392(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2393(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2394(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate869(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate870(.a(gate189inter0), .b(s_46), .O(gate189inter1));
  and2  gate871(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate872(.a(s_46), .O(gate189inter3));
  inv1  gate873(.a(s_47), .O(gate189inter4));
  nand2 gate874(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate875(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate876(.a(G578), .O(gate189inter7));
  inv1  gate877(.a(G579), .O(gate189inter8));
  nand2 gate878(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate879(.a(s_47), .b(gate189inter3), .O(gate189inter10));
  nor2  gate880(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate881(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate882(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate995(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate996(.a(gate193inter0), .b(s_64), .O(gate193inter1));
  and2  gate997(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate998(.a(s_64), .O(gate193inter3));
  inv1  gate999(.a(s_65), .O(gate193inter4));
  nand2 gate1000(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1001(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1002(.a(G586), .O(gate193inter7));
  inv1  gate1003(.a(G587), .O(gate193inter8));
  nand2 gate1004(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1005(.a(s_65), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1006(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1007(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1008(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1485(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1486(.a(gate197inter0), .b(s_134), .O(gate197inter1));
  and2  gate1487(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1488(.a(s_134), .O(gate197inter3));
  inv1  gate1489(.a(s_135), .O(gate197inter4));
  nand2 gate1490(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1491(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1492(.a(G594), .O(gate197inter7));
  inv1  gate1493(.a(G595), .O(gate197inter8));
  nand2 gate1494(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1495(.a(s_135), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1496(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1497(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1498(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1625(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1626(.a(gate199inter0), .b(s_154), .O(gate199inter1));
  and2  gate1627(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1628(.a(s_154), .O(gate199inter3));
  inv1  gate1629(.a(s_155), .O(gate199inter4));
  nand2 gate1630(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1631(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1632(.a(G598), .O(gate199inter7));
  inv1  gate1633(.a(G599), .O(gate199inter8));
  nand2 gate1634(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1635(.a(s_155), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1636(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1637(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1638(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2199(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2200(.a(gate201inter0), .b(s_236), .O(gate201inter1));
  and2  gate2201(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2202(.a(s_236), .O(gate201inter3));
  inv1  gate2203(.a(s_237), .O(gate201inter4));
  nand2 gate2204(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2205(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2206(.a(G602), .O(gate201inter7));
  inv1  gate2207(.a(G607), .O(gate201inter8));
  nand2 gate2208(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2209(.a(s_237), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2210(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2211(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2212(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1023(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1024(.a(gate203inter0), .b(s_68), .O(gate203inter1));
  and2  gate1025(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1026(.a(s_68), .O(gate203inter3));
  inv1  gate1027(.a(s_69), .O(gate203inter4));
  nand2 gate1028(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1029(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1030(.a(G602), .O(gate203inter7));
  inv1  gate1031(.a(G612), .O(gate203inter8));
  nand2 gate1032(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1033(.a(s_69), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1034(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1035(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1036(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1051(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1052(.a(gate206inter0), .b(s_72), .O(gate206inter1));
  and2  gate1053(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1054(.a(s_72), .O(gate206inter3));
  inv1  gate1055(.a(s_73), .O(gate206inter4));
  nand2 gate1056(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1057(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1058(.a(G632), .O(gate206inter7));
  inv1  gate1059(.a(G637), .O(gate206inter8));
  nand2 gate1060(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1061(.a(s_73), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1062(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1063(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1064(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1443(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1444(.a(gate210inter0), .b(s_128), .O(gate210inter1));
  and2  gate1445(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1446(.a(s_128), .O(gate210inter3));
  inv1  gate1447(.a(s_129), .O(gate210inter4));
  nand2 gate1448(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1449(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1450(.a(G607), .O(gate210inter7));
  inv1  gate1451(.a(G666), .O(gate210inter8));
  nand2 gate1452(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1453(.a(s_129), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1454(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1455(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1456(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1345(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1346(.a(gate211inter0), .b(s_114), .O(gate211inter1));
  and2  gate1347(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1348(.a(s_114), .O(gate211inter3));
  inv1  gate1349(.a(s_115), .O(gate211inter4));
  nand2 gate1350(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1351(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1352(.a(G612), .O(gate211inter7));
  inv1  gate1353(.a(G669), .O(gate211inter8));
  nand2 gate1354(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1355(.a(s_115), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1356(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1357(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1358(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate911(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate912(.a(gate214inter0), .b(s_52), .O(gate214inter1));
  and2  gate913(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate914(.a(s_52), .O(gate214inter3));
  inv1  gate915(.a(s_53), .O(gate214inter4));
  nand2 gate916(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate917(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate918(.a(G612), .O(gate214inter7));
  inv1  gate919(.a(G672), .O(gate214inter8));
  nand2 gate920(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate921(.a(s_53), .b(gate214inter3), .O(gate214inter10));
  nor2  gate922(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate923(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate924(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1667(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1668(.a(gate215inter0), .b(s_160), .O(gate215inter1));
  and2  gate1669(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1670(.a(s_160), .O(gate215inter3));
  inv1  gate1671(.a(s_161), .O(gate215inter4));
  nand2 gate1672(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1673(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1674(.a(G607), .O(gate215inter7));
  inv1  gate1675(.a(G675), .O(gate215inter8));
  nand2 gate1676(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1677(.a(s_161), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1678(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1679(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1680(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2101(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2102(.a(gate217inter0), .b(s_222), .O(gate217inter1));
  and2  gate2103(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2104(.a(s_222), .O(gate217inter3));
  inv1  gate2105(.a(s_223), .O(gate217inter4));
  nand2 gate2106(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2107(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2108(.a(G622), .O(gate217inter7));
  inv1  gate2109(.a(G678), .O(gate217inter8));
  nand2 gate2110(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2111(.a(s_223), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2112(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2113(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2114(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate2549(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2550(.a(gate219inter0), .b(s_286), .O(gate219inter1));
  and2  gate2551(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2552(.a(s_286), .O(gate219inter3));
  inv1  gate2553(.a(s_287), .O(gate219inter4));
  nand2 gate2554(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2555(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2556(.a(G632), .O(gate219inter7));
  inv1  gate2557(.a(G681), .O(gate219inter8));
  nand2 gate2558(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2559(.a(s_287), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2560(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2561(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2562(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2717(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2718(.a(gate220inter0), .b(s_310), .O(gate220inter1));
  and2  gate2719(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2720(.a(s_310), .O(gate220inter3));
  inv1  gate2721(.a(s_311), .O(gate220inter4));
  nand2 gate2722(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2723(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2724(.a(G637), .O(gate220inter7));
  inv1  gate2725(.a(G681), .O(gate220inter8));
  nand2 gate2726(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2727(.a(s_311), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2728(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2729(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2730(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate2241(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate2242(.a(gate221inter0), .b(s_242), .O(gate221inter1));
  and2  gate2243(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate2244(.a(s_242), .O(gate221inter3));
  inv1  gate2245(.a(s_243), .O(gate221inter4));
  nand2 gate2246(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate2247(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate2248(.a(G622), .O(gate221inter7));
  inv1  gate2249(.a(G684), .O(gate221inter8));
  nand2 gate2250(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate2251(.a(s_243), .b(gate221inter3), .O(gate221inter10));
  nor2  gate2252(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate2253(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate2254(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1401(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1402(.a(gate222inter0), .b(s_122), .O(gate222inter1));
  and2  gate1403(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1404(.a(s_122), .O(gate222inter3));
  inv1  gate1405(.a(s_123), .O(gate222inter4));
  nand2 gate1406(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1407(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1408(.a(G632), .O(gate222inter7));
  inv1  gate1409(.a(G684), .O(gate222inter8));
  nand2 gate1410(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1411(.a(s_123), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1412(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1413(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1414(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2045(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2046(.a(gate224inter0), .b(s_214), .O(gate224inter1));
  and2  gate2047(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2048(.a(s_214), .O(gate224inter3));
  inv1  gate2049(.a(s_215), .O(gate224inter4));
  nand2 gate2050(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2051(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2052(.a(G637), .O(gate224inter7));
  inv1  gate2053(.a(G687), .O(gate224inter8));
  nand2 gate2054(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2055(.a(s_215), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2056(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2057(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2058(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1037(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1038(.a(gate226inter0), .b(s_70), .O(gate226inter1));
  and2  gate1039(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1040(.a(s_70), .O(gate226inter3));
  inv1  gate1041(.a(s_71), .O(gate226inter4));
  nand2 gate1042(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1043(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1044(.a(G692), .O(gate226inter7));
  inv1  gate1045(.a(G693), .O(gate226inter8));
  nand2 gate1046(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1047(.a(s_71), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1048(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1049(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1050(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate617(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate618(.a(gate227inter0), .b(s_10), .O(gate227inter1));
  and2  gate619(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate620(.a(s_10), .O(gate227inter3));
  inv1  gate621(.a(s_11), .O(gate227inter4));
  nand2 gate622(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate623(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate624(.a(G694), .O(gate227inter7));
  inv1  gate625(.a(G695), .O(gate227inter8));
  nand2 gate626(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate627(.a(s_11), .b(gate227inter3), .O(gate227inter10));
  nor2  gate628(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate629(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate630(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2353(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2354(.a(gate229inter0), .b(s_258), .O(gate229inter1));
  and2  gate2355(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2356(.a(s_258), .O(gate229inter3));
  inv1  gate2357(.a(s_259), .O(gate229inter4));
  nand2 gate2358(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2359(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2360(.a(G698), .O(gate229inter7));
  inv1  gate2361(.a(G699), .O(gate229inter8));
  nand2 gate2362(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2363(.a(s_259), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2364(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2365(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2366(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1233(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1234(.a(gate234inter0), .b(s_98), .O(gate234inter1));
  and2  gate1235(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1236(.a(s_98), .O(gate234inter3));
  inv1  gate1237(.a(s_99), .O(gate234inter4));
  nand2 gate1238(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1239(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1240(.a(G245), .O(gate234inter7));
  inv1  gate1241(.a(G721), .O(gate234inter8));
  nand2 gate1242(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1243(.a(s_99), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1244(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1245(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1246(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1905(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1906(.a(gate237inter0), .b(s_194), .O(gate237inter1));
  and2  gate1907(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1908(.a(s_194), .O(gate237inter3));
  inv1  gate1909(.a(s_195), .O(gate237inter4));
  nand2 gate1910(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1911(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1912(.a(G254), .O(gate237inter7));
  inv1  gate1913(.a(G706), .O(gate237inter8));
  nand2 gate1914(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1915(.a(s_195), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1916(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1917(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1918(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1163(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1164(.a(gate238inter0), .b(s_88), .O(gate238inter1));
  and2  gate1165(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1166(.a(s_88), .O(gate238inter3));
  inv1  gate1167(.a(s_89), .O(gate238inter4));
  nand2 gate1168(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1169(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1170(.a(G257), .O(gate238inter7));
  inv1  gate1171(.a(G709), .O(gate238inter8));
  nand2 gate1172(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1173(.a(s_89), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1174(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1175(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1176(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1639(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1640(.a(gate242inter0), .b(s_156), .O(gate242inter1));
  and2  gate1641(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1642(.a(s_156), .O(gate242inter3));
  inv1  gate1643(.a(s_157), .O(gate242inter4));
  nand2 gate1644(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1645(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1646(.a(G718), .O(gate242inter7));
  inv1  gate1647(.a(G730), .O(gate242inter8));
  nand2 gate1648(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1649(.a(s_157), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1650(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1651(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1652(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate2227(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2228(.a(gate243inter0), .b(s_240), .O(gate243inter1));
  and2  gate2229(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2230(.a(s_240), .O(gate243inter3));
  inv1  gate2231(.a(s_241), .O(gate243inter4));
  nand2 gate2232(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2233(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2234(.a(G245), .O(gate243inter7));
  inv1  gate2235(.a(G733), .O(gate243inter8));
  nand2 gate2236(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2237(.a(s_241), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2238(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2239(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2240(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2815(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2816(.a(gate245inter0), .b(s_324), .O(gate245inter1));
  and2  gate2817(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2818(.a(s_324), .O(gate245inter3));
  inv1  gate2819(.a(s_325), .O(gate245inter4));
  nand2 gate2820(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2821(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2822(.a(G248), .O(gate245inter7));
  inv1  gate2823(.a(G736), .O(gate245inter8));
  nand2 gate2824(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2825(.a(s_325), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2826(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2827(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2828(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate561(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate562(.a(gate248inter0), .b(s_2), .O(gate248inter1));
  and2  gate563(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate564(.a(s_2), .O(gate248inter3));
  inv1  gate565(.a(s_3), .O(gate248inter4));
  nand2 gate566(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate567(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate568(.a(G727), .O(gate248inter7));
  inv1  gate569(.a(G739), .O(gate248inter8));
  nand2 gate570(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate571(.a(s_3), .b(gate248inter3), .O(gate248inter10));
  nor2  gate572(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate573(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate574(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2423(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2424(.a(gate250inter0), .b(s_268), .O(gate250inter1));
  and2  gate2425(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2426(.a(s_268), .O(gate250inter3));
  inv1  gate2427(.a(s_269), .O(gate250inter4));
  nand2 gate2428(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2429(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2430(.a(G706), .O(gate250inter7));
  inv1  gate2431(.a(G742), .O(gate250inter8));
  nand2 gate2432(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2433(.a(s_269), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2434(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2435(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2436(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1219(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1220(.a(gate251inter0), .b(s_96), .O(gate251inter1));
  and2  gate1221(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1222(.a(s_96), .O(gate251inter3));
  inv1  gate1223(.a(s_97), .O(gate251inter4));
  nand2 gate1224(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1225(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1226(.a(G257), .O(gate251inter7));
  inv1  gate1227(.a(G745), .O(gate251inter8));
  nand2 gate1228(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1229(.a(s_97), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1230(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1231(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1232(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1513(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1514(.a(gate253inter0), .b(s_138), .O(gate253inter1));
  and2  gate1515(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1516(.a(s_138), .O(gate253inter3));
  inv1  gate1517(.a(s_139), .O(gate253inter4));
  nand2 gate1518(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1519(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1520(.a(G260), .O(gate253inter7));
  inv1  gate1521(.a(G748), .O(gate253inter8));
  nand2 gate1522(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1523(.a(s_139), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1524(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1525(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1526(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate2647(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2648(.a(gate254inter0), .b(s_300), .O(gate254inter1));
  and2  gate2649(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2650(.a(s_300), .O(gate254inter3));
  inv1  gate2651(.a(s_301), .O(gate254inter4));
  nand2 gate2652(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2653(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2654(.a(G712), .O(gate254inter7));
  inv1  gate2655(.a(G748), .O(gate254inter8));
  nand2 gate2656(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2657(.a(s_301), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2658(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2659(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2660(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1793(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1794(.a(gate255inter0), .b(s_178), .O(gate255inter1));
  and2  gate1795(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1796(.a(s_178), .O(gate255inter3));
  inv1  gate1797(.a(s_179), .O(gate255inter4));
  nand2 gate1798(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1799(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1800(.a(G263), .O(gate255inter7));
  inv1  gate1801(.a(G751), .O(gate255inter8));
  nand2 gate1802(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1803(.a(s_179), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1804(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1805(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1806(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1359(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1360(.a(gate256inter0), .b(s_116), .O(gate256inter1));
  and2  gate1361(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1362(.a(s_116), .O(gate256inter3));
  inv1  gate1363(.a(s_117), .O(gate256inter4));
  nand2 gate1364(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1365(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1366(.a(G715), .O(gate256inter7));
  inv1  gate1367(.a(G751), .O(gate256inter8));
  nand2 gate1368(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1369(.a(s_117), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1370(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1371(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1372(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate2437(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2438(.a(gate259inter0), .b(s_270), .O(gate259inter1));
  and2  gate2439(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2440(.a(s_270), .O(gate259inter3));
  inv1  gate2441(.a(s_271), .O(gate259inter4));
  nand2 gate2442(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2443(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2444(.a(G758), .O(gate259inter7));
  inv1  gate2445(.a(G759), .O(gate259inter8));
  nand2 gate2446(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2447(.a(s_271), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2448(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2449(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2450(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1317(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1318(.a(gate260inter0), .b(s_110), .O(gate260inter1));
  and2  gate1319(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1320(.a(s_110), .O(gate260inter3));
  inv1  gate1321(.a(s_111), .O(gate260inter4));
  nand2 gate1322(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1323(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1324(.a(G760), .O(gate260inter7));
  inv1  gate1325(.a(G761), .O(gate260inter8));
  nand2 gate1326(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1327(.a(s_111), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1328(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1329(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1330(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1205(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1206(.a(gate261inter0), .b(s_94), .O(gate261inter1));
  and2  gate1207(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1208(.a(s_94), .O(gate261inter3));
  inv1  gate1209(.a(s_95), .O(gate261inter4));
  nand2 gate1210(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1211(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1212(.a(G762), .O(gate261inter7));
  inv1  gate1213(.a(G763), .O(gate261inter8));
  nand2 gate1214(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1215(.a(s_95), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1216(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1217(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1218(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2773(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2774(.a(gate264inter0), .b(s_318), .O(gate264inter1));
  and2  gate2775(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2776(.a(s_318), .O(gate264inter3));
  inv1  gate2777(.a(s_319), .O(gate264inter4));
  nand2 gate2778(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2779(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2780(.a(G768), .O(gate264inter7));
  inv1  gate2781(.a(G769), .O(gate264inter8));
  nand2 gate2782(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2783(.a(s_319), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2784(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2785(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2786(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate673(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate674(.a(gate266inter0), .b(s_18), .O(gate266inter1));
  and2  gate675(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate676(.a(s_18), .O(gate266inter3));
  inv1  gate677(.a(s_19), .O(gate266inter4));
  nand2 gate678(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate679(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate680(.a(G645), .O(gate266inter7));
  inv1  gate681(.a(G773), .O(gate266inter8));
  nand2 gate682(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate683(.a(s_19), .b(gate266inter3), .O(gate266inter10));
  nor2  gate684(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate685(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate686(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2535(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2536(.a(gate267inter0), .b(s_284), .O(gate267inter1));
  and2  gate2537(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2538(.a(s_284), .O(gate267inter3));
  inv1  gate2539(.a(s_285), .O(gate267inter4));
  nand2 gate2540(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2541(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2542(.a(G648), .O(gate267inter7));
  inv1  gate2543(.a(G776), .O(gate267inter8));
  nand2 gate2544(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2545(.a(s_285), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2546(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2547(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2548(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2787(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2788(.a(gate268inter0), .b(s_320), .O(gate268inter1));
  and2  gate2789(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2790(.a(s_320), .O(gate268inter3));
  inv1  gate2791(.a(s_321), .O(gate268inter4));
  nand2 gate2792(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2793(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2794(.a(G651), .O(gate268inter7));
  inv1  gate2795(.a(G779), .O(gate268inter8));
  nand2 gate2796(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2797(.a(s_321), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2798(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2799(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2800(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1835(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1836(.a(gate270inter0), .b(s_184), .O(gate270inter1));
  and2  gate1837(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1838(.a(s_184), .O(gate270inter3));
  inv1  gate1839(.a(s_185), .O(gate270inter4));
  nand2 gate1840(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1841(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1842(.a(G657), .O(gate270inter7));
  inv1  gate1843(.a(G785), .O(gate270inter8));
  nand2 gate1844(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1845(.a(s_185), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1846(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1847(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1848(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate827(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate828(.a(gate271inter0), .b(s_40), .O(gate271inter1));
  and2  gate829(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate830(.a(s_40), .O(gate271inter3));
  inv1  gate831(.a(s_41), .O(gate271inter4));
  nand2 gate832(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate833(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate834(.a(G660), .O(gate271inter7));
  inv1  gate835(.a(G788), .O(gate271inter8));
  nand2 gate836(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate837(.a(s_41), .b(gate271inter3), .O(gate271inter10));
  nor2  gate838(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate839(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate840(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1779(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1780(.a(gate273inter0), .b(s_176), .O(gate273inter1));
  and2  gate1781(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1782(.a(s_176), .O(gate273inter3));
  inv1  gate1783(.a(s_177), .O(gate273inter4));
  nand2 gate1784(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1785(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1786(.a(G642), .O(gate273inter7));
  inv1  gate1787(.a(G794), .O(gate273inter8));
  nand2 gate1788(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1789(.a(s_177), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1790(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1791(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1792(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1415(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1416(.a(gate274inter0), .b(s_124), .O(gate274inter1));
  and2  gate1417(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1418(.a(s_124), .O(gate274inter3));
  inv1  gate1419(.a(s_125), .O(gate274inter4));
  nand2 gate1420(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1421(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1422(.a(G770), .O(gate274inter7));
  inv1  gate1423(.a(G794), .O(gate274inter8));
  nand2 gate1424(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1425(.a(s_125), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1426(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1427(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1428(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2409(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2410(.a(gate275inter0), .b(s_266), .O(gate275inter1));
  and2  gate2411(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2412(.a(s_266), .O(gate275inter3));
  inv1  gate2413(.a(s_267), .O(gate275inter4));
  nand2 gate2414(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2415(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2416(.a(G645), .O(gate275inter7));
  inv1  gate2417(.a(G797), .O(gate275inter8));
  nand2 gate2418(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2419(.a(s_267), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2420(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2421(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2422(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate2843(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2844(.a(gate276inter0), .b(s_328), .O(gate276inter1));
  and2  gate2845(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2846(.a(s_328), .O(gate276inter3));
  inv1  gate2847(.a(s_329), .O(gate276inter4));
  nand2 gate2848(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2849(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2850(.a(G773), .O(gate276inter7));
  inv1  gate2851(.a(G797), .O(gate276inter8));
  nand2 gate2852(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2853(.a(s_329), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2854(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2855(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2856(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1471(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1472(.a(gate278inter0), .b(s_132), .O(gate278inter1));
  and2  gate1473(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1474(.a(s_132), .O(gate278inter3));
  inv1  gate1475(.a(s_133), .O(gate278inter4));
  nand2 gate1476(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1477(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1478(.a(G776), .O(gate278inter7));
  inv1  gate1479(.a(G800), .O(gate278inter8));
  nand2 gate1480(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1481(.a(s_133), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1482(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1483(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1484(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2143(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2144(.a(gate280inter0), .b(s_228), .O(gate280inter1));
  and2  gate2145(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2146(.a(s_228), .O(gate280inter3));
  inv1  gate2147(.a(s_229), .O(gate280inter4));
  nand2 gate2148(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2149(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2150(.a(G779), .O(gate280inter7));
  inv1  gate2151(.a(G803), .O(gate280inter8));
  nand2 gate2152(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2153(.a(s_229), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2154(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2155(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2156(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2311(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2312(.a(gate285inter0), .b(s_252), .O(gate285inter1));
  and2  gate2313(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2314(.a(s_252), .O(gate285inter3));
  inv1  gate2315(.a(s_253), .O(gate285inter4));
  nand2 gate2316(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2317(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2318(.a(G660), .O(gate285inter7));
  inv1  gate2319(.a(G812), .O(gate285inter8));
  nand2 gate2320(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2321(.a(s_253), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2322(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2323(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2324(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2115(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2116(.a(gate286inter0), .b(s_224), .O(gate286inter1));
  and2  gate2117(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2118(.a(s_224), .O(gate286inter3));
  inv1  gate2119(.a(s_225), .O(gate286inter4));
  nand2 gate2120(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2121(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2122(.a(G788), .O(gate286inter7));
  inv1  gate2123(.a(G812), .O(gate286inter8));
  nand2 gate2124(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2125(.a(s_225), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2126(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2127(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2128(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2577(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2578(.a(gate288inter0), .b(s_290), .O(gate288inter1));
  and2  gate2579(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2580(.a(s_290), .O(gate288inter3));
  inv1  gate2581(.a(s_291), .O(gate288inter4));
  nand2 gate2582(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2583(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2584(.a(G791), .O(gate288inter7));
  inv1  gate2585(.a(G815), .O(gate288inter8));
  nand2 gate2586(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2587(.a(s_291), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2588(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2589(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2590(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2157(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2158(.a(gate292inter0), .b(s_230), .O(gate292inter1));
  and2  gate2159(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2160(.a(s_230), .O(gate292inter3));
  inv1  gate2161(.a(s_231), .O(gate292inter4));
  nand2 gate2162(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2163(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2164(.a(G824), .O(gate292inter7));
  inv1  gate2165(.a(G825), .O(gate292inter8));
  nand2 gate2166(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2167(.a(s_231), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2168(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2169(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2170(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1303(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1304(.a(gate293inter0), .b(s_108), .O(gate293inter1));
  and2  gate1305(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1306(.a(s_108), .O(gate293inter3));
  inv1  gate1307(.a(s_109), .O(gate293inter4));
  nand2 gate1308(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1309(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1310(.a(G828), .O(gate293inter7));
  inv1  gate1311(.a(G829), .O(gate293inter8));
  nand2 gate1312(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1313(.a(s_109), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1314(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1315(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1316(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1275(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1276(.a(gate390inter0), .b(s_104), .O(gate390inter1));
  and2  gate1277(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1278(.a(s_104), .O(gate390inter3));
  inv1  gate1279(.a(s_105), .O(gate390inter4));
  nand2 gate1280(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1281(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1282(.a(G4), .O(gate390inter7));
  inv1  gate1283(.a(G1045), .O(gate390inter8));
  nand2 gate1284(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1285(.a(s_105), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1286(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1287(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1288(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2521(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2522(.a(gate393inter0), .b(s_282), .O(gate393inter1));
  and2  gate2523(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2524(.a(s_282), .O(gate393inter3));
  inv1  gate2525(.a(s_283), .O(gate393inter4));
  nand2 gate2526(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2527(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2528(.a(G7), .O(gate393inter7));
  inv1  gate2529(.a(G1054), .O(gate393inter8));
  nand2 gate2530(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2531(.a(s_283), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2532(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2533(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2534(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1177(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1178(.a(gate396inter0), .b(s_90), .O(gate396inter1));
  and2  gate1179(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1180(.a(s_90), .O(gate396inter3));
  inv1  gate1181(.a(s_91), .O(gate396inter4));
  nand2 gate1182(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1183(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1184(.a(G10), .O(gate396inter7));
  inv1  gate1185(.a(G1063), .O(gate396inter8));
  nand2 gate1186(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1187(.a(s_91), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1188(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1189(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1190(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2171(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2172(.a(gate401inter0), .b(s_232), .O(gate401inter1));
  and2  gate2173(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2174(.a(s_232), .O(gate401inter3));
  inv1  gate2175(.a(s_233), .O(gate401inter4));
  nand2 gate2176(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2177(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2178(.a(G15), .O(gate401inter7));
  inv1  gate2179(.a(G1078), .O(gate401inter8));
  nand2 gate2180(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2181(.a(s_233), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2182(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2183(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2184(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2451(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2452(.a(gate403inter0), .b(s_272), .O(gate403inter1));
  and2  gate2453(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2454(.a(s_272), .O(gate403inter3));
  inv1  gate2455(.a(s_273), .O(gate403inter4));
  nand2 gate2456(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2457(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2458(.a(G17), .O(gate403inter7));
  inv1  gate2459(.a(G1084), .O(gate403inter8));
  nand2 gate2460(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2461(.a(s_273), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2462(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2463(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2464(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1653(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1654(.a(gate404inter0), .b(s_158), .O(gate404inter1));
  and2  gate1655(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1656(.a(s_158), .O(gate404inter3));
  inv1  gate1657(.a(s_159), .O(gate404inter4));
  nand2 gate1658(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1659(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1660(.a(G18), .O(gate404inter7));
  inv1  gate1661(.a(G1087), .O(gate404inter8));
  nand2 gate1662(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1663(.a(s_159), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1664(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1665(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1666(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2619(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2620(.a(gate406inter0), .b(s_296), .O(gate406inter1));
  and2  gate2621(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2622(.a(s_296), .O(gate406inter3));
  inv1  gate2623(.a(s_297), .O(gate406inter4));
  nand2 gate2624(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2625(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2626(.a(G20), .O(gate406inter7));
  inv1  gate2627(.a(G1093), .O(gate406inter8));
  nand2 gate2628(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2629(.a(s_297), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2630(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2631(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2632(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1527(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1528(.a(gate411inter0), .b(s_140), .O(gate411inter1));
  and2  gate1529(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1530(.a(s_140), .O(gate411inter3));
  inv1  gate1531(.a(s_141), .O(gate411inter4));
  nand2 gate1532(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1533(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1534(.a(G25), .O(gate411inter7));
  inv1  gate1535(.a(G1108), .O(gate411inter8));
  nand2 gate1536(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1537(.a(s_141), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1538(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1539(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1540(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1135(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1136(.a(gate420inter0), .b(s_84), .O(gate420inter1));
  and2  gate1137(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1138(.a(s_84), .O(gate420inter3));
  inv1  gate1139(.a(s_85), .O(gate420inter4));
  nand2 gate1140(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1141(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1142(.a(G1036), .O(gate420inter7));
  inv1  gate1143(.a(G1132), .O(gate420inter8));
  nand2 gate1144(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1145(.a(s_85), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1146(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1147(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1148(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate701(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate702(.a(gate421inter0), .b(s_22), .O(gate421inter1));
  and2  gate703(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate704(.a(s_22), .O(gate421inter3));
  inv1  gate705(.a(s_23), .O(gate421inter4));
  nand2 gate706(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate707(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate708(.a(G2), .O(gate421inter7));
  inv1  gate709(.a(G1135), .O(gate421inter8));
  nand2 gate710(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate711(.a(s_23), .b(gate421inter3), .O(gate421inter10));
  nor2  gate712(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate713(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate714(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1583(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1584(.a(gate424inter0), .b(s_148), .O(gate424inter1));
  and2  gate1585(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1586(.a(s_148), .O(gate424inter3));
  inv1  gate1587(.a(s_149), .O(gate424inter4));
  nand2 gate1588(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1589(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1590(.a(G1042), .O(gate424inter7));
  inv1  gate1591(.a(G1138), .O(gate424inter8));
  nand2 gate1592(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1593(.a(s_149), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1594(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1595(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1596(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate925(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate926(.a(gate426inter0), .b(s_54), .O(gate426inter1));
  and2  gate927(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate928(.a(s_54), .O(gate426inter3));
  inv1  gate929(.a(s_55), .O(gate426inter4));
  nand2 gate930(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate931(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate932(.a(G1045), .O(gate426inter7));
  inv1  gate933(.a(G1141), .O(gate426inter8));
  nand2 gate934(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate935(.a(s_55), .b(gate426inter3), .O(gate426inter10));
  nor2  gate936(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate937(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate938(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1919(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1920(.a(gate428inter0), .b(s_196), .O(gate428inter1));
  and2  gate1921(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1922(.a(s_196), .O(gate428inter3));
  inv1  gate1923(.a(s_197), .O(gate428inter4));
  nand2 gate1924(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1925(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1926(.a(G1048), .O(gate428inter7));
  inv1  gate1927(.a(G1144), .O(gate428inter8));
  nand2 gate1928(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1929(.a(s_197), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1930(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1931(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1932(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2031(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2032(.a(gate430inter0), .b(s_212), .O(gate430inter1));
  and2  gate2033(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2034(.a(s_212), .O(gate430inter3));
  inv1  gate2035(.a(s_213), .O(gate430inter4));
  nand2 gate2036(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2037(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2038(.a(G1051), .O(gate430inter7));
  inv1  gate2039(.a(G1147), .O(gate430inter8));
  nand2 gate2040(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2041(.a(s_213), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2042(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2043(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2044(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate547(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate548(.a(gate432inter0), .b(s_0), .O(gate432inter1));
  and2  gate549(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate550(.a(s_0), .O(gate432inter3));
  inv1  gate551(.a(s_1), .O(gate432inter4));
  nand2 gate552(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate553(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate554(.a(G1054), .O(gate432inter7));
  inv1  gate555(.a(G1150), .O(gate432inter8));
  nand2 gate556(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate557(.a(s_1), .b(gate432inter3), .O(gate432inter10));
  nor2  gate558(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate559(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate560(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1765(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1766(.a(gate433inter0), .b(s_174), .O(gate433inter1));
  and2  gate1767(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1768(.a(s_174), .O(gate433inter3));
  inv1  gate1769(.a(s_175), .O(gate433inter4));
  nand2 gate1770(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1771(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1772(.a(G8), .O(gate433inter7));
  inv1  gate1773(.a(G1153), .O(gate433inter8));
  nand2 gate1774(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1775(.a(s_175), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1776(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1777(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1778(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate2801(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2802(.a(gate434inter0), .b(s_322), .O(gate434inter1));
  and2  gate2803(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2804(.a(s_322), .O(gate434inter3));
  inv1  gate2805(.a(s_323), .O(gate434inter4));
  nand2 gate2806(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2807(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2808(.a(G1057), .O(gate434inter7));
  inv1  gate2809(.a(G1153), .O(gate434inter8));
  nand2 gate2810(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2811(.a(s_323), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2812(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2813(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2814(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2661(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2662(.a(gate435inter0), .b(s_302), .O(gate435inter1));
  and2  gate2663(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2664(.a(s_302), .O(gate435inter3));
  inv1  gate2665(.a(s_303), .O(gate435inter4));
  nand2 gate2666(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2667(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2668(.a(G9), .O(gate435inter7));
  inv1  gate2669(.a(G1156), .O(gate435inter8));
  nand2 gate2670(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2671(.a(s_303), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2672(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2673(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2674(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2465(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2466(.a(gate440inter0), .b(s_274), .O(gate440inter1));
  and2  gate2467(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2468(.a(s_274), .O(gate440inter3));
  inv1  gate2469(.a(s_275), .O(gate440inter4));
  nand2 gate2470(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2471(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2472(.a(G1066), .O(gate440inter7));
  inv1  gate2473(.a(G1162), .O(gate440inter8));
  nand2 gate2474(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2475(.a(s_275), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2476(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2477(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2478(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1191(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1192(.a(gate443inter0), .b(s_92), .O(gate443inter1));
  and2  gate1193(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1194(.a(s_92), .O(gate443inter3));
  inv1  gate1195(.a(s_93), .O(gate443inter4));
  nand2 gate1196(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1197(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1198(.a(G13), .O(gate443inter7));
  inv1  gate1199(.a(G1168), .O(gate443inter8));
  nand2 gate1200(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1201(.a(s_93), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1202(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1203(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1204(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2325(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2326(.a(gate445inter0), .b(s_254), .O(gate445inter1));
  and2  gate2327(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2328(.a(s_254), .O(gate445inter3));
  inv1  gate2329(.a(s_255), .O(gate445inter4));
  nand2 gate2330(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2331(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2332(.a(G14), .O(gate445inter7));
  inv1  gate2333(.a(G1171), .O(gate445inter8));
  nand2 gate2334(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2335(.a(s_255), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2336(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2337(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2338(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1709(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1710(.a(gate447inter0), .b(s_166), .O(gate447inter1));
  and2  gate1711(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1712(.a(s_166), .O(gate447inter3));
  inv1  gate1713(.a(s_167), .O(gate447inter4));
  nand2 gate1714(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1715(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1716(.a(G15), .O(gate447inter7));
  inv1  gate1717(.a(G1174), .O(gate447inter8));
  nand2 gate1718(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1719(.a(s_167), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1720(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1721(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1722(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2479(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2480(.a(gate452inter0), .b(s_276), .O(gate452inter1));
  and2  gate2481(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2482(.a(s_276), .O(gate452inter3));
  inv1  gate2483(.a(s_277), .O(gate452inter4));
  nand2 gate2484(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2485(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2486(.a(G1084), .O(gate452inter7));
  inv1  gate2487(.a(G1180), .O(gate452inter8));
  nand2 gate2488(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2489(.a(s_277), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2490(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2491(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2492(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1751(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1752(.a(gate454inter0), .b(s_172), .O(gate454inter1));
  and2  gate1753(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1754(.a(s_172), .O(gate454inter3));
  inv1  gate1755(.a(s_173), .O(gate454inter4));
  nand2 gate1756(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1757(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1758(.a(G1087), .O(gate454inter7));
  inv1  gate1759(.a(G1183), .O(gate454inter8));
  nand2 gate1760(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1761(.a(s_173), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1762(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1763(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1764(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate2017(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2018(.a(gate455inter0), .b(s_210), .O(gate455inter1));
  and2  gate2019(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2020(.a(s_210), .O(gate455inter3));
  inv1  gate2021(.a(s_211), .O(gate455inter4));
  nand2 gate2022(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2023(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2024(.a(G19), .O(gate455inter7));
  inv1  gate2025(.a(G1186), .O(gate455inter8));
  nand2 gate2026(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2027(.a(s_211), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2028(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2029(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2030(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2703(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2704(.a(gate459inter0), .b(s_308), .O(gate459inter1));
  and2  gate2705(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2706(.a(s_308), .O(gate459inter3));
  inv1  gate2707(.a(s_309), .O(gate459inter4));
  nand2 gate2708(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2709(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2710(.a(G21), .O(gate459inter7));
  inv1  gate2711(.a(G1192), .O(gate459inter8));
  nand2 gate2712(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2713(.a(s_309), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2714(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2715(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2716(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1569(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1570(.a(gate461inter0), .b(s_146), .O(gate461inter1));
  and2  gate1571(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1572(.a(s_146), .O(gate461inter3));
  inv1  gate1573(.a(s_147), .O(gate461inter4));
  nand2 gate1574(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1575(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1576(.a(G22), .O(gate461inter7));
  inv1  gate1577(.a(G1195), .O(gate461inter8));
  nand2 gate1578(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1579(.a(s_147), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1580(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1581(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1582(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2493(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2494(.a(gate464inter0), .b(s_278), .O(gate464inter1));
  and2  gate2495(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2496(.a(s_278), .O(gate464inter3));
  inv1  gate2497(.a(s_279), .O(gate464inter4));
  nand2 gate2498(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2499(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2500(.a(G1102), .O(gate464inter7));
  inv1  gate2501(.a(G1198), .O(gate464inter8));
  nand2 gate2502(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2503(.a(s_279), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2504(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2505(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2506(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2395(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2396(.a(gate467inter0), .b(s_264), .O(gate467inter1));
  and2  gate2397(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2398(.a(s_264), .O(gate467inter3));
  inv1  gate2399(.a(s_265), .O(gate467inter4));
  nand2 gate2400(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2401(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2402(.a(G25), .O(gate467inter7));
  inv1  gate2403(.a(G1204), .O(gate467inter8));
  nand2 gate2404(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2405(.a(s_265), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2406(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2407(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2408(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2633(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2634(.a(gate472inter0), .b(s_298), .O(gate472inter1));
  and2  gate2635(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2636(.a(s_298), .O(gate472inter3));
  inv1  gate2637(.a(s_299), .O(gate472inter4));
  nand2 gate2638(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2639(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2640(.a(G1114), .O(gate472inter7));
  inv1  gate2641(.a(G1210), .O(gate472inter8));
  nand2 gate2642(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2643(.a(s_299), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2644(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2645(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2646(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate2563(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2564(.a(gate473inter0), .b(s_288), .O(gate473inter1));
  and2  gate2565(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2566(.a(s_288), .O(gate473inter3));
  inv1  gate2567(.a(s_289), .O(gate473inter4));
  nand2 gate2568(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2569(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2570(.a(G28), .O(gate473inter7));
  inv1  gate2571(.a(G1213), .O(gate473inter8));
  nand2 gate2572(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2573(.a(s_289), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2574(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2575(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2576(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate981(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate982(.a(gate477inter0), .b(s_62), .O(gate477inter1));
  and2  gate983(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate984(.a(s_62), .O(gate477inter3));
  inv1  gate985(.a(s_63), .O(gate477inter4));
  nand2 gate986(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate987(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate988(.a(G30), .O(gate477inter7));
  inv1  gate989(.a(G1219), .O(gate477inter8));
  nand2 gate990(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate991(.a(s_63), .b(gate477inter3), .O(gate477inter10));
  nor2  gate992(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate993(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate994(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate2297(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2298(.a(gate481inter0), .b(s_250), .O(gate481inter1));
  and2  gate2299(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2300(.a(s_250), .O(gate481inter3));
  inv1  gate2301(.a(s_251), .O(gate481inter4));
  nand2 gate2302(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2303(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2304(.a(G32), .O(gate481inter7));
  inv1  gate2305(.a(G1225), .O(gate481inter8));
  nand2 gate2306(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2307(.a(s_251), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2308(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2309(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2310(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate715(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate716(.a(gate482inter0), .b(s_24), .O(gate482inter1));
  and2  gate717(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate718(.a(s_24), .O(gate482inter3));
  inv1  gate719(.a(s_25), .O(gate482inter4));
  nand2 gate720(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate721(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate722(.a(G1129), .O(gate482inter7));
  inv1  gate723(.a(G1225), .O(gate482inter8));
  nand2 gate724(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate725(.a(s_25), .b(gate482inter3), .O(gate482inter10));
  nor2  gate726(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate727(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate728(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2367(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2368(.a(gate485inter0), .b(s_260), .O(gate485inter1));
  and2  gate2369(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2370(.a(s_260), .O(gate485inter3));
  inv1  gate2371(.a(s_261), .O(gate485inter4));
  nand2 gate2372(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2373(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2374(.a(G1232), .O(gate485inter7));
  inv1  gate2375(.a(G1233), .O(gate485inter8));
  nand2 gate2376(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2377(.a(s_261), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2378(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2379(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2380(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1373(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1374(.a(gate487inter0), .b(s_118), .O(gate487inter1));
  and2  gate1375(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1376(.a(s_118), .O(gate487inter3));
  inv1  gate1377(.a(s_119), .O(gate487inter4));
  nand2 gate1378(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1379(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1380(.a(G1236), .O(gate487inter7));
  inv1  gate1381(.a(G1237), .O(gate487inter8));
  nand2 gate1382(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1383(.a(s_119), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1384(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1385(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1386(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2283(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2284(.a(gate490inter0), .b(s_248), .O(gate490inter1));
  and2  gate2285(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2286(.a(s_248), .O(gate490inter3));
  inv1  gate2287(.a(s_249), .O(gate490inter4));
  nand2 gate2288(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2289(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2290(.a(G1242), .O(gate490inter7));
  inv1  gate2291(.a(G1243), .O(gate490inter8));
  nand2 gate2292(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2293(.a(s_249), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2294(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2295(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2296(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1961(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1962(.a(gate500inter0), .b(s_202), .O(gate500inter1));
  and2  gate1963(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1964(.a(s_202), .O(gate500inter3));
  inv1  gate1965(.a(s_203), .O(gate500inter4));
  nand2 gate1966(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1967(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1968(.a(G1262), .O(gate500inter7));
  inv1  gate1969(.a(G1263), .O(gate500inter8));
  nand2 gate1970(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1971(.a(s_203), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1972(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1973(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1974(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1429(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1430(.a(gate501inter0), .b(s_126), .O(gate501inter1));
  and2  gate1431(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1432(.a(s_126), .O(gate501inter3));
  inv1  gate1433(.a(s_127), .O(gate501inter4));
  nand2 gate1434(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1435(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1436(.a(G1264), .O(gate501inter7));
  inv1  gate1437(.a(G1265), .O(gate501inter8));
  nand2 gate1438(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1439(.a(s_127), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1440(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1441(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1442(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2731(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2732(.a(gate503inter0), .b(s_312), .O(gate503inter1));
  and2  gate2733(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2734(.a(s_312), .O(gate503inter3));
  inv1  gate2735(.a(s_313), .O(gate503inter4));
  nand2 gate2736(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2737(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2738(.a(G1268), .O(gate503inter7));
  inv1  gate2739(.a(G1269), .O(gate503inter8));
  nand2 gate2740(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2741(.a(s_313), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2742(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2743(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2744(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate757(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate758(.a(gate508inter0), .b(s_30), .O(gate508inter1));
  and2  gate759(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate760(.a(s_30), .O(gate508inter3));
  inv1  gate761(.a(s_31), .O(gate508inter4));
  nand2 gate762(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate763(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate764(.a(G1278), .O(gate508inter7));
  inv1  gate765(.a(G1279), .O(gate508inter8));
  nand2 gate766(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate767(.a(s_31), .b(gate508inter3), .O(gate508inter10));
  nor2  gate768(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate769(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate770(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate645(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate646(.a(gate512inter0), .b(s_14), .O(gate512inter1));
  and2  gate647(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate648(.a(s_14), .O(gate512inter3));
  inv1  gate649(.a(s_15), .O(gate512inter4));
  nand2 gate650(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate651(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate652(.a(G1286), .O(gate512inter7));
  inv1  gate653(.a(G1287), .O(gate512inter8));
  nand2 gate654(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate655(.a(s_15), .b(gate512inter3), .O(gate512inter10));
  nor2  gate656(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate657(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate658(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1821(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1822(.a(gate513inter0), .b(s_182), .O(gate513inter1));
  and2  gate1823(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1824(.a(s_182), .O(gate513inter3));
  inv1  gate1825(.a(s_183), .O(gate513inter4));
  nand2 gate1826(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1827(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1828(.a(G1288), .O(gate513inter7));
  inv1  gate1829(.a(G1289), .O(gate513inter8));
  nand2 gate1830(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1831(.a(s_183), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1832(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1833(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1834(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1261(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1262(.a(gate514inter0), .b(s_102), .O(gate514inter1));
  and2  gate1263(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1264(.a(s_102), .O(gate514inter3));
  inv1  gate1265(.a(s_103), .O(gate514inter4));
  nand2 gate1266(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1267(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1268(.a(G1290), .O(gate514inter7));
  inv1  gate1269(.a(G1291), .O(gate514inter8));
  nand2 gate1270(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1271(.a(s_103), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1272(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1273(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1274(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule