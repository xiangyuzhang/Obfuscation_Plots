module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2801(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2802(.a(gate9inter0), .b(s_322), .O(gate9inter1));
  and2  gate2803(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2804(.a(s_322), .O(gate9inter3));
  inv1  gate2805(.a(s_323), .O(gate9inter4));
  nand2 gate2806(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2807(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2808(.a(G1), .O(gate9inter7));
  inv1  gate2809(.a(G2), .O(gate9inter8));
  nand2 gate2810(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2811(.a(s_323), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2812(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2813(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2814(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2829(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2830(.a(gate14inter0), .b(s_326), .O(gate14inter1));
  and2  gate2831(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2832(.a(s_326), .O(gate14inter3));
  inv1  gate2833(.a(s_327), .O(gate14inter4));
  nand2 gate2834(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2835(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2836(.a(G11), .O(gate14inter7));
  inv1  gate2837(.a(G12), .O(gate14inter8));
  nand2 gate2838(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2839(.a(s_327), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2840(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2841(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2842(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1219(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1220(.a(gate15inter0), .b(s_96), .O(gate15inter1));
  and2  gate1221(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1222(.a(s_96), .O(gate15inter3));
  inv1  gate1223(.a(s_97), .O(gate15inter4));
  nand2 gate1224(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1225(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1226(.a(G13), .O(gate15inter7));
  inv1  gate1227(.a(G14), .O(gate15inter8));
  nand2 gate1228(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1229(.a(s_97), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1230(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1231(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1232(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2507(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2508(.a(gate16inter0), .b(s_280), .O(gate16inter1));
  and2  gate2509(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2510(.a(s_280), .O(gate16inter3));
  inv1  gate2511(.a(s_281), .O(gate16inter4));
  nand2 gate2512(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2513(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2514(.a(G15), .O(gate16inter7));
  inv1  gate2515(.a(G16), .O(gate16inter8));
  nand2 gate2516(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2517(.a(s_281), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2518(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2519(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2520(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate701(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate702(.a(gate18inter0), .b(s_22), .O(gate18inter1));
  and2  gate703(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate704(.a(s_22), .O(gate18inter3));
  inv1  gate705(.a(s_23), .O(gate18inter4));
  nand2 gate706(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate707(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate708(.a(G19), .O(gate18inter7));
  inv1  gate709(.a(G20), .O(gate18inter8));
  nand2 gate710(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate711(.a(s_23), .b(gate18inter3), .O(gate18inter10));
  nor2  gate712(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate713(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate714(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate897(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate898(.a(gate19inter0), .b(s_50), .O(gate19inter1));
  and2  gate899(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate900(.a(s_50), .O(gate19inter3));
  inv1  gate901(.a(s_51), .O(gate19inter4));
  nand2 gate902(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate903(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate904(.a(G21), .O(gate19inter7));
  inv1  gate905(.a(G22), .O(gate19inter8));
  nand2 gate906(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate907(.a(s_51), .b(gate19inter3), .O(gate19inter10));
  nor2  gate908(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate909(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate910(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1247(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1248(.a(gate20inter0), .b(s_100), .O(gate20inter1));
  and2  gate1249(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1250(.a(s_100), .O(gate20inter3));
  inv1  gate1251(.a(s_101), .O(gate20inter4));
  nand2 gate1252(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1253(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1254(.a(G23), .O(gate20inter7));
  inv1  gate1255(.a(G24), .O(gate20inter8));
  nand2 gate1256(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1257(.a(s_101), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1258(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1259(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1260(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1457(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1458(.a(gate21inter0), .b(s_130), .O(gate21inter1));
  and2  gate1459(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1460(.a(s_130), .O(gate21inter3));
  inv1  gate1461(.a(s_131), .O(gate21inter4));
  nand2 gate1462(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1463(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1464(.a(G25), .O(gate21inter7));
  inv1  gate1465(.a(G26), .O(gate21inter8));
  nand2 gate1466(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1467(.a(s_131), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1468(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1469(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1470(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate631(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate632(.a(gate27inter0), .b(s_12), .O(gate27inter1));
  and2  gate633(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate634(.a(s_12), .O(gate27inter3));
  inv1  gate635(.a(s_13), .O(gate27inter4));
  nand2 gate636(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate637(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate638(.a(G2), .O(gate27inter7));
  inv1  gate639(.a(G6), .O(gate27inter8));
  nand2 gate640(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate641(.a(s_13), .b(gate27inter3), .O(gate27inter10));
  nor2  gate642(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate643(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate644(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1919(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1920(.a(gate34inter0), .b(s_196), .O(gate34inter1));
  and2  gate1921(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1922(.a(s_196), .O(gate34inter3));
  inv1  gate1923(.a(s_197), .O(gate34inter4));
  nand2 gate1924(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1925(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1926(.a(G25), .O(gate34inter7));
  inv1  gate1927(.a(G29), .O(gate34inter8));
  nand2 gate1928(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1929(.a(s_197), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1930(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1931(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1932(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2605(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2606(.a(gate37inter0), .b(s_294), .O(gate37inter1));
  and2  gate2607(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2608(.a(s_294), .O(gate37inter3));
  inv1  gate2609(.a(s_295), .O(gate37inter4));
  nand2 gate2610(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2611(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2612(.a(G19), .O(gate37inter7));
  inv1  gate2613(.a(G23), .O(gate37inter8));
  nand2 gate2614(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2615(.a(s_295), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2616(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2617(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2618(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1499(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1500(.a(gate41inter0), .b(s_136), .O(gate41inter1));
  and2  gate1501(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1502(.a(s_136), .O(gate41inter3));
  inv1  gate1503(.a(s_137), .O(gate41inter4));
  nand2 gate1504(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1505(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1506(.a(G1), .O(gate41inter7));
  inv1  gate1507(.a(G266), .O(gate41inter8));
  nand2 gate1508(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1509(.a(s_137), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1510(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1511(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1512(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2913(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2914(.a(gate44inter0), .b(s_338), .O(gate44inter1));
  and2  gate2915(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2916(.a(s_338), .O(gate44inter3));
  inv1  gate2917(.a(s_339), .O(gate44inter4));
  nand2 gate2918(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2919(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2920(.a(G4), .O(gate44inter7));
  inv1  gate2921(.a(G269), .O(gate44inter8));
  nand2 gate2922(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2923(.a(s_339), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2924(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2925(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2926(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2045(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2046(.a(gate48inter0), .b(s_214), .O(gate48inter1));
  and2  gate2047(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2048(.a(s_214), .O(gate48inter3));
  inv1  gate2049(.a(s_215), .O(gate48inter4));
  nand2 gate2050(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2051(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2052(.a(G8), .O(gate48inter7));
  inv1  gate2053(.a(G275), .O(gate48inter8));
  nand2 gate2054(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2055(.a(s_215), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2056(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2057(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2058(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1037(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1038(.a(gate49inter0), .b(s_70), .O(gate49inter1));
  and2  gate1039(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1040(.a(s_70), .O(gate49inter3));
  inv1  gate1041(.a(s_71), .O(gate49inter4));
  nand2 gate1042(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1043(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1044(.a(G9), .O(gate49inter7));
  inv1  gate1045(.a(G278), .O(gate49inter8));
  nand2 gate1046(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1047(.a(s_71), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1048(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1049(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1050(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate645(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate646(.a(gate50inter0), .b(s_14), .O(gate50inter1));
  and2  gate647(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate648(.a(s_14), .O(gate50inter3));
  inv1  gate649(.a(s_15), .O(gate50inter4));
  nand2 gate650(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate651(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate652(.a(G10), .O(gate50inter7));
  inv1  gate653(.a(G278), .O(gate50inter8));
  nand2 gate654(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate655(.a(s_15), .b(gate50inter3), .O(gate50inter10));
  nor2  gate656(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate657(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate658(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1821(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1822(.a(gate51inter0), .b(s_182), .O(gate51inter1));
  and2  gate1823(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1824(.a(s_182), .O(gate51inter3));
  inv1  gate1825(.a(s_183), .O(gate51inter4));
  nand2 gate1826(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1827(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1828(.a(G11), .O(gate51inter7));
  inv1  gate1829(.a(G281), .O(gate51inter8));
  nand2 gate1830(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1831(.a(s_183), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1832(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1833(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1834(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1135(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1136(.a(gate52inter0), .b(s_84), .O(gate52inter1));
  and2  gate1137(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1138(.a(s_84), .O(gate52inter3));
  inv1  gate1139(.a(s_85), .O(gate52inter4));
  nand2 gate1140(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1141(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1142(.a(G12), .O(gate52inter7));
  inv1  gate1143(.a(G281), .O(gate52inter8));
  nand2 gate1144(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1145(.a(s_85), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1146(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1147(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1148(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1597(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1598(.a(gate56inter0), .b(s_150), .O(gate56inter1));
  and2  gate1599(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1600(.a(s_150), .O(gate56inter3));
  inv1  gate1601(.a(s_151), .O(gate56inter4));
  nand2 gate1602(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1603(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1604(.a(G16), .O(gate56inter7));
  inv1  gate1605(.a(G287), .O(gate56inter8));
  nand2 gate1606(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1607(.a(s_151), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1608(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1609(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1610(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1737(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1738(.a(gate59inter0), .b(s_170), .O(gate59inter1));
  and2  gate1739(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1740(.a(s_170), .O(gate59inter3));
  inv1  gate1741(.a(s_171), .O(gate59inter4));
  nand2 gate1742(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1743(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1744(.a(G19), .O(gate59inter7));
  inv1  gate1745(.a(G293), .O(gate59inter8));
  nand2 gate1746(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1747(.a(s_171), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1748(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1749(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1750(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate925(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate926(.a(gate60inter0), .b(s_54), .O(gate60inter1));
  and2  gate927(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate928(.a(s_54), .O(gate60inter3));
  inv1  gate929(.a(s_55), .O(gate60inter4));
  nand2 gate930(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate931(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate932(.a(G20), .O(gate60inter7));
  inv1  gate933(.a(G293), .O(gate60inter8));
  nand2 gate934(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate935(.a(s_55), .b(gate60inter3), .O(gate60inter10));
  nor2  gate936(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate937(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate938(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2479(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2480(.a(gate62inter0), .b(s_276), .O(gate62inter1));
  and2  gate2481(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2482(.a(s_276), .O(gate62inter3));
  inv1  gate2483(.a(s_277), .O(gate62inter4));
  nand2 gate2484(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2485(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2486(.a(G22), .O(gate62inter7));
  inv1  gate2487(.a(G296), .O(gate62inter8));
  nand2 gate2488(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2489(.a(s_277), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2490(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2491(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2492(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2143(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2144(.a(gate63inter0), .b(s_228), .O(gate63inter1));
  and2  gate2145(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2146(.a(s_228), .O(gate63inter3));
  inv1  gate2147(.a(s_229), .O(gate63inter4));
  nand2 gate2148(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2149(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2150(.a(G23), .O(gate63inter7));
  inv1  gate2151(.a(G299), .O(gate63inter8));
  nand2 gate2152(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2153(.a(s_229), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2154(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2155(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2156(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1275(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1276(.a(gate66inter0), .b(s_104), .O(gate66inter1));
  and2  gate1277(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1278(.a(s_104), .O(gate66inter3));
  inv1  gate1279(.a(s_105), .O(gate66inter4));
  nand2 gate1280(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1281(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1282(.a(G26), .O(gate66inter7));
  inv1  gate1283(.a(G302), .O(gate66inter8));
  nand2 gate1284(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1285(.a(s_105), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1286(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1287(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1288(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1863(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1864(.a(gate67inter0), .b(s_188), .O(gate67inter1));
  and2  gate1865(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1866(.a(s_188), .O(gate67inter3));
  inv1  gate1867(.a(s_189), .O(gate67inter4));
  nand2 gate1868(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1869(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1870(.a(G27), .O(gate67inter7));
  inv1  gate1871(.a(G305), .O(gate67inter8));
  nand2 gate1872(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1873(.a(s_189), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1874(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1875(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1876(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1303(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1304(.a(gate71inter0), .b(s_108), .O(gate71inter1));
  and2  gate1305(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1306(.a(s_108), .O(gate71inter3));
  inv1  gate1307(.a(s_109), .O(gate71inter4));
  nand2 gate1308(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1309(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1310(.a(G31), .O(gate71inter7));
  inv1  gate1311(.a(G311), .O(gate71inter8));
  nand2 gate1312(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1313(.a(s_109), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1314(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1315(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1316(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate603(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate604(.a(gate78inter0), .b(s_8), .O(gate78inter1));
  and2  gate605(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate606(.a(s_8), .O(gate78inter3));
  inv1  gate607(.a(s_9), .O(gate78inter4));
  nand2 gate608(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate609(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate610(.a(G6), .O(gate78inter7));
  inv1  gate611(.a(G320), .O(gate78inter8));
  nand2 gate612(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate613(.a(s_9), .b(gate78inter3), .O(gate78inter10));
  nor2  gate614(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate615(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate616(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2395(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2396(.a(gate79inter0), .b(s_264), .O(gate79inter1));
  and2  gate2397(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2398(.a(s_264), .O(gate79inter3));
  inv1  gate2399(.a(s_265), .O(gate79inter4));
  nand2 gate2400(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2401(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2402(.a(G10), .O(gate79inter7));
  inv1  gate2403(.a(G323), .O(gate79inter8));
  nand2 gate2404(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2405(.a(s_265), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2406(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2407(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2408(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate673(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate674(.a(gate83inter0), .b(s_18), .O(gate83inter1));
  and2  gate675(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate676(.a(s_18), .O(gate83inter3));
  inv1  gate677(.a(s_19), .O(gate83inter4));
  nand2 gate678(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate679(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate680(.a(G11), .O(gate83inter7));
  inv1  gate681(.a(G329), .O(gate83inter8));
  nand2 gate682(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate683(.a(s_19), .b(gate83inter3), .O(gate83inter10));
  nor2  gate684(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate685(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate686(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate2871(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2872(.a(gate84inter0), .b(s_332), .O(gate84inter1));
  and2  gate2873(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2874(.a(s_332), .O(gate84inter3));
  inv1  gate2875(.a(s_333), .O(gate84inter4));
  nand2 gate2876(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2877(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2878(.a(G15), .O(gate84inter7));
  inv1  gate2879(.a(G329), .O(gate84inter8));
  nand2 gate2880(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2881(.a(s_333), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2882(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2883(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2884(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1751(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1752(.a(gate85inter0), .b(s_172), .O(gate85inter1));
  and2  gate1753(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1754(.a(s_172), .O(gate85inter3));
  inv1  gate1755(.a(s_173), .O(gate85inter4));
  nand2 gate1756(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1757(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1758(.a(G4), .O(gate85inter7));
  inv1  gate1759(.a(G332), .O(gate85inter8));
  nand2 gate1760(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1761(.a(s_173), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1762(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1763(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1764(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1793(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1794(.a(gate89inter0), .b(s_178), .O(gate89inter1));
  and2  gate1795(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1796(.a(s_178), .O(gate89inter3));
  inv1  gate1797(.a(s_179), .O(gate89inter4));
  nand2 gate1798(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1799(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1800(.a(G17), .O(gate89inter7));
  inv1  gate1801(.a(G338), .O(gate89inter8));
  nand2 gate1802(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1803(.a(s_179), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1804(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1805(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1806(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate2423(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2424(.a(gate90inter0), .b(s_268), .O(gate90inter1));
  and2  gate2425(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2426(.a(s_268), .O(gate90inter3));
  inv1  gate2427(.a(s_269), .O(gate90inter4));
  nand2 gate2428(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2429(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2430(.a(G21), .O(gate90inter7));
  inv1  gate2431(.a(G338), .O(gate90inter8));
  nand2 gate2432(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2433(.a(s_269), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2434(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2435(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2436(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate2353(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2354(.a(gate91inter0), .b(s_258), .O(gate91inter1));
  and2  gate2355(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2356(.a(s_258), .O(gate91inter3));
  inv1  gate2357(.a(s_259), .O(gate91inter4));
  nand2 gate2358(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2359(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2360(.a(G25), .O(gate91inter7));
  inv1  gate2361(.a(G341), .O(gate91inter8));
  nand2 gate2362(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2363(.a(s_259), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2364(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2365(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2366(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2633(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2634(.a(gate93inter0), .b(s_298), .O(gate93inter1));
  and2  gate2635(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2636(.a(s_298), .O(gate93inter3));
  inv1  gate2637(.a(s_299), .O(gate93inter4));
  nand2 gate2638(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2639(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2640(.a(G18), .O(gate93inter7));
  inv1  gate2641(.a(G344), .O(gate93inter8));
  nand2 gate2642(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2643(.a(s_299), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2644(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2645(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2646(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1387(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1388(.a(gate94inter0), .b(s_120), .O(gate94inter1));
  and2  gate1389(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1390(.a(s_120), .O(gate94inter3));
  inv1  gate1391(.a(s_121), .O(gate94inter4));
  nand2 gate1392(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1393(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1394(.a(G22), .O(gate94inter7));
  inv1  gate1395(.a(G344), .O(gate94inter8));
  nand2 gate1396(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1397(.a(s_121), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1398(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1399(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1400(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1009(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1010(.a(gate98inter0), .b(s_66), .O(gate98inter1));
  and2  gate1011(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1012(.a(s_66), .O(gate98inter3));
  inv1  gate1013(.a(s_67), .O(gate98inter4));
  nand2 gate1014(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1015(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1016(.a(G23), .O(gate98inter7));
  inv1  gate1017(.a(G350), .O(gate98inter8));
  nand2 gate1018(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1019(.a(s_67), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1020(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1021(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1022(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate2549(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate2550(.a(gate101inter0), .b(s_286), .O(gate101inter1));
  and2  gate2551(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate2552(.a(s_286), .O(gate101inter3));
  inv1  gate2553(.a(s_287), .O(gate101inter4));
  nand2 gate2554(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate2555(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate2556(.a(G20), .O(gate101inter7));
  inv1  gate2557(.a(G356), .O(gate101inter8));
  nand2 gate2558(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate2559(.a(s_287), .b(gate101inter3), .O(gate101inter10));
  nor2  gate2560(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate2561(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate2562(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1611(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1612(.a(gate104inter0), .b(s_152), .O(gate104inter1));
  and2  gate1613(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1614(.a(s_152), .O(gate104inter3));
  inv1  gate1615(.a(s_153), .O(gate104inter4));
  nand2 gate1616(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1617(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1618(.a(G32), .O(gate104inter7));
  inv1  gate1619(.a(G359), .O(gate104inter8));
  nand2 gate1620(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1621(.a(s_153), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1622(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1623(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1624(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2521(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2522(.a(gate106inter0), .b(s_282), .O(gate106inter1));
  and2  gate2523(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2524(.a(s_282), .O(gate106inter3));
  inv1  gate2525(.a(s_283), .O(gate106inter4));
  nand2 gate2526(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2527(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2528(.a(G364), .O(gate106inter7));
  inv1  gate2529(.a(G365), .O(gate106inter8));
  nand2 gate2530(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2531(.a(s_283), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2532(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2533(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2534(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2255(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2256(.a(gate107inter0), .b(s_244), .O(gate107inter1));
  and2  gate2257(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2258(.a(s_244), .O(gate107inter3));
  inv1  gate2259(.a(s_245), .O(gate107inter4));
  nand2 gate2260(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2261(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2262(.a(G366), .O(gate107inter7));
  inv1  gate2263(.a(G367), .O(gate107inter8));
  nand2 gate2264(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2265(.a(s_245), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2266(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2267(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2268(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1807(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1808(.a(gate109inter0), .b(s_180), .O(gate109inter1));
  and2  gate1809(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1810(.a(s_180), .O(gate109inter3));
  inv1  gate1811(.a(s_181), .O(gate109inter4));
  nand2 gate1812(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1813(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1814(.a(G370), .O(gate109inter7));
  inv1  gate1815(.a(G371), .O(gate109inter8));
  nand2 gate1816(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1817(.a(s_181), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1818(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1819(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1820(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate2199(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2200(.a(gate110inter0), .b(s_236), .O(gate110inter1));
  and2  gate2201(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2202(.a(s_236), .O(gate110inter3));
  inv1  gate2203(.a(s_237), .O(gate110inter4));
  nand2 gate2204(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2205(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2206(.a(G372), .O(gate110inter7));
  inv1  gate2207(.a(G373), .O(gate110inter8));
  nand2 gate2208(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2209(.a(s_237), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2210(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2211(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2212(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate883(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate884(.a(gate115inter0), .b(s_48), .O(gate115inter1));
  and2  gate885(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate886(.a(s_48), .O(gate115inter3));
  inv1  gate887(.a(s_49), .O(gate115inter4));
  nand2 gate888(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate889(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate890(.a(G382), .O(gate115inter7));
  inv1  gate891(.a(G383), .O(gate115inter8));
  nand2 gate892(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate893(.a(s_49), .b(gate115inter3), .O(gate115inter10));
  nor2  gate894(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate895(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate896(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate589(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate590(.a(gate116inter0), .b(s_6), .O(gate116inter1));
  and2  gate591(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate592(.a(s_6), .O(gate116inter3));
  inv1  gate593(.a(s_7), .O(gate116inter4));
  nand2 gate594(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate595(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate596(.a(G384), .O(gate116inter7));
  inv1  gate597(.a(G385), .O(gate116inter8));
  nand2 gate598(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate599(.a(s_7), .b(gate116inter3), .O(gate116inter10));
  nor2  gate600(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate601(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate602(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate2773(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2774(.a(gate117inter0), .b(s_318), .O(gate117inter1));
  and2  gate2775(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2776(.a(s_318), .O(gate117inter3));
  inv1  gate2777(.a(s_319), .O(gate117inter4));
  nand2 gate2778(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2779(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2780(.a(G386), .O(gate117inter7));
  inv1  gate2781(.a(G387), .O(gate117inter8));
  nand2 gate2782(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2783(.a(s_319), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2784(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2785(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2786(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1555(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1556(.a(gate119inter0), .b(s_144), .O(gate119inter1));
  and2  gate1557(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1558(.a(s_144), .O(gate119inter3));
  inv1  gate1559(.a(s_145), .O(gate119inter4));
  nand2 gate1560(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1561(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1562(.a(G390), .O(gate119inter7));
  inv1  gate1563(.a(G391), .O(gate119inter8));
  nand2 gate1564(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1565(.a(s_145), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1566(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1567(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1568(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2675(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2676(.a(gate122inter0), .b(s_304), .O(gate122inter1));
  and2  gate2677(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2678(.a(s_304), .O(gate122inter3));
  inv1  gate2679(.a(s_305), .O(gate122inter4));
  nand2 gate2680(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2681(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2682(.a(G396), .O(gate122inter7));
  inv1  gate2683(.a(G397), .O(gate122inter8));
  nand2 gate2684(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2685(.a(s_305), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2686(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2687(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2688(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate995(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate996(.a(gate126inter0), .b(s_64), .O(gate126inter1));
  and2  gate997(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate998(.a(s_64), .O(gate126inter3));
  inv1  gate999(.a(s_65), .O(gate126inter4));
  nand2 gate1000(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1001(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1002(.a(G404), .O(gate126inter7));
  inv1  gate1003(.a(G405), .O(gate126inter8));
  nand2 gate1004(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1005(.a(s_65), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1006(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1007(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1008(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate813(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate814(.a(gate131inter0), .b(s_38), .O(gate131inter1));
  and2  gate815(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate816(.a(s_38), .O(gate131inter3));
  inv1  gate817(.a(s_39), .O(gate131inter4));
  nand2 gate818(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate819(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate820(.a(G414), .O(gate131inter7));
  inv1  gate821(.a(G415), .O(gate131inter8));
  nand2 gate822(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate823(.a(s_39), .b(gate131inter3), .O(gate131inter10));
  nor2  gate824(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate825(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate826(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1079(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1080(.a(gate132inter0), .b(s_76), .O(gate132inter1));
  and2  gate1081(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1082(.a(s_76), .O(gate132inter3));
  inv1  gate1083(.a(s_77), .O(gate132inter4));
  nand2 gate1084(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1085(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1086(.a(G416), .O(gate132inter7));
  inv1  gate1087(.a(G417), .O(gate132inter8));
  nand2 gate1088(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1089(.a(s_77), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1090(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1091(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1092(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1625(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1626(.a(gate136inter0), .b(s_154), .O(gate136inter1));
  and2  gate1627(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1628(.a(s_154), .O(gate136inter3));
  inv1  gate1629(.a(s_155), .O(gate136inter4));
  nand2 gate1630(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1631(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1632(.a(G424), .O(gate136inter7));
  inv1  gate1633(.a(G425), .O(gate136inter8));
  nand2 gate1634(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1635(.a(s_155), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1636(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1637(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1638(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2563(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2564(.a(gate137inter0), .b(s_288), .O(gate137inter1));
  and2  gate2565(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2566(.a(s_288), .O(gate137inter3));
  inv1  gate2567(.a(s_289), .O(gate137inter4));
  nand2 gate2568(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2569(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2570(.a(G426), .O(gate137inter7));
  inv1  gate2571(.a(G429), .O(gate137inter8));
  nand2 gate2572(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2573(.a(s_289), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2574(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2575(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2576(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2297(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2298(.a(gate140inter0), .b(s_250), .O(gate140inter1));
  and2  gate2299(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2300(.a(s_250), .O(gate140inter3));
  inv1  gate2301(.a(s_251), .O(gate140inter4));
  nand2 gate2302(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2303(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2304(.a(G444), .O(gate140inter7));
  inv1  gate2305(.a(G447), .O(gate140inter8));
  nand2 gate2306(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2307(.a(s_251), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2308(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2309(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2310(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1765(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1766(.a(gate142inter0), .b(s_174), .O(gate142inter1));
  and2  gate1767(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1768(.a(s_174), .O(gate142inter3));
  inv1  gate1769(.a(s_175), .O(gate142inter4));
  nand2 gate1770(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1771(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1772(.a(G456), .O(gate142inter7));
  inv1  gate1773(.a(G459), .O(gate142inter8));
  nand2 gate1774(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1775(.a(s_175), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1776(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1777(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1778(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2703(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2704(.a(gate148inter0), .b(s_308), .O(gate148inter1));
  and2  gate2705(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2706(.a(s_308), .O(gate148inter3));
  inv1  gate2707(.a(s_309), .O(gate148inter4));
  nand2 gate2708(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2709(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2710(.a(G492), .O(gate148inter7));
  inv1  gate2711(.a(G495), .O(gate148inter8));
  nand2 gate2712(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2713(.a(s_309), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2714(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2715(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2716(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1415(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1416(.a(gate150inter0), .b(s_124), .O(gate150inter1));
  and2  gate1417(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1418(.a(s_124), .O(gate150inter3));
  inv1  gate1419(.a(s_125), .O(gate150inter4));
  nand2 gate1420(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1421(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1422(.a(G504), .O(gate150inter7));
  inv1  gate1423(.a(G507), .O(gate150inter8));
  nand2 gate1424(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1425(.a(s_125), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1426(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1427(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1428(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2745(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2746(.a(gate151inter0), .b(s_314), .O(gate151inter1));
  and2  gate2747(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2748(.a(s_314), .O(gate151inter3));
  inv1  gate2749(.a(s_315), .O(gate151inter4));
  nand2 gate2750(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2751(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2752(.a(G510), .O(gate151inter7));
  inv1  gate2753(.a(G513), .O(gate151inter8));
  nand2 gate2754(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2755(.a(s_315), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2756(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2757(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2758(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate841(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate842(.a(gate154inter0), .b(s_42), .O(gate154inter1));
  and2  gate843(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate844(.a(s_42), .O(gate154inter3));
  inv1  gate845(.a(s_43), .O(gate154inter4));
  nand2 gate846(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate847(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate848(.a(G429), .O(gate154inter7));
  inv1  gate849(.a(G522), .O(gate154inter8));
  nand2 gate850(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate851(.a(s_43), .b(gate154inter3), .O(gate154inter10));
  nor2  gate852(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate853(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate854(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2815(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2816(.a(gate157inter0), .b(s_324), .O(gate157inter1));
  and2  gate2817(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2818(.a(s_324), .O(gate157inter3));
  inv1  gate2819(.a(s_325), .O(gate157inter4));
  nand2 gate2820(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2821(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2822(.a(G438), .O(gate157inter7));
  inv1  gate2823(.a(G528), .O(gate157inter8));
  nand2 gate2824(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2825(.a(s_325), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2826(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2827(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2828(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1023(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1024(.a(gate158inter0), .b(s_68), .O(gate158inter1));
  and2  gate1025(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1026(.a(s_68), .O(gate158inter3));
  inv1  gate1027(.a(s_69), .O(gate158inter4));
  nand2 gate1028(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1029(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1030(.a(G441), .O(gate158inter7));
  inv1  gate1031(.a(G528), .O(gate158inter8));
  nand2 gate1032(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1033(.a(s_69), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1034(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1035(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1036(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate2899(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2900(.a(gate160inter0), .b(s_336), .O(gate160inter1));
  and2  gate2901(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2902(.a(s_336), .O(gate160inter3));
  inv1  gate2903(.a(s_337), .O(gate160inter4));
  nand2 gate2904(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2905(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2906(.a(G447), .O(gate160inter7));
  inv1  gate2907(.a(G531), .O(gate160inter8));
  nand2 gate2908(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2909(.a(s_337), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2910(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2911(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2912(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate2059(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2060(.a(gate161inter0), .b(s_216), .O(gate161inter1));
  and2  gate2061(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2062(.a(s_216), .O(gate161inter3));
  inv1  gate2063(.a(s_217), .O(gate161inter4));
  nand2 gate2064(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2065(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2066(.a(G450), .O(gate161inter7));
  inv1  gate2067(.a(G534), .O(gate161inter8));
  nand2 gate2068(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2069(.a(s_217), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2070(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2071(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2072(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2213(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2214(.a(gate167inter0), .b(s_238), .O(gate167inter1));
  and2  gate2215(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2216(.a(s_238), .O(gate167inter3));
  inv1  gate2217(.a(s_239), .O(gate167inter4));
  nand2 gate2218(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2219(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2220(.a(G468), .O(gate167inter7));
  inv1  gate2221(.a(G543), .O(gate167inter8));
  nand2 gate2222(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2223(.a(s_239), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2224(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2225(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2226(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate687(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate688(.a(gate168inter0), .b(s_20), .O(gate168inter1));
  and2  gate689(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate690(.a(s_20), .O(gate168inter3));
  inv1  gate691(.a(s_21), .O(gate168inter4));
  nand2 gate692(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate693(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate694(.a(G471), .O(gate168inter7));
  inv1  gate695(.a(G543), .O(gate168inter8));
  nand2 gate696(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate697(.a(s_21), .b(gate168inter3), .O(gate168inter10));
  nor2  gate698(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate699(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate700(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1121(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1122(.a(gate169inter0), .b(s_82), .O(gate169inter1));
  and2  gate1123(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1124(.a(s_82), .O(gate169inter3));
  inv1  gate1125(.a(s_83), .O(gate169inter4));
  nand2 gate1126(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1127(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1128(.a(G474), .O(gate169inter7));
  inv1  gate1129(.a(G546), .O(gate169inter8));
  nand2 gate1130(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1131(.a(s_83), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1132(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1133(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1134(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1401(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1402(.a(gate175inter0), .b(s_122), .O(gate175inter1));
  and2  gate1403(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1404(.a(s_122), .O(gate175inter3));
  inv1  gate1405(.a(s_123), .O(gate175inter4));
  nand2 gate1406(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1407(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1408(.a(G492), .O(gate175inter7));
  inv1  gate1409(.a(G555), .O(gate175inter8));
  nand2 gate1410(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1411(.a(s_123), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1412(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1413(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1414(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate2311(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2312(.a(gate176inter0), .b(s_252), .O(gate176inter1));
  and2  gate2313(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2314(.a(s_252), .O(gate176inter3));
  inv1  gate2315(.a(s_253), .O(gate176inter4));
  nand2 gate2316(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2317(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2318(.a(G495), .O(gate176inter7));
  inv1  gate2319(.a(G555), .O(gate176inter8));
  nand2 gate2320(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2321(.a(s_253), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2322(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2323(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2324(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1905(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1906(.a(gate178inter0), .b(s_194), .O(gate178inter1));
  and2  gate1907(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1908(.a(s_194), .O(gate178inter3));
  inv1  gate1909(.a(s_195), .O(gate178inter4));
  nand2 gate1910(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1911(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1912(.a(G501), .O(gate178inter7));
  inv1  gate1913(.a(G558), .O(gate178inter8));
  nand2 gate1914(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1915(.a(s_195), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1916(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1917(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1918(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2689(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2690(.a(gate180inter0), .b(s_306), .O(gate180inter1));
  and2  gate2691(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2692(.a(s_306), .O(gate180inter3));
  inv1  gate2693(.a(s_307), .O(gate180inter4));
  nand2 gate2694(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2695(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2696(.a(G507), .O(gate180inter7));
  inv1  gate2697(.a(G561), .O(gate180inter8));
  nand2 gate2698(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2699(.a(s_307), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2700(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2701(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2702(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2409(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2410(.a(gate182inter0), .b(s_266), .O(gate182inter1));
  and2  gate2411(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2412(.a(s_266), .O(gate182inter3));
  inv1  gate2413(.a(s_267), .O(gate182inter4));
  nand2 gate2414(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2415(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2416(.a(G513), .O(gate182inter7));
  inv1  gate2417(.a(G564), .O(gate182inter8));
  nand2 gate2418(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2419(.a(s_267), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2420(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2421(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2422(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate827(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate828(.a(gate184inter0), .b(s_40), .O(gate184inter1));
  and2  gate829(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate830(.a(s_40), .O(gate184inter3));
  inv1  gate831(.a(s_41), .O(gate184inter4));
  nand2 gate832(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate833(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate834(.a(G519), .O(gate184inter7));
  inv1  gate835(.a(G567), .O(gate184inter8));
  nand2 gate836(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate837(.a(s_41), .b(gate184inter3), .O(gate184inter10));
  nor2  gate838(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate839(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate840(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1709(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1710(.a(gate186inter0), .b(s_166), .O(gate186inter1));
  and2  gate1711(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1712(.a(s_166), .O(gate186inter3));
  inv1  gate1713(.a(s_167), .O(gate186inter4));
  nand2 gate1714(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1715(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1716(.a(G572), .O(gate186inter7));
  inv1  gate1717(.a(G573), .O(gate186inter8));
  nand2 gate1718(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1719(.a(s_167), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1720(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1721(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1722(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate2157(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2158(.a(gate187inter0), .b(s_230), .O(gate187inter1));
  and2  gate2159(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2160(.a(s_230), .O(gate187inter3));
  inv1  gate2161(.a(s_231), .O(gate187inter4));
  nand2 gate2162(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2163(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2164(.a(G574), .O(gate187inter7));
  inv1  gate2165(.a(G575), .O(gate187inter8));
  nand2 gate2166(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2167(.a(s_231), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2168(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2169(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2170(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1205(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1206(.a(gate189inter0), .b(s_94), .O(gate189inter1));
  and2  gate1207(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1208(.a(s_94), .O(gate189inter3));
  inv1  gate1209(.a(s_95), .O(gate189inter4));
  nand2 gate1210(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1211(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1212(.a(G578), .O(gate189inter7));
  inv1  gate1213(.a(G579), .O(gate189inter8));
  nand2 gate1214(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1215(.a(s_95), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1216(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1217(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1218(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate967(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate968(.a(gate192inter0), .b(s_60), .O(gate192inter1));
  and2  gate969(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate970(.a(s_60), .O(gate192inter3));
  inv1  gate971(.a(s_61), .O(gate192inter4));
  nand2 gate972(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate973(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate974(.a(G584), .O(gate192inter7));
  inv1  gate975(.a(G585), .O(gate192inter8));
  nand2 gate976(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate977(.a(s_61), .b(gate192inter3), .O(gate192inter10));
  nor2  gate978(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate979(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate980(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1891(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1892(.a(gate197inter0), .b(s_192), .O(gate197inter1));
  and2  gate1893(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1894(.a(s_192), .O(gate197inter3));
  inv1  gate1895(.a(s_193), .O(gate197inter4));
  nand2 gate1896(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1897(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1898(.a(G594), .O(gate197inter7));
  inv1  gate1899(.a(G595), .O(gate197inter8));
  nand2 gate1900(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1901(.a(s_193), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1902(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1903(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1904(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1849(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1850(.a(gate200inter0), .b(s_186), .O(gate200inter1));
  and2  gate1851(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1852(.a(s_186), .O(gate200inter3));
  inv1  gate1853(.a(s_187), .O(gate200inter4));
  nand2 gate1854(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1855(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1856(.a(G600), .O(gate200inter7));
  inv1  gate1857(.a(G601), .O(gate200inter8));
  nand2 gate1858(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1859(.a(s_187), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1860(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1861(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1862(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2885(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2886(.a(gate205inter0), .b(s_334), .O(gate205inter1));
  and2  gate2887(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2888(.a(s_334), .O(gate205inter3));
  inv1  gate2889(.a(s_335), .O(gate205inter4));
  nand2 gate2890(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2891(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2892(.a(G622), .O(gate205inter7));
  inv1  gate2893(.a(G627), .O(gate205inter8));
  nand2 gate2894(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2895(.a(s_335), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2896(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2897(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2898(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate715(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate716(.a(gate206inter0), .b(s_24), .O(gate206inter1));
  and2  gate717(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate718(.a(s_24), .O(gate206inter3));
  inv1  gate719(.a(s_25), .O(gate206inter4));
  nand2 gate720(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate721(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate722(.a(G632), .O(gate206inter7));
  inv1  gate723(.a(G637), .O(gate206inter8));
  nand2 gate724(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate725(.a(s_25), .b(gate206inter3), .O(gate206inter10));
  nor2  gate726(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate727(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate728(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1065(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1066(.a(gate212inter0), .b(s_74), .O(gate212inter1));
  and2  gate1067(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1068(.a(s_74), .O(gate212inter3));
  inv1  gate1069(.a(s_75), .O(gate212inter4));
  nand2 gate1070(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1071(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1072(.a(G617), .O(gate212inter7));
  inv1  gate1073(.a(G669), .O(gate212inter8));
  nand2 gate1074(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1075(.a(s_75), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1076(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1077(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1078(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1681(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1682(.a(gate213inter0), .b(s_162), .O(gate213inter1));
  and2  gate1683(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1684(.a(s_162), .O(gate213inter3));
  inv1  gate1685(.a(s_163), .O(gate213inter4));
  nand2 gate1686(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1687(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1688(.a(G602), .O(gate213inter7));
  inv1  gate1689(.a(G672), .O(gate213inter8));
  nand2 gate1690(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1691(.a(s_163), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1692(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1693(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1694(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1989(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1990(.a(gate214inter0), .b(s_206), .O(gate214inter1));
  and2  gate1991(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1992(.a(s_206), .O(gate214inter3));
  inv1  gate1993(.a(s_207), .O(gate214inter4));
  nand2 gate1994(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1995(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1996(.a(G612), .O(gate214inter7));
  inv1  gate1997(.a(G672), .O(gate214inter8));
  nand2 gate1998(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1999(.a(s_207), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2000(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2001(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2002(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1485(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1486(.a(gate217inter0), .b(s_134), .O(gate217inter1));
  and2  gate1487(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1488(.a(s_134), .O(gate217inter3));
  inv1  gate1489(.a(s_135), .O(gate217inter4));
  nand2 gate1490(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1491(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1492(.a(G622), .O(gate217inter7));
  inv1  gate1493(.a(G678), .O(gate217inter8));
  nand2 gate1494(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1495(.a(s_135), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1496(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1497(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1498(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1429(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1430(.a(gate219inter0), .b(s_126), .O(gate219inter1));
  and2  gate1431(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1432(.a(s_126), .O(gate219inter3));
  inv1  gate1433(.a(s_127), .O(gate219inter4));
  nand2 gate1434(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1435(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1436(.a(G632), .O(gate219inter7));
  inv1  gate1437(.a(G681), .O(gate219inter8));
  nand2 gate1438(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1439(.a(s_127), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1440(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1441(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1442(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2843(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2844(.a(gate220inter0), .b(s_328), .O(gate220inter1));
  and2  gate2845(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2846(.a(s_328), .O(gate220inter3));
  inv1  gate2847(.a(s_329), .O(gate220inter4));
  nand2 gate2848(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2849(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2850(.a(G637), .O(gate220inter7));
  inv1  gate2851(.a(G681), .O(gate220inter8));
  nand2 gate2852(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2853(.a(s_329), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2854(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2855(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2856(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1331(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1332(.a(gate221inter0), .b(s_112), .O(gate221inter1));
  and2  gate1333(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1334(.a(s_112), .O(gate221inter3));
  inv1  gate1335(.a(s_113), .O(gate221inter4));
  nand2 gate1336(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1337(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1338(.a(G622), .O(gate221inter7));
  inv1  gate1339(.a(G684), .O(gate221inter8));
  nand2 gate1340(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1341(.a(s_113), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1342(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1343(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1344(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate2927(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2928(.a(gate222inter0), .b(s_340), .O(gate222inter1));
  and2  gate2929(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2930(.a(s_340), .O(gate222inter3));
  inv1  gate2931(.a(s_341), .O(gate222inter4));
  nand2 gate2932(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2933(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2934(.a(G632), .O(gate222inter7));
  inv1  gate2935(.a(G684), .O(gate222inter8));
  nand2 gate2936(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2937(.a(s_341), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2938(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2939(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2940(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2381(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2382(.a(gate225inter0), .b(s_262), .O(gate225inter1));
  and2  gate2383(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2384(.a(s_262), .O(gate225inter3));
  inv1  gate2385(.a(s_263), .O(gate225inter4));
  nand2 gate2386(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2387(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2388(.a(G690), .O(gate225inter7));
  inv1  gate2389(.a(G691), .O(gate225inter8));
  nand2 gate2390(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2391(.a(s_263), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2392(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2393(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2394(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate617(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate618(.a(gate226inter0), .b(s_10), .O(gate226inter1));
  and2  gate619(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate620(.a(s_10), .O(gate226inter3));
  inv1  gate621(.a(s_11), .O(gate226inter4));
  nand2 gate622(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate623(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate624(.a(G692), .O(gate226inter7));
  inv1  gate625(.a(G693), .O(gate226inter8));
  nand2 gate626(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate627(.a(s_11), .b(gate226inter3), .O(gate226inter10));
  nor2  gate628(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate629(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate630(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2283(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2284(.a(gate229inter0), .b(s_248), .O(gate229inter1));
  and2  gate2285(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2286(.a(s_248), .O(gate229inter3));
  inv1  gate2287(.a(s_249), .O(gate229inter4));
  nand2 gate2288(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2289(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2290(.a(G698), .O(gate229inter7));
  inv1  gate2291(.a(G699), .O(gate229inter8));
  nand2 gate2292(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2293(.a(s_249), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2294(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2295(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2296(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate2339(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2340(.a(gate230inter0), .b(s_256), .O(gate230inter1));
  and2  gate2341(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2342(.a(s_256), .O(gate230inter3));
  inv1  gate2343(.a(s_257), .O(gate230inter4));
  nand2 gate2344(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2345(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2346(.a(G700), .O(gate230inter7));
  inv1  gate2347(.a(G701), .O(gate230inter8));
  nand2 gate2348(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2349(.a(s_257), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2350(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2351(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2352(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2857(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2858(.a(gate231inter0), .b(s_330), .O(gate231inter1));
  and2  gate2859(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2860(.a(s_330), .O(gate231inter3));
  inv1  gate2861(.a(s_331), .O(gate231inter4));
  nand2 gate2862(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2863(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2864(.a(G702), .O(gate231inter7));
  inv1  gate2865(.a(G703), .O(gate231inter8));
  nand2 gate2866(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2867(.a(s_331), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2868(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2869(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2870(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1289(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1290(.a(gate232inter0), .b(s_106), .O(gate232inter1));
  and2  gate1291(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1292(.a(s_106), .O(gate232inter3));
  inv1  gate1293(.a(s_107), .O(gate232inter4));
  nand2 gate1294(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1295(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1296(.a(G704), .O(gate232inter7));
  inv1  gate1297(.a(G705), .O(gate232inter8));
  nand2 gate1298(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1299(.a(s_107), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1300(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1301(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1302(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2661(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2662(.a(gate234inter0), .b(s_302), .O(gate234inter1));
  and2  gate2663(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2664(.a(s_302), .O(gate234inter3));
  inv1  gate2665(.a(s_303), .O(gate234inter4));
  nand2 gate2666(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2667(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2668(.a(G245), .O(gate234inter7));
  inv1  gate2669(.a(G721), .O(gate234inter8));
  nand2 gate2670(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2671(.a(s_303), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2672(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2673(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2674(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2227(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2228(.a(gate235inter0), .b(s_240), .O(gate235inter1));
  and2  gate2229(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2230(.a(s_240), .O(gate235inter3));
  inv1  gate2231(.a(s_241), .O(gate235inter4));
  nand2 gate2232(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2233(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2234(.a(G248), .O(gate235inter7));
  inv1  gate2235(.a(G724), .O(gate235inter8));
  nand2 gate2236(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2237(.a(s_241), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2238(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2239(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2240(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate1051(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1052(.a(gate236inter0), .b(s_72), .O(gate236inter1));
  and2  gate1053(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1054(.a(s_72), .O(gate236inter3));
  inv1  gate1055(.a(s_73), .O(gate236inter4));
  nand2 gate1056(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1057(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1058(.a(G251), .O(gate236inter7));
  inv1  gate1059(.a(G727), .O(gate236inter8));
  nand2 gate1060(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1061(.a(s_73), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1062(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1063(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1064(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate2017(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2018(.a(gate237inter0), .b(s_210), .O(gate237inter1));
  and2  gate2019(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2020(.a(s_210), .O(gate237inter3));
  inv1  gate2021(.a(s_211), .O(gate237inter4));
  nand2 gate2022(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2023(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2024(.a(G254), .O(gate237inter7));
  inv1  gate2025(.a(G706), .O(gate237inter8));
  nand2 gate2026(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2027(.a(s_211), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2028(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2029(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2030(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate757(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate758(.a(gate239inter0), .b(s_30), .O(gate239inter1));
  and2  gate759(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate760(.a(s_30), .O(gate239inter3));
  inv1  gate761(.a(s_31), .O(gate239inter4));
  nand2 gate762(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate763(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate764(.a(G260), .O(gate239inter7));
  inv1  gate765(.a(G712), .O(gate239inter8));
  nand2 gate766(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate767(.a(s_31), .b(gate239inter3), .O(gate239inter10));
  nor2  gate768(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate769(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate770(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2787(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2788(.a(gate244inter0), .b(s_320), .O(gate244inter1));
  and2  gate2789(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2790(.a(s_320), .O(gate244inter3));
  inv1  gate2791(.a(s_321), .O(gate244inter4));
  nand2 gate2792(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2793(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2794(.a(G721), .O(gate244inter7));
  inv1  gate2795(.a(G733), .O(gate244inter8));
  nand2 gate2796(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2797(.a(s_321), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2798(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2799(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2800(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2325(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2326(.a(gate249inter0), .b(s_254), .O(gate249inter1));
  and2  gate2327(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2328(.a(s_254), .O(gate249inter3));
  inv1  gate2329(.a(s_255), .O(gate249inter4));
  nand2 gate2330(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2331(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2332(.a(G254), .O(gate249inter7));
  inv1  gate2333(.a(G742), .O(gate249inter8));
  nand2 gate2334(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2335(.a(s_255), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2336(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2337(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2338(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate729(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate730(.a(gate251inter0), .b(s_26), .O(gate251inter1));
  and2  gate731(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate732(.a(s_26), .O(gate251inter3));
  inv1  gate733(.a(s_27), .O(gate251inter4));
  nand2 gate734(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate735(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate736(.a(G257), .O(gate251inter7));
  inv1  gate737(.a(G745), .O(gate251inter8));
  nand2 gate738(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate739(.a(s_27), .b(gate251inter3), .O(gate251inter10));
  nor2  gate740(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate741(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate742(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate785(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate786(.a(gate255inter0), .b(s_34), .O(gate255inter1));
  and2  gate787(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate788(.a(s_34), .O(gate255inter3));
  inv1  gate789(.a(s_35), .O(gate255inter4));
  nand2 gate790(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate791(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate792(.a(G263), .O(gate255inter7));
  inv1  gate793(.a(G751), .O(gate255inter8));
  nand2 gate794(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate795(.a(s_35), .b(gate255inter3), .O(gate255inter10));
  nor2  gate796(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate797(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate798(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate799(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate800(.a(gate256inter0), .b(s_36), .O(gate256inter1));
  and2  gate801(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate802(.a(s_36), .O(gate256inter3));
  inv1  gate803(.a(s_37), .O(gate256inter4));
  nand2 gate804(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate805(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate806(.a(G715), .O(gate256inter7));
  inv1  gate807(.a(G751), .O(gate256inter8));
  nand2 gate808(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate809(.a(s_37), .b(gate256inter3), .O(gate256inter10));
  nor2  gate810(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate811(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate812(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1093(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1094(.a(gate258inter0), .b(s_78), .O(gate258inter1));
  and2  gate1095(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1096(.a(s_78), .O(gate258inter3));
  inv1  gate1097(.a(s_79), .O(gate258inter4));
  nand2 gate1098(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1099(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1100(.a(G756), .O(gate258inter7));
  inv1  gate1101(.a(G757), .O(gate258inter8));
  nand2 gate1102(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1103(.a(s_79), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1104(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1105(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1106(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1779(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1780(.a(gate259inter0), .b(s_176), .O(gate259inter1));
  and2  gate1781(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1782(.a(s_176), .O(gate259inter3));
  inv1  gate1783(.a(s_177), .O(gate259inter4));
  nand2 gate1784(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1785(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1786(.a(G758), .O(gate259inter7));
  inv1  gate1787(.a(G759), .O(gate259inter8));
  nand2 gate1788(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1789(.a(s_177), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1790(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1791(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1792(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2717(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2718(.a(gate261inter0), .b(s_310), .O(gate261inter1));
  and2  gate2719(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2720(.a(s_310), .O(gate261inter3));
  inv1  gate2721(.a(s_311), .O(gate261inter4));
  nand2 gate2722(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2723(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2724(.a(G762), .O(gate261inter7));
  inv1  gate2725(.a(G763), .O(gate261inter8));
  nand2 gate2726(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2727(.a(s_311), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2728(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2729(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2730(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1345(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1346(.a(gate265inter0), .b(s_114), .O(gate265inter1));
  and2  gate1347(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1348(.a(s_114), .O(gate265inter3));
  inv1  gate1349(.a(s_115), .O(gate265inter4));
  nand2 gate1350(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1351(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1352(.a(G642), .O(gate265inter7));
  inv1  gate1353(.a(G770), .O(gate265inter8));
  nand2 gate1354(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1355(.a(s_115), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1356(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1357(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1358(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate743(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate744(.a(gate267inter0), .b(s_28), .O(gate267inter1));
  and2  gate745(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate746(.a(s_28), .O(gate267inter3));
  inv1  gate747(.a(s_29), .O(gate267inter4));
  nand2 gate748(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate749(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate750(.a(G648), .O(gate267inter7));
  inv1  gate751(.a(G776), .O(gate267inter8));
  nand2 gate752(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate753(.a(s_29), .b(gate267inter3), .O(gate267inter10));
  nor2  gate754(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate755(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate756(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate547(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate548(.a(gate270inter0), .b(s_0), .O(gate270inter1));
  and2  gate549(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate550(.a(s_0), .O(gate270inter3));
  inv1  gate551(.a(s_1), .O(gate270inter4));
  nand2 gate552(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate553(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate554(.a(G657), .O(gate270inter7));
  inv1  gate555(.a(G785), .O(gate270inter8));
  nand2 gate556(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate557(.a(s_1), .b(gate270inter3), .O(gate270inter10));
  nor2  gate558(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate559(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate560(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1471(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1472(.a(gate279inter0), .b(s_132), .O(gate279inter1));
  and2  gate1473(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1474(.a(s_132), .O(gate279inter3));
  inv1  gate1475(.a(s_133), .O(gate279inter4));
  nand2 gate1476(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1477(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1478(.a(G651), .O(gate279inter7));
  inv1  gate1479(.a(G803), .O(gate279inter8));
  nand2 gate1480(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1481(.a(s_133), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1482(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1483(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1484(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate2731(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2732(.a(gate280inter0), .b(s_312), .O(gate280inter1));
  and2  gate2733(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2734(.a(s_312), .O(gate280inter3));
  inv1  gate2735(.a(s_313), .O(gate280inter4));
  nand2 gate2736(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2737(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2738(.a(G779), .O(gate280inter7));
  inv1  gate2739(.a(G803), .O(gate280inter8));
  nand2 gate2740(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2741(.a(s_313), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2742(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2743(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2744(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1877(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1878(.a(gate281inter0), .b(s_190), .O(gate281inter1));
  and2  gate1879(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1880(.a(s_190), .O(gate281inter3));
  inv1  gate1881(.a(s_191), .O(gate281inter4));
  nand2 gate1882(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1883(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1884(.a(G654), .O(gate281inter7));
  inv1  gate1885(.a(G806), .O(gate281inter8));
  nand2 gate1886(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1887(.a(s_191), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1888(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1889(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1890(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2493(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2494(.a(gate286inter0), .b(s_278), .O(gate286inter1));
  and2  gate2495(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2496(.a(s_278), .O(gate286inter3));
  inv1  gate2497(.a(s_279), .O(gate286inter4));
  nand2 gate2498(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2499(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2500(.a(G788), .O(gate286inter7));
  inv1  gate2501(.a(G812), .O(gate286inter8));
  nand2 gate2502(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2503(.a(s_279), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2504(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2505(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2506(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2465(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2466(.a(gate288inter0), .b(s_274), .O(gate288inter1));
  and2  gate2467(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2468(.a(s_274), .O(gate288inter3));
  inv1  gate2469(.a(s_275), .O(gate288inter4));
  nand2 gate2470(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2471(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2472(.a(G791), .O(gate288inter7));
  inv1  gate2473(.a(G815), .O(gate288inter8));
  nand2 gate2474(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2475(.a(s_275), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2476(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2477(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2478(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate2619(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2620(.a(gate289inter0), .b(s_296), .O(gate289inter1));
  and2  gate2621(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2622(.a(s_296), .O(gate289inter3));
  inv1  gate2623(.a(s_297), .O(gate289inter4));
  nand2 gate2624(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2625(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2626(.a(G818), .O(gate289inter7));
  inv1  gate2627(.a(G819), .O(gate289inter8));
  nand2 gate2628(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2629(.a(s_297), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2630(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2631(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2632(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate869(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate870(.a(gate290inter0), .b(s_46), .O(gate290inter1));
  and2  gate871(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate872(.a(s_46), .O(gate290inter3));
  inv1  gate873(.a(s_47), .O(gate290inter4));
  nand2 gate874(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate875(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate876(.a(G820), .O(gate290inter7));
  inv1  gate877(.a(G821), .O(gate290inter8));
  nand2 gate878(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate879(.a(s_47), .b(gate290inter3), .O(gate290inter10));
  nor2  gate880(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate881(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate882(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1149(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1150(.a(gate292inter0), .b(s_86), .O(gate292inter1));
  and2  gate1151(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1152(.a(s_86), .O(gate292inter3));
  inv1  gate1153(.a(s_87), .O(gate292inter4));
  nand2 gate1154(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1155(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1156(.a(G824), .O(gate292inter7));
  inv1  gate1157(.a(G825), .O(gate292inter8));
  nand2 gate1158(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1159(.a(s_87), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1160(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1161(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1162(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate561(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate562(.a(gate293inter0), .b(s_2), .O(gate293inter1));
  and2  gate563(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate564(.a(s_2), .O(gate293inter3));
  inv1  gate565(.a(s_3), .O(gate293inter4));
  nand2 gate566(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate567(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate568(.a(G828), .O(gate293inter7));
  inv1  gate569(.a(G829), .O(gate293inter8));
  nand2 gate570(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate571(.a(s_3), .b(gate293inter3), .O(gate293inter10));
  nor2  gate572(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate573(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate574(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1975(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1976(.a(gate387inter0), .b(s_204), .O(gate387inter1));
  and2  gate1977(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1978(.a(s_204), .O(gate387inter3));
  inv1  gate1979(.a(s_205), .O(gate387inter4));
  nand2 gate1980(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1981(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1982(.a(G1), .O(gate387inter7));
  inv1  gate1983(.a(G1036), .O(gate387inter8));
  nand2 gate1984(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1985(.a(s_205), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1986(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1987(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1988(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2115(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2116(.a(gate389inter0), .b(s_224), .O(gate389inter1));
  and2  gate2117(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2118(.a(s_224), .O(gate389inter3));
  inv1  gate2119(.a(s_225), .O(gate389inter4));
  nand2 gate2120(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2121(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2122(.a(G3), .O(gate389inter7));
  inv1  gate2123(.a(G1042), .O(gate389inter8));
  nand2 gate2124(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2125(.a(s_225), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2126(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2127(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2128(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2073(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2074(.a(gate393inter0), .b(s_218), .O(gate393inter1));
  and2  gate2075(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2076(.a(s_218), .O(gate393inter3));
  inv1  gate2077(.a(s_219), .O(gate393inter4));
  nand2 gate2078(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2079(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2080(.a(G7), .O(gate393inter7));
  inv1  gate2081(.a(G1054), .O(gate393inter8));
  nand2 gate2082(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2083(.a(s_219), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2084(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2085(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2086(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1359(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1360(.a(gate395inter0), .b(s_116), .O(gate395inter1));
  and2  gate1361(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1362(.a(s_116), .O(gate395inter3));
  inv1  gate1363(.a(s_117), .O(gate395inter4));
  nand2 gate1364(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1365(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1366(.a(G9), .O(gate395inter7));
  inv1  gate1367(.a(G1060), .O(gate395inter8));
  nand2 gate1368(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1369(.a(s_117), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1370(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1371(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1372(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1443(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1444(.a(gate396inter0), .b(s_128), .O(gate396inter1));
  and2  gate1445(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1446(.a(s_128), .O(gate396inter3));
  inv1  gate1447(.a(s_129), .O(gate396inter4));
  nand2 gate1448(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1449(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1450(.a(G10), .O(gate396inter7));
  inv1  gate1451(.a(G1063), .O(gate396inter8));
  nand2 gate1452(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1453(.a(s_129), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1454(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1455(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1456(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1177(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1178(.a(gate398inter0), .b(s_90), .O(gate398inter1));
  and2  gate1179(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1180(.a(s_90), .O(gate398inter3));
  inv1  gate1181(.a(s_91), .O(gate398inter4));
  nand2 gate1182(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1183(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1184(.a(G12), .O(gate398inter7));
  inv1  gate1185(.a(G1069), .O(gate398inter8));
  nand2 gate1186(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1187(.a(s_91), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1188(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1189(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1190(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate953(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate954(.a(gate399inter0), .b(s_58), .O(gate399inter1));
  and2  gate955(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate956(.a(s_58), .O(gate399inter3));
  inv1  gate957(.a(s_59), .O(gate399inter4));
  nand2 gate958(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate959(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate960(.a(G13), .O(gate399inter7));
  inv1  gate961(.a(G1072), .O(gate399inter8));
  nand2 gate962(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate963(.a(s_59), .b(gate399inter3), .O(gate399inter10));
  nor2  gate964(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate965(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate966(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate2129(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2130(.a(gate400inter0), .b(s_226), .O(gate400inter1));
  and2  gate2131(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2132(.a(s_226), .O(gate400inter3));
  inv1  gate2133(.a(s_227), .O(gate400inter4));
  nand2 gate2134(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2135(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2136(.a(G14), .O(gate400inter7));
  inv1  gate2137(.a(G1075), .O(gate400inter8));
  nand2 gate2138(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2139(.a(s_227), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2140(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2141(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2142(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate575(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate576(.a(gate401inter0), .b(s_4), .O(gate401inter1));
  and2  gate577(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate578(.a(s_4), .O(gate401inter3));
  inv1  gate579(.a(s_5), .O(gate401inter4));
  nand2 gate580(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate581(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate582(.a(G15), .O(gate401inter7));
  inv1  gate583(.a(G1078), .O(gate401inter8));
  nand2 gate584(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate585(.a(s_5), .b(gate401inter3), .O(gate401inter10));
  nor2  gate586(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate587(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate588(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1695(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1696(.a(gate402inter0), .b(s_164), .O(gate402inter1));
  and2  gate1697(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1698(.a(s_164), .O(gate402inter3));
  inv1  gate1699(.a(s_165), .O(gate402inter4));
  nand2 gate1700(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1701(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1702(.a(G16), .O(gate402inter7));
  inv1  gate1703(.a(G1081), .O(gate402inter8));
  nand2 gate1704(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1705(.a(s_165), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1706(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1707(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1708(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate2003(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2004(.a(gate403inter0), .b(s_208), .O(gate403inter1));
  and2  gate2005(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2006(.a(s_208), .O(gate403inter3));
  inv1  gate2007(.a(s_209), .O(gate403inter4));
  nand2 gate2008(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2009(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2010(.a(G17), .O(gate403inter7));
  inv1  gate2011(.a(G1084), .O(gate403inter8));
  nand2 gate2012(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2013(.a(s_209), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2014(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2015(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2016(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2241(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2242(.a(gate408inter0), .b(s_242), .O(gate408inter1));
  and2  gate2243(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2244(.a(s_242), .O(gate408inter3));
  inv1  gate2245(.a(s_243), .O(gate408inter4));
  nand2 gate2246(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2247(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2248(.a(G22), .O(gate408inter7));
  inv1  gate2249(.a(G1099), .O(gate408inter8));
  nand2 gate2250(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2251(.a(s_243), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2252(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2253(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2254(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2101(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2102(.a(gate412inter0), .b(s_222), .O(gate412inter1));
  and2  gate2103(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2104(.a(s_222), .O(gate412inter3));
  inv1  gate2105(.a(s_223), .O(gate412inter4));
  nand2 gate2106(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2107(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2108(.a(G26), .O(gate412inter7));
  inv1  gate2109(.a(G1111), .O(gate412inter8));
  nand2 gate2110(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2111(.a(s_223), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2112(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2113(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2114(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1191(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1192(.a(gate415inter0), .b(s_92), .O(gate415inter1));
  and2  gate1193(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1194(.a(s_92), .O(gate415inter3));
  inv1  gate1195(.a(s_93), .O(gate415inter4));
  nand2 gate1196(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1197(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1198(.a(G29), .O(gate415inter7));
  inv1  gate1199(.a(G1120), .O(gate415inter8));
  nand2 gate1200(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1201(.a(s_93), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1202(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1203(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1204(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate855(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate856(.a(gate416inter0), .b(s_44), .O(gate416inter1));
  and2  gate857(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate858(.a(s_44), .O(gate416inter3));
  inv1  gate859(.a(s_45), .O(gate416inter4));
  nand2 gate860(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate861(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate862(.a(G30), .O(gate416inter7));
  inv1  gate863(.a(G1123), .O(gate416inter8));
  nand2 gate864(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate865(.a(s_45), .b(gate416inter3), .O(gate416inter10));
  nor2  gate866(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate867(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate868(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1947(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1948(.a(gate417inter0), .b(s_200), .O(gate417inter1));
  and2  gate1949(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1950(.a(s_200), .O(gate417inter3));
  inv1  gate1951(.a(s_201), .O(gate417inter4));
  nand2 gate1952(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1953(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1954(.a(G31), .O(gate417inter7));
  inv1  gate1955(.a(G1126), .O(gate417inter8));
  nand2 gate1956(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1957(.a(s_201), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1958(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1959(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1960(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1667(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1668(.a(gate419inter0), .b(s_160), .O(gate419inter1));
  and2  gate1669(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1670(.a(s_160), .O(gate419inter3));
  inv1  gate1671(.a(s_161), .O(gate419inter4));
  nand2 gate1672(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1673(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1674(.a(G1), .O(gate419inter7));
  inv1  gate1675(.a(G1132), .O(gate419inter8));
  nand2 gate1676(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1677(.a(s_161), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1678(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1679(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1680(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1233(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1234(.a(gate427inter0), .b(s_98), .O(gate427inter1));
  and2  gate1235(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1236(.a(s_98), .O(gate427inter3));
  inv1  gate1237(.a(s_99), .O(gate427inter4));
  nand2 gate1238(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1239(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1240(.a(G5), .O(gate427inter7));
  inv1  gate1241(.a(G1144), .O(gate427inter8));
  nand2 gate1242(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1243(.a(s_99), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1244(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1245(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1246(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2367(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2368(.a(gate430inter0), .b(s_260), .O(gate430inter1));
  and2  gate2369(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2370(.a(s_260), .O(gate430inter3));
  inv1  gate2371(.a(s_261), .O(gate430inter4));
  nand2 gate2372(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2373(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2374(.a(G1051), .O(gate430inter7));
  inv1  gate2375(.a(G1147), .O(gate430inter8));
  nand2 gate2376(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2377(.a(s_261), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2378(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2379(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2380(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1317(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1318(.a(gate435inter0), .b(s_110), .O(gate435inter1));
  and2  gate1319(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1320(.a(s_110), .O(gate435inter3));
  inv1  gate1321(.a(s_111), .O(gate435inter4));
  nand2 gate1322(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1323(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1324(.a(G9), .O(gate435inter7));
  inv1  gate1325(.a(G1156), .O(gate435inter8));
  nand2 gate1326(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1327(.a(s_111), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1328(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1329(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1330(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate911(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate912(.a(gate437inter0), .b(s_52), .O(gate437inter1));
  and2  gate913(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate914(.a(s_52), .O(gate437inter3));
  inv1  gate915(.a(s_53), .O(gate437inter4));
  nand2 gate916(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate917(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate918(.a(G10), .O(gate437inter7));
  inv1  gate919(.a(G1159), .O(gate437inter8));
  nand2 gate920(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate921(.a(s_53), .b(gate437inter3), .O(gate437inter10));
  nor2  gate922(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate923(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate924(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1653(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1654(.a(gate438inter0), .b(s_158), .O(gate438inter1));
  and2  gate1655(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1656(.a(s_158), .O(gate438inter3));
  inv1  gate1657(.a(s_159), .O(gate438inter4));
  nand2 gate1658(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1659(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1660(.a(G1063), .O(gate438inter7));
  inv1  gate1661(.a(G1159), .O(gate438inter8));
  nand2 gate1662(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1663(.a(s_159), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1664(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1665(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1666(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1163(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1164(.a(gate440inter0), .b(s_88), .O(gate440inter1));
  and2  gate1165(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1166(.a(s_88), .O(gate440inter3));
  inv1  gate1167(.a(s_89), .O(gate440inter4));
  nand2 gate1168(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1169(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1170(.a(G1066), .O(gate440inter7));
  inv1  gate1171(.a(G1162), .O(gate440inter8));
  nand2 gate1172(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1173(.a(s_89), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1174(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1175(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1176(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1527(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1528(.a(gate441inter0), .b(s_140), .O(gate441inter1));
  and2  gate1529(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1530(.a(s_140), .O(gate441inter3));
  inv1  gate1531(.a(s_141), .O(gate441inter4));
  nand2 gate1532(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1533(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1534(.a(G12), .O(gate441inter7));
  inv1  gate1535(.a(G1165), .O(gate441inter8));
  nand2 gate1536(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1537(.a(s_141), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1538(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1539(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1540(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1933(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1934(.a(gate450inter0), .b(s_198), .O(gate450inter1));
  and2  gate1935(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1936(.a(s_198), .O(gate450inter3));
  inv1  gate1937(.a(s_199), .O(gate450inter4));
  nand2 gate1938(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1939(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1940(.a(G1081), .O(gate450inter7));
  inv1  gate1941(.a(G1177), .O(gate450inter8));
  nand2 gate1942(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1943(.a(s_199), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1944(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1945(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1946(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2171(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2172(.a(gate453inter0), .b(s_232), .O(gate453inter1));
  and2  gate2173(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2174(.a(s_232), .O(gate453inter3));
  inv1  gate2175(.a(s_233), .O(gate453inter4));
  nand2 gate2176(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2177(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2178(.a(G18), .O(gate453inter7));
  inv1  gate2179(.a(G1183), .O(gate453inter8));
  nand2 gate2180(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2181(.a(s_233), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2182(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2183(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2184(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate2437(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2438(.a(gate454inter0), .b(s_270), .O(gate454inter1));
  and2  gate2439(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2440(.a(s_270), .O(gate454inter3));
  inv1  gate2441(.a(s_271), .O(gate454inter4));
  nand2 gate2442(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2443(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2444(.a(G1087), .O(gate454inter7));
  inv1  gate2445(.a(G1183), .O(gate454inter8));
  nand2 gate2446(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2447(.a(s_271), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2448(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2449(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2450(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2535(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2536(.a(gate456inter0), .b(s_284), .O(gate456inter1));
  and2  gate2537(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2538(.a(s_284), .O(gate456inter3));
  inv1  gate2539(.a(s_285), .O(gate456inter4));
  nand2 gate2540(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2541(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2542(.a(G1090), .O(gate456inter7));
  inv1  gate2543(.a(G1186), .O(gate456inter8));
  nand2 gate2544(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2545(.a(s_285), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2546(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2547(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2548(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2451(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2452(.a(gate458inter0), .b(s_272), .O(gate458inter1));
  and2  gate2453(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2454(.a(s_272), .O(gate458inter3));
  inv1  gate2455(.a(s_273), .O(gate458inter4));
  nand2 gate2456(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2457(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2458(.a(G1093), .O(gate458inter7));
  inv1  gate2459(.a(G1189), .O(gate458inter8));
  nand2 gate2460(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2461(.a(s_273), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2462(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2463(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2464(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate2647(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2648(.a(gate459inter0), .b(s_300), .O(gate459inter1));
  and2  gate2649(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2650(.a(s_300), .O(gate459inter3));
  inv1  gate2651(.a(s_301), .O(gate459inter4));
  nand2 gate2652(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2653(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2654(.a(G21), .O(gate459inter7));
  inv1  gate2655(.a(G1192), .O(gate459inter8));
  nand2 gate2656(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2657(.a(s_301), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2658(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2659(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2660(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate2185(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2186(.a(gate460inter0), .b(s_234), .O(gate460inter1));
  and2  gate2187(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2188(.a(s_234), .O(gate460inter3));
  inv1  gate2189(.a(s_235), .O(gate460inter4));
  nand2 gate2190(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2191(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2192(.a(G1096), .O(gate460inter7));
  inv1  gate2193(.a(G1192), .O(gate460inter8));
  nand2 gate2194(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2195(.a(s_235), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2196(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2197(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2198(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2269(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2270(.a(gate462inter0), .b(s_246), .O(gate462inter1));
  and2  gate2271(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2272(.a(s_246), .O(gate462inter3));
  inv1  gate2273(.a(s_247), .O(gate462inter4));
  nand2 gate2274(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2275(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2276(.a(G1099), .O(gate462inter7));
  inv1  gate2277(.a(G1195), .O(gate462inter8));
  nand2 gate2278(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2279(.a(s_247), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2280(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2281(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2282(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2759(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2760(.a(gate464inter0), .b(s_316), .O(gate464inter1));
  and2  gate2761(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2762(.a(s_316), .O(gate464inter3));
  inv1  gate2763(.a(s_317), .O(gate464inter4));
  nand2 gate2764(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2765(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2766(.a(G1102), .O(gate464inter7));
  inv1  gate2767(.a(G1198), .O(gate464inter8));
  nand2 gate2768(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2769(.a(s_317), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2770(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2771(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2772(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2087(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2088(.a(gate467inter0), .b(s_220), .O(gate467inter1));
  and2  gate2089(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2090(.a(s_220), .O(gate467inter3));
  inv1  gate2091(.a(s_221), .O(gate467inter4));
  nand2 gate2092(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2093(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2094(.a(G25), .O(gate467inter7));
  inv1  gate2095(.a(G1204), .O(gate467inter8));
  nand2 gate2096(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2097(.a(s_221), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2098(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2099(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2100(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate659(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate660(.a(gate468inter0), .b(s_16), .O(gate468inter1));
  and2  gate661(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate662(.a(s_16), .O(gate468inter3));
  inv1  gate663(.a(s_17), .O(gate468inter4));
  nand2 gate664(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate665(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate666(.a(G1108), .O(gate468inter7));
  inv1  gate667(.a(G1204), .O(gate468inter8));
  nand2 gate668(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate669(.a(s_17), .b(gate468inter3), .O(gate468inter10));
  nor2  gate670(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate671(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate672(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1373(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1374(.a(gate470inter0), .b(s_118), .O(gate470inter1));
  and2  gate1375(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1376(.a(s_118), .O(gate470inter3));
  inv1  gate1377(.a(s_119), .O(gate470inter4));
  nand2 gate1378(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1379(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1380(.a(G1111), .O(gate470inter7));
  inv1  gate1381(.a(G1207), .O(gate470inter8));
  nand2 gate1382(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1383(.a(s_119), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1384(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1385(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1386(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1723(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1724(.a(gate472inter0), .b(s_168), .O(gate472inter1));
  and2  gate1725(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1726(.a(s_168), .O(gate472inter3));
  inv1  gate1727(.a(s_169), .O(gate472inter4));
  nand2 gate1728(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1729(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1730(.a(G1114), .O(gate472inter7));
  inv1  gate1731(.a(G1210), .O(gate472inter8));
  nand2 gate1732(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1733(.a(s_169), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1734(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1735(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1736(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1569(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1570(.a(gate473inter0), .b(s_146), .O(gate473inter1));
  and2  gate1571(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1572(.a(s_146), .O(gate473inter3));
  inv1  gate1573(.a(s_147), .O(gate473inter4));
  nand2 gate1574(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1575(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1576(.a(G28), .O(gate473inter7));
  inv1  gate1577(.a(G1213), .O(gate473inter8));
  nand2 gate1578(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1579(.a(s_147), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1580(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1581(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1582(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1835(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1836(.a(gate477inter0), .b(s_184), .O(gate477inter1));
  and2  gate1837(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1838(.a(s_184), .O(gate477inter3));
  inv1  gate1839(.a(s_185), .O(gate477inter4));
  nand2 gate1840(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1841(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1842(.a(G30), .O(gate477inter7));
  inv1  gate1843(.a(G1219), .O(gate477inter8));
  nand2 gate1844(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1845(.a(s_185), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1846(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1847(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1848(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate2031(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2032(.a(gate478inter0), .b(s_212), .O(gate478inter1));
  and2  gate2033(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2034(.a(s_212), .O(gate478inter3));
  inv1  gate2035(.a(s_213), .O(gate478inter4));
  nand2 gate2036(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2037(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2038(.a(G1123), .O(gate478inter7));
  inv1  gate2039(.a(G1219), .O(gate478inter8));
  nand2 gate2040(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2041(.a(s_213), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2042(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2043(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2044(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1961(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1962(.a(gate486inter0), .b(s_202), .O(gate486inter1));
  and2  gate1963(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1964(.a(s_202), .O(gate486inter3));
  inv1  gate1965(.a(s_203), .O(gate486inter4));
  nand2 gate1966(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1967(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1968(.a(G1234), .O(gate486inter7));
  inv1  gate1969(.a(G1235), .O(gate486inter8));
  nand2 gate1970(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1971(.a(s_203), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1972(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1973(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1974(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1261(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1262(.a(gate487inter0), .b(s_102), .O(gate487inter1));
  and2  gate1263(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1264(.a(s_102), .O(gate487inter3));
  inv1  gate1265(.a(s_103), .O(gate487inter4));
  nand2 gate1266(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1267(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1268(.a(G1236), .O(gate487inter7));
  inv1  gate1269(.a(G1237), .O(gate487inter8));
  nand2 gate1270(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1271(.a(s_103), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1272(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1273(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1274(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1541(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1542(.a(gate489inter0), .b(s_142), .O(gate489inter1));
  and2  gate1543(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1544(.a(s_142), .O(gate489inter3));
  inv1  gate1545(.a(s_143), .O(gate489inter4));
  nand2 gate1546(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1547(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1548(.a(G1240), .O(gate489inter7));
  inv1  gate1549(.a(G1241), .O(gate489inter8));
  nand2 gate1550(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1551(.a(s_143), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1552(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1553(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1554(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2591(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2592(.a(gate493inter0), .b(s_292), .O(gate493inter1));
  and2  gate2593(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2594(.a(s_292), .O(gate493inter3));
  inv1  gate2595(.a(s_293), .O(gate493inter4));
  nand2 gate2596(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2597(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2598(.a(G1248), .O(gate493inter7));
  inv1  gate2599(.a(G1249), .O(gate493inter8));
  nand2 gate2600(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2601(.a(s_293), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2602(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2603(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2604(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1107(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1108(.a(gate494inter0), .b(s_80), .O(gate494inter1));
  and2  gate1109(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1110(.a(s_80), .O(gate494inter3));
  inv1  gate1111(.a(s_81), .O(gate494inter4));
  nand2 gate1112(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1113(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1114(.a(G1250), .O(gate494inter7));
  inv1  gate1115(.a(G1251), .O(gate494inter8));
  nand2 gate1116(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1117(.a(s_81), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1118(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1119(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1120(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate939(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate940(.a(gate497inter0), .b(s_56), .O(gate497inter1));
  and2  gate941(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate942(.a(s_56), .O(gate497inter3));
  inv1  gate943(.a(s_57), .O(gate497inter4));
  nand2 gate944(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate945(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate946(.a(G1256), .O(gate497inter7));
  inv1  gate947(.a(G1257), .O(gate497inter8));
  nand2 gate948(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate949(.a(s_57), .b(gate497inter3), .O(gate497inter10));
  nor2  gate950(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate951(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate952(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate771(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate772(.a(gate498inter0), .b(s_32), .O(gate498inter1));
  and2  gate773(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate774(.a(s_32), .O(gate498inter3));
  inv1  gate775(.a(s_33), .O(gate498inter4));
  nand2 gate776(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate777(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate778(.a(G1258), .O(gate498inter7));
  inv1  gate779(.a(G1259), .O(gate498inter8));
  nand2 gate780(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate781(.a(s_33), .b(gate498inter3), .O(gate498inter10));
  nor2  gate782(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate783(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate784(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1583(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1584(.a(gate502inter0), .b(s_148), .O(gate502inter1));
  and2  gate1585(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1586(.a(s_148), .O(gate502inter3));
  inv1  gate1587(.a(s_149), .O(gate502inter4));
  nand2 gate1588(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1589(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1590(.a(G1266), .O(gate502inter7));
  inv1  gate1591(.a(G1267), .O(gate502inter8));
  nand2 gate1592(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1593(.a(s_149), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1594(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1595(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1596(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1639(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1640(.a(gate505inter0), .b(s_156), .O(gate505inter1));
  and2  gate1641(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1642(.a(s_156), .O(gate505inter3));
  inv1  gate1643(.a(s_157), .O(gate505inter4));
  nand2 gate1644(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1645(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1646(.a(G1272), .O(gate505inter7));
  inv1  gate1647(.a(G1273), .O(gate505inter8));
  nand2 gate1648(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1649(.a(s_157), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1650(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1651(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1652(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1513(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1514(.a(gate506inter0), .b(s_138), .O(gate506inter1));
  and2  gate1515(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1516(.a(s_138), .O(gate506inter3));
  inv1  gate1517(.a(s_139), .O(gate506inter4));
  nand2 gate1518(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1519(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1520(.a(G1274), .O(gate506inter7));
  inv1  gate1521(.a(G1275), .O(gate506inter8));
  nand2 gate1522(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1523(.a(s_139), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1524(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1525(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1526(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate981(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate982(.a(gate511inter0), .b(s_62), .O(gate511inter1));
  and2  gate983(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate984(.a(s_62), .O(gate511inter3));
  inv1  gate985(.a(s_63), .O(gate511inter4));
  nand2 gate986(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate987(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate988(.a(G1284), .O(gate511inter7));
  inv1  gate989(.a(G1285), .O(gate511inter8));
  nand2 gate990(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate991(.a(s_63), .b(gate511inter3), .O(gate511inter10));
  nor2  gate992(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate993(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate994(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2577(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2578(.a(gate514inter0), .b(s_290), .O(gate514inter1));
  and2  gate2579(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2580(.a(s_290), .O(gate514inter3));
  inv1  gate2581(.a(s_291), .O(gate514inter4));
  nand2 gate2582(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2583(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2584(.a(G1290), .O(gate514inter7));
  inv1  gate2585(.a(G1291), .O(gate514inter8));
  nand2 gate2586(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2587(.a(s_291), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2588(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2589(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2590(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule