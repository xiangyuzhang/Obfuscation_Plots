module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1653(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1654(.a(gate16inter0), .b(s_158), .O(gate16inter1));
  and2  gate1655(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1656(.a(s_158), .O(gate16inter3));
  inv1  gate1657(.a(s_159), .O(gate16inter4));
  nand2 gate1658(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1659(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1660(.a(G15), .O(gate16inter7));
  inv1  gate1661(.a(G16), .O(gate16inter8));
  nand2 gate1662(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1663(.a(s_159), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1664(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1665(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1666(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate813(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate814(.a(gate22inter0), .b(s_38), .O(gate22inter1));
  and2  gate815(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate816(.a(s_38), .O(gate22inter3));
  inv1  gate817(.a(s_39), .O(gate22inter4));
  nand2 gate818(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate819(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate820(.a(G27), .O(gate22inter7));
  inv1  gate821(.a(G28), .O(gate22inter8));
  nand2 gate822(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate823(.a(s_39), .b(gate22inter3), .O(gate22inter10));
  nor2  gate824(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate825(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate826(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2143(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2144(.a(gate24inter0), .b(s_228), .O(gate24inter1));
  and2  gate2145(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2146(.a(s_228), .O(gate24inter3));
  inv1  gate2147(.a(s_229), .O(gate24inter4));
  nand2 gate2148(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2149(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2150(.a(G31), .O(gate24inter7));
  inv1  gate2151(.a(G32), .O(gate24inter8));
  nand2 gate2152(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2153(.a(s_229), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2154(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2155(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2156(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate2171(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2172(.a(gate25inter0), .b(s_232), .O(gate25inter1));
  and2  gate2173(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2174(.a(s_232), .O(gate25inter3));
  inv1  gate2175(.a(s_233), .O(gate25inter4));
  nand2 gate2176(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2177(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2178(.a(G1), .O(gate25inter7));
  inv1  gate2179(.a(G5), .O(gate25inter8));
  nand2 gate2180(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2181(.a(s_233), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2182(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2183(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2184(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate939(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate940(.a(gate26inter0), .b(s_56), .O(gate26inter1));
  and2  gate941(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate942(.a(s_56), .O(gate26inter3));
  inv1  gate943(.a(s_57), .O(gate26inter4));
  nand2 gate944(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate945(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate946(.a(G9), .O(gate26inter7));
  inv1  gate947(.a(G13), .O(gate26inter8));
  nand2 gate948(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate949(.a(s_57), .b(gate26inter3), .O(gate26inter10));
  nor2  gate950(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate951(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate952(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate841(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate842(.a(gate28inter0), .b(s_42), .O(gate28inter1));
  and2  gate843(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate844(.a(s_42), .O(gate28inter3));
  inv1  gate845(.a(s_43), .O(gate28inter4));
  nand2 gate846(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate847(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate848(.a(G10), .O(gate28inter7));
  inv1  gate849(.a(G14), .O(gate28inter8));
  nand2 gate850(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate851(.a(s_43), .b(gate28inter3), .O(gate28inter10));
  nor2  gate852(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate853(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate854(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2927(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2928(.a(gate29inter0), .b(s_340), .O(gate29inter1));
  and2  gate2929(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2930(.a(s_340), .O(gate29inter3));
  inv1  gate2931(.a(s_341), .O(gate29inter4));
  nand2 gate2932(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2933(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2934(.a(G3), .O(gate29inter7));
  inv1  gate2935(.a(G7), .O(gate29inter8));
  nand2 gate2936(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2937(.a(s_341), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2938(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2939(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2940(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1009(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1010(.a(gate36inter0), .b(s_66), .O(gate36inter1));
  and2  gate1011(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1012(.a(s_66), .O(gate36inter3));
  inv1  gate1013(.a(s_67), .O(gate36inter4));
  nand2 gate1014(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1015(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1016(.a(G26), .O(gate36inter7));
  inv1  gate1017(.a(G30), .O(gate36inter8));
  nand2 gate1018(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1019(.a(s_67), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1020(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1021(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1022(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate883(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate884(.a(gate37inter0), .b(s_48), .O(gate37inter1));
  and2  gate885(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate886(.a(s_48), .O(gate37inter3));
  inv1  gate887(.a(s_49), .O(gate37inter4));
  nand2 gate888(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate889(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate890(.a(G19), .O(gate37inter7));
  inv1  gate891(.a(G23), .O(gate37inter8));
  nand2 gate892(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate893(.a(s_49), .b(gate37inter3), .O(gate37inter10));
  nor2  gate894(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate895(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate896(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate3179(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate3180(.a(gate41inter0), .b(s_376), .O(gate41inter1));
  and2  gate3181(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate3182(.a(s_376), .O(gate41inter3));
  inv1  gate3183(.a(s_377), .O(gate41inter4));
  nand2 gate3184(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate3185(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate3186(.a(G1), .O(gate41inter7));
  inv1  gate3187(.a(G266), .O(gate41inter8));
  nand2 gate3188(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate3189(.a(s_377), .b(gate41inter3), .O(gate41inter10));
  nor2  gate3190(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate3191(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate3192(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1219(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1220(.a(gate42inter0), .b(s_96), .O(gate42inter1));
  and2  gate1221(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1222(.a(s_96), .O(gate42inter3));
  inv1  gate1223(.a(s_97), .O(gate42inter4));
  nand2 gate1224(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1225(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1226(.a(G2), .O(gate42inter7));
  inv1  gate1227(.a(G266), .O(gate42inter8));
  nand2 gate1228(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1229(.a(s_97), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1230(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1231(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1232(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate2843(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2844(.a(gate43inter0), .b(s_328), .O(gate43inter1));
  and2  gate2845(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2846(.a(s_328), .O(gate43inter3));
  inv1  gate2847(.a(s_329), .O(gate43inter4));
  nand2 gate2848(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2849(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2850(.a(G3), .O(gate43inter7));
  inv1  gate2851(.a(G269), .O(gate43inter8));
  nand2 gate2852(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2853(.a(s_329), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2854(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2855(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2856(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate603(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate604(.a(gate44inter0), .b(s_8), .O(gate44inter1));
  and2  gate605(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate606(.a(s_8), .O(gate44inter3));
  inv1  gate607(.a(s_9), .O(gate44inter4));
  nand2 gate608(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate609(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate610(.a(G4), .O(gate44inter7));
  inv1  gate611(.a(G269), .O(gate44inter8));
  nand2 gate612(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate613(.a(s_9), .b(gate44inter3), .O(gate44inter10));
  nor2  gate614(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate615(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate616(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1037(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1038(.a(gate45inter0), .b(s_70), .O(gate45inter1));
  and2  gate1039(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1040(.a(s_70), .O(gate45inter3));
  inv1  gate1041(.a(s_71), .O(gate45inter4));
  nand2 gate1042(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1043(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1044(.a(G5), .O(gate45inter7));
  inv1  gate1045(.a(G272), .O(gate45inter8));
  nand2 gate1046(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1047(.a(s_71), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1048(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1049(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1050(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2577(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2578(.a(gate49inter0), .b(s_290), .O(gate49inter1));
  and2  gate2579(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2580(.a(s_290), .O(gate49inter3));
  inv1  gate2581(.a(s_291), .O(gate49inter4));
  nand2 gate2582(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2583(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2584(.a(G9), .O(gate49inter7));
  inv1  gate2585(.a(G278), .O(gate49inter8));
  nand2 gate2586(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2587(.a(s_291), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2588(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2589(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2590(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate1905(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1906(.a(gate50inter0), .b(s_194), .O(gate50inter1));
  and2  gate1907(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1908(.a(s_194), .O(gate50inter3));
  inv1  gate1909(.a(s_195), .O(gate50inter4));
  nand2 gate1910(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1911(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1912(.a(G10), .O(gate50inter7));
  inv1  gate1913(.a(G278), .O(gate50inter8));
  nand2 gate1914(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1915(.a(s_195), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1916(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1917(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1918(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate2675(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2676(.a(gate51inter0), .b(s_304), .O(gate51inter1));
  and2  gate2677(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2678(.a(s_304), .O(gate51inter3));
  inv1  gate2679(.a(s_305), .O(gate51inter4));
  nand2 gate2680(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2681(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2682(.a(G11), .O(gate51inter7));
  inv1  gate2683(.a(G281), .O(gate51inter8));
  nand2 gate2684(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2685(.a(s_305), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2686(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2687(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2688(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate3109(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate3110(.a(gate56inter0), .b(s_366), .O(gate56inter1));
  and2  gate3111(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate3112(.a(s_366), .O(gate56inter3));
  inv1  gate3113(.a(s_367), .O(gate56inter4));
  nand2 gate3114(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate3115(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate3116(.a(G16), .O(gate56inter7));
  inv1  gate3117(.a(G287), .O(gate56inter8));
  nand2 gate3118(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate3119(.a(s_367), .b(gate56inter3), .O(gate56inter10));
  nor2  gate3120(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate3121(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate3122(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1751(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1752(.a(gate57inter0), .b(s_172), .O(gate57inter1));
  and2  gate1753(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1754(.a(s_172), .O(gate57inter3));
  inv1  gate1755(.a(s_173), .O(gate57inter4));
  nand2 gate1756(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1757(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1758(.a(G17), .O(gate57inter7));
  inv1  gate1759(.a(G290), .O(gate57inter8));
  nand2 gate1760(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1761(.a(s_173), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1762(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1763(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1764(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate2787(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2788(.a(gate58inter0), .b(s_320), .O(gate58inter1));
  and2  gate2789(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2790(.a(s_320), .O(gate58inter3));
  inv1  gate2791(.a(s_321), .O(gate58inter4));
  nand2 gate2792(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2793(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2794(.a(G18), .O(gate58inter7));
  inv1  gate2795(.a(G290), .O(gate58inter8));
  nand2 gate2796(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2797(.a(s_321), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2798(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2799(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2800(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2003(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2004(.a(gate61inter0), .b(s_208), .O(gate61inter1));
  and2  gate2005(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2006(.a(s_208), .O(gate61inter3));
  inv1  gate2007(.a(s_209), .O(gate61inter4));
  nand2 gate2008(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2009(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2010(.a(G21), .O(gate61inter7));
  inv1  gate2011(.a(G296), .O(gate61inter8));
  nand2 gate2012(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2013(.a(s_209), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2014(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2015(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2016(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1513(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1514(.a(gate64inter0), .b(s_138), .O(gate64inter1));
  and2  gate1515(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1516(.a(s_138), .O(gate64inter3));
  inv1  gate1517(.a(s_139), .O(gate64inter4));
  nand2 gate1518(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1519(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1520(.a(G24), .O(gate64inter7));
  inv1  gate1521(.a(G299), .O(gate64inter8));
  nand2 gate1522(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1523(.a(s_139), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1524(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1525(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1526(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1457(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1458(.a(gate66inter0), .b(s_130), .O(gate66inter1));
  and2  gate1459(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1460(.a(s_130), .O(gate66inter3));
  inv1  gate1461(.a(s_131), .O(gate66inter4));
  nand2 gate1462(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1463(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1464(.a(G26), .O(gate66inter7));
  inv1  gate1465(.a(G302), .O(gate66inter8));
  nand2 gate1466(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1467(.a(s_131), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1468(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1469(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1470(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2479(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2480(.a(gate69inter0), .b(s_276), .O(gate69inter1));
  and2  gate2481(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2482(.a(s_276), .O(gate69inter3));
  inv1  gate2483(.a(s_277), .O(gate69inter4));
  nand2 gate2484(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2485(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2486(.a(G29), .O(gate69inter7));
  inv1  gate2487(.a(G308), .O(gate69inter8));
  nand2 gate2488(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2489(.a(s_277), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2490(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2491(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2492(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2801(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2802(.a(gate72inter0), .b(s_322), .O(gate72inter1));
  and2  gate2803(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2804(.a(s_322), .O(gate72inter3));
  inv1  gate2805(.a(s_323), .O(gate72inter4));
  nand2 gate2806(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2807(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2808(.a(G32), .O(gate72inter7));
  inv1  gate2809(.a(G311), .O(gate72inter8));
  nand2 gate2810(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2811(.a(s_323), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2812(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2813(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2814(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1891(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1892(.a(gate73inter0), .b(s_192), .O(gate73inter1));
  and2  gate1893(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1894(.a(s_192), .O(gate73inter3));
  inv1  gate1895(.a(s_193), .O(gate73inter4));
  nand2 gate1896(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1897(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1898(.a(G1), .O(gate73inter7));
  inv1  gate1899(.a(G314), .O(gate73inter8));
  nand2 gate1900(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1901(.a(s_193), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1902(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1903(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1904(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2661(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2662(.a(gate74inter0), .b(s_302), .O(gate74inter1));
  and2  gate2663(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2664(.a(s_302), .O(gate74inter3));
  inv1  gate2665(.a(s_303), .O(gate74inter4));
  nand2 gate2666(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2667(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2668(.a(G5), .O(gate74inter7));
  inv1  gate2669(.a(G314), .O(gate74inter8));
  nand2 gate2670(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2671(.a(s_303), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2672(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2673(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2674(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1709(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1710(.a(gate80inter0), .b(s_166), .O(gate80inter1));
  and2  gate1711(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1712(.a(s_166), .O(gate80inter3));
  inv1  gate1713(.a(s_167), .O(gate80inter4));
  nand2 gate1714(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1715(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1716(.a(G14), .O(gate80inter7));
  inv1  gate1717(.a(G323), .O(gate80inter8));
  nand2 gate1718(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1719(.a(s_167), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1720(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1721(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1722(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2717(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2718(.a(gate81inter0), .b(s_310), .O(gate81inter1));
  and2  gate2719(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2720(.a(s_310), .O(gate81inter3));
  inv1  gate2721(.a(s_311), .O(gate81inter4));
  nand2 gate2722(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2723(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2724(.a(G3), .O(gate81inter7));
  inv1  gate2725(.a(G326), .O(gate81inter8));
  nand2 gate2726(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2727(.a(s_311), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2728(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2729(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2730(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate3011(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate3012(.a(gate82inter0), .b(s_352), .O(gate82inter1));
  and2  gate3013(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate3014(.a(s_352), .O(gate82inter3));
  inv1  gate3015(.a(s_353), .O(gate82inter4));
  nand2 gate3016(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate3017(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate3018(.a(G7), .O(gate82inter7));
  inv1  gate3019(.a(G326), .O(gate82inter8));
  nand2 gate3020(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate3021(.a(s_353), .b(gate82inter3), .O(gate82inter10));
  nor2  gate3022(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate3023(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate3024(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1541(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1542(.a(gate85inter0), .b(s_142), .O(gate85inter1));
  and2  gate1543(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1544(.a(s_142), .O(gate85inter3));
  inv1  gate1545(.a(s_143), .O(gate85inter4));
  nand2 gate1546(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1547(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1548(.a(G4), .O(gate85inter7));
  inv1  gate1549(.a(G332), .O(gate85inter8));
  nand2 gate1550(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1551(.a(s_143), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1552(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1553(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1554(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2969(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2970(.a(gate88inter0), .b(s_346), .O(gate88inter1));
  and2  gate2971(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2972(.a(s_346), .O(gate88inter3));
  inv1  gate2973(.a(s_347), .O(gate88inter4));
  nand2 gate2974(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2975(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2976(.a(G16), .O(gate88inter7));
  inv1  gate2977(.a(G335), .O(gate88inter8));
  nand2 gate2978(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2979(.a(s_347), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2980(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2981(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2982(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1863(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1864(.a(gate89inter0), .b(s_188), .O(gate89inter1));
  and2  gate1865(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1866(.a(s_188), .O(gate89inter3));
  inv1  gate1867(.a(s_189), .O(gate89inter4));
  nand2 gate1868(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1869(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1870(.a(G17), .O(gate89inter7));
  inv1  gate1871(.a(G338), .O(gate89inter8));
  nand2 gate1872(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1873(.a(s_189), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1874(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1875(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1876(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate3151(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate3152(.a(gate91inter0), .b(s_372), .O(gate91inter1));
  and2  gate3153(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate3154(.a(s_372), .O(gate91inter3));
  inv1  gate3155(.a(s_373), .O(gate91inter4));
  nand2 gate3156(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate3157(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate3158(.a(G25), .O(gate91inter7));
  inv1  gate3159(.a(G341), .O(gate91inter8));
  nand2 gate3160(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate3161(.a(s_373), .b(gate91inter3), .O(gate91inter10));
  nor2  gate3162(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate3163(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate3164(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate729(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate730(.a(gate93inter0), .b(s_26), .O(gate93inter1));
  and2  gate731(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate732(.a(s_26), .O(gate93inter3));
  inv1  gate733(.a(s_27), .O(gate93inter4));
  nand2 gate734(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate735(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate736(.a(G18), .O(gate93inter7));
  inv1  gate737(.a(G344), .O(gate93inter8));
  nand2 gate738(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate739(.a(s_27), .b(gate93inter3), .O(gate93inter10));
  nor2  gate740(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate741(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate742(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate575(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate576(.a(gate94inter0), .b(s_4), .O(gate94inter1));
  and2  gate577(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate578(.a(s_4), .O(gate94inter3));
  inv1  gate579(.a(s_5), .O(gate94inter4));
  nand2 gate580(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate581(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate582(.a(G22), .O(gate94inter7));
  inv1  gate583(.a(G344), .O(gate94inter8));
  nand2 gate584(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate585(.a(s_5), .b(gate94inter3), .O(gate94inter10));
  nor2  gate586(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate587(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate588(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1471(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1472(.a(gate100inter0), .b(s_132), .O(gate100inter1));
  and2  gate1473(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1474(.a(s_132), .O(gate100inter3));
  inv1  gate1475(.a(s_133), .O(gate100inter4));
  nand2 gate1476(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1477(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1478(.a(G31), .O(gate100inter7));
  inv1  gate1479(.a(G353), .O(gate100inter8));
  nand2 gate1480(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1481(.a(s_133), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1482(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1483(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1484(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate911(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate912(.a(gate101inter0), .b(s_52), .O(gate101inter1));
  and2  gate913(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate914(.a(s_52), .O(gate101inter3));
  inv1  gate915(.a(s_53), .O(gate101inter4));
  nand2 gate916(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate917(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate918(.a(G20), .O(gate101inter7));
  inv1  gate919(.a(G356), .O(gate101inter8));
  nand2 gate920(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate921(.a(s_53), .b(gate101inter3), .O(gate101inter10));
  nor2  gate922(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate923(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate924(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate869(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate870(.a(gate102inter0), .b(s_46), .O(gate102inter1));
  and2  gate871(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate872(.a(s_46), .O(gate102inter3));
  inv1  gate873(.a(s_47), .O(gate102inter4));
  nand2 gate874(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate875(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate876(.a(G24), .O(gate102inter7));
  inv1  gate877(.a(G356), .O(gate102inter8));
  nand2 gate878(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate879(.a(s_47), .b(gate102inter3), .O(gate102inter10));
  nor2  gate880(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate881(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate882(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1485(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1486(.a(gate103inter0), .b(s_134), .O(gate103inter1));
  and2  gate1487(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1488(.a(s_134), .O(gate103inter3));
  inv1  gate1489(.a(s_135), .O(gate103inter4));
  nand2 gate1490(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1491(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1492(.a(G28), .O(gate103inter7));
  inv1  gate1493(.a(G359), .O(gate103inter8));
  nand2 gate1494(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1495(.a(s_135), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1496(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1497(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1498(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1233(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1234(.a(gate107inter0), .b(s_98), .O(gate107inter1));
  and2  gate1235(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1236(.a(s_98), .O(gate107inter3));
  inv1  gate1237(.a(s_99), .O(gate107inter4));
  nand2 gate1238(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1239(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1240(.a(G366), .O(gate107inter7));
  inv1  gate1241(.a(G367), .O(gate107inter8));
  nand2 gate1242(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1243(.a(s_99), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1244(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1245(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1246(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2241(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2242(.a(gate111inter0), .b(s_242), .O(gate111inter1));
  and2  gate2243(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2244(.a(s_242), .O(gate111inter3));
  inv1  gate2245(.a(s_243), .O(gate111inter4));
  nand2 gate2246(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2247(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2248(.a(G374), .O(gate111inter7));
  inv1  gate2249(.a(G375), .O(gate111inter8));
  nand2 gate2250(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2251(.a(s_243), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2252(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2253(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2254(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1807(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1808(.a(gate112inter0), .b(s_180), .O(gate112inter1));
  and2  gate1809(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1810(.a(s_180), .O(gate112inter3));
  inv1  gate1811(.a(s_181), .O(gate112inter4));
  nand2 gate1812(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1813(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1814(.a(G376), .O(gate112inter7));
  inv1  gate1815(.a(G377), .O(gate112inter8));
  nand2 gate1816(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1817(.a(s_181), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1818(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1819(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1820(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1387(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1388(.a(gate114inter0), .b(s_120), .O(gate114inter1));
  and2  gate1389(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1390(.a(s_120), .O(gate114inter3));
  inv1  gate1391(.a(s_121), .O(gate114inter4));
  nand2 gate1392(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1393(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1394(.a(G380), .O(gate114inter7));
  inv1  gate1395(.a(G381), .O(gate114inter8));
  nand2 gate1396(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1397(.a(s_121), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1398(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1399(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1400(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2549(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2550(.a(gate120inter0), .b(s_286), .O(gate120inter1));
  and2  gate2551(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2552(.a(s_286), .O(gate120inter3));
  inv1  gate2553(.a(s_287), .O(gate120inter4));
  nand2 gate2554(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2555(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2556(.a(G392), .O(gate120inter7));
  inv1  gate2557(.a(G393), .O(gate120inter8));
  nand2 gate2558(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2559(.a(s_287), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2560(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2561(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2562(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1919(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1920(.a(gate123inter0), .b(s_196), .O(gate123inter1));
  and2  gate1921(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1922(.a(s_196), .O(gate123inter3));
  inv1  gate1923(.a(s_197), .O(gate123inter4));
  nand2 gate1924(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1925(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1926(.a(G398), .O(gate123inter7));
  inv1  gate1927(.a(G399), .O(gate123inter8));
  nand2 gate1928(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1929(.a(s_197), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1930(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1931(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1932(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1275(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1276(.a(gate125inter0), .b(s_104), .O(gate125inter1));
  and2  gate1277(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1278(.a(s_104), .O(gate125inter3));
  inv1  gate1279(.a(s_105), .O(gate125inter4));
  nand2 gate1280(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1281(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1282(.a(G402), .O(gate125inter7));
  inv1  gate1283(.a(G403), .O(gate125inter8));
  nand2 gate1284(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1285(.a(s_105), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1286(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1287(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1288(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1793(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1794(.a(gate130inter0), .b(s_178), .O(gate130inter1));
  and2  gate1795(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1796(.a(s_178), .O(gate130inter3));
  inv1  gate1797(.a(s_179), .O(gate130inter4));
  nand2 gate1798(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1799(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1800(.a(G412), .O(gate130inter7));
  inv1  gate1801(.a(G413), .O(gate130inter8));
  nand2 gate1802(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1803(.a(s_179), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1804(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1805(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1806(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1191(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1192(.a(gate133inter0), .b(s_92), .O(gate133inter1));
  and2  gate1193(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1194(.a(s_92), .O(gate133inter3));
  inv1  gate1195(.a(s_93), .O(gate133inter4));
  nand2 gate1196(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1197(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1198(.a(G418), .O(gate133inter7));
  inv1  gate1199(.a(G419), .O(gate133inter8));
  nand2 gate1200(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1201(.a(s_93), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1202(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1203(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1204(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1247(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1248(.a(gate134inter0), .b(s_100), .O(gate134inter1));
  and2  gate1249(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1250(.a(s_100), .O(gate134inter3));
  inv1  gate1251(.a(s_101), .O(gate134inter4));
  nand2 gate1252(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1253(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1254(.a(G420), .O(gate134inter7));
  inv1  gate1255(.a(G421), .O(gate134inter8));
  nand2 gate1256(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1257(.a(s_101), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1258(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1259(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1260(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2297(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2298(.a(gate135inter0), .b(s_250), .O(gate135inter1));
  and2  gate2299(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2300(.a(s_250), .O(gate135inter3));
  inv1  gate2301(.a(s_251), .O(gate135inter4));
  nand2 gate2302(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2303(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2304(.a(G422), .O(gate135inter7));
  inv1  gate2305(.a(G423), .O(gate135inter8));
  nand2 gate2306(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2307(.a(s_251), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2308(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2309(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2310(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1289(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1290(.a(gate138inter0), .b(s_106), .O(gate138inter1));
  and2  gate1291(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1292(.a(s_106), .O(gate138inter3));
  inv1  gate1293(.a(s_107), .O(gate138inter4));
  nand2 gate1294(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1295(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1296(.a(G432), .O(gate138inter7));
  inv1  gate1297(.a(G435), .O(gate138inter8));
  nand2 gate1298(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1299(.a(s_107), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1300(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1301(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1302(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1079(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1080(.a(gate139inter0), .b(s_76), .O(gate139inter1));
  and2  gate1081(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1082(.a(s_76), .O(gate139inter3));
  inv1  gate1083(.a(s_77), .O(gate139inter4));
  nand2 gate1084(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1085(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1086(.a(G438), .O(gate139inter7));
  inv1  gate1087(.a(G441), .O(gate139inter8));
  nand2 gate1088(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1089(.a(s_77), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1090(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1091(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1092(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2227(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2228(.a(gate140inter0), .b(s_240), .O(gate140inter1));
  and2  gate2229(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2230(.a(s_240), .O(gate140inter3));
  inv1  gate2231(.a(s_241), .O(gate140inter4));
  nand2 gate2232(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2233(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2234(.a(G444), .O(gate140inter7));
  inv1  gate2235(.a(G447), .O(gate140inter8));
  nand2 gate2236(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2237(.a(s_241), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2238(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2239(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2240(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate855(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate856(.a(gate143inter0), .b(s_44), .O(gate143inter1));
  and2  gate857(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate858(.a(s_44), .O(gate143inter3));
  inv1  gate859(.a(s_45), .O(gate143inter4));
  nand2 gate860(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate861(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate862(.a(G462), .O(gate143inter7));
  inv1  gate863(.a(G465), .O(gate143inter8));
  nand2 gate864(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate865(.a(s_45), .b(gate143inter3), .O(gate143inter10));
  nor2  gate866(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate867(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate868(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate3207(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate3208(.a(gate144inter0), .b(s_380), .O(gate144inter1));
  and2  gate3209(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate3210(.a(s_380), .O(gate144inter3));
  inv1  gate3211(.a(s_381), .O(gate144inter4));
  nand2 gate3212(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate3213(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate3214(.a(G468), .O(gate144inter7));
  inv1  gate3215(.a(G471), .O(gate144inter8));
  nand2 gate3216(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate3217(.a(s_381), .b(gate144inter3), .O(gate144inter10));
  nor2  gate3218(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate3219(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate3220(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate3053(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate3054(.a(gate145inter0), .b(s_358), .O(gate145inter1));
  and2  gate3055(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate3056(.a(s_358), .O(gate145inter3));
  inv1  gate3057(.a(s_359), .O(gate145inter4));
  nand2 gate3058(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate3059(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate3060(.a(G474), .O(gate145inter7));
  inv1  gate3061(.a(G477), .O(gate145inter8));
  nand2 gate3062(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate3063(.a(s_359), .b(gate145inter3), .O(gate145inter10));
  nor2  gate3064(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate3065(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate3066(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate3067(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate3068(.a(gate147inter0), .b(s_360), .O(gate147inter1));
  and2  gate3069(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate3070(.a(s_360), .O(gate147inter3));
  inv1  gate3071(.a(s_361), .O(gate147inter4));
  nand2 gate3072(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate3073(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate3074(.a(G486), .O(gate147inter7));
  inv1  gate3075(.a(G489), .O(gate147inter8));
  nand2 gate3076(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate3077(.a(s_361), .b(gate147inter3), .O(gate147inter10));
  nor2  gate3078(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate3079(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate3080(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2759(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2760(.a(gate149inter0), .b(s_316), .O(gate149inter1));
  and2  gate2761(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2762(.a(s_316), .O(gate149inter3));
  inv1  gate2763(.a(s_317), .O(gate149inter4));
  nand2 gate2764(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2765(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2766(.a(G498), .O(gate149inter7));
  inv1  gate2767(.a(G501), .O(gate149inter8));
  nand2 gate2768(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2769(.a(s_317), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2770(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2771(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2772(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2101(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2102(.a(gate150inter0), .b(s_222), .O(gate150inter1));
  and2  gate2103(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2104(.a(s_222), .O(gate150inter3));
  inv1  gate2105(.a(s_223), .O(gate150inter4));
  nand2 gate2106(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2107(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2108(.a(G504), .O(gate150inter7));
  inv1  gate2109(.a(G507), .O(gate150inter8));
  nand2 gate2110(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2111(.a(s_223), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2112(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2113(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2114(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1583(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1584(.a(gate152inter0), .b(s_148), .O(gate152inter1));
  and2  gate1585(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1586(.a(s_148), .O(gate152inter3));
  inv1  gate1587(.a(s_149), .O(gate152inter4));
  nand2 gate1588(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1589(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1590(.a(G516), .O(gate152inter7));
  inv1  gate1591(.a(G519), .O(gate152inter8));
  nand2 gate1592(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1593(.a(s_149), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1594(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1595(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1596(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2535(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2536(.a(gate157inter0), .b(s_284), .O(gate157inter1));
  and2  gate2537(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2538(.a(s_284), .O(gate157inter3));
  inv1  gate2539(.a(s_285), .O(gate157inter4));
  nand2 gate2540(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2541(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2542(.a(G438), .O(gate157inter7));
  inv1  gate2543(.a(G528), .O(gate157inter8));
  nand2 gate2544(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2545(.a(s_285), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2546(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2547(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2548(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2339(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2340(.a(gate161inter0), .b(s_256), .O(gate161inter1));
  and2  gate2341(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2342(.a(s_256), .O(gate161inter3));
  inv1  gate2343(.a(s_257), .O(gate161inter4));
  nand2 gate2344(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2345(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2346(.a(G450), .O(gate161inter7));
  inv1  gate2347(.a(G534), .O(gate161inter8));
  nand2 gate2348(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2349(.a(s_257), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2350(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2351(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2352(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate2073(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2074(.a(gate162inter0), .b(s_218), .O(gate162inter1));
  and2  gate2075(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2076(.a(s_218), .O(gate162inter3));
  inv1  gate2077(.a(s_219), .O(gate162inter4));
  nand2 gate2078(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2079(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2080(.a(G453), .O(gate162inter7));
  inv1  gate2081(.a(G534), .O(gate162inter8));
  nand2 gate2082(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2083(.a(s_219), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2084(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2085(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2086(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1821(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1822(.a(gate164inter0), .b(s_182), .O(gate164inter1));
  and2  gate1823(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1824(.a(s_182), .O(gate164inter3));
  inv1  gate1825(.a(s_183), .O(gate164inter4));
  nand2 gate1826(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1827(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1828(.a(G459), .O(gate164inter7));
  inv1  gate1829(.a(G537), .O(gate164inter8));
  nand2 gate1830(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1831(.a(s_183), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1832(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1833(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1834(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate925(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate926(.a(gate165inter0), .b(s_54), .O(gate165inter1));
  and2  gate927(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate928(.a(s_54), .O(gate165inter3));
  inv1  gate929(.a(s_55), .O(gate165inter4));
  nand2 gate930(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate931(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate932(.a(G462), .O(gate165inter7));
  inv1  gate933(.a(G540), .O(gate165inter8));
  nand2 gate934(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate935(.a(s_55), .b(gate165inter3), .O(gate165inter10));
  nor2  gate936(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate937(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate938(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate2885(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2886(.a(gate167inter0), .b(s_334), .O(gate167inter1));
  and2  gate2887(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2888(.a(s_334), .O(gate167inter3));
  inv1  gate2889(.a(s_335), .O(gate167inter4));
  nand2 gate2890(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2891(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2892(.a(G468), .O(gate167inter7));
  inv1  gate2893(.a(G543), .O(gate167inter8));
  nand2 gate2894(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2895(.a(s_335), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2896(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2897(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2898(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate659(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate660(.a(gate168inter0), .b(s_16), .O(gate168inter1));
  and2  gate661(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate662(.a(s_16), .O(gate168inter3));
  inv1  gate663(.a(s_17), .O(gate168inter4));
  nand2 gate664(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate665(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate666(.a(G471), .O(gate168inter7));
  inv1  gate667(.a(G543), .O(gate168inter8));
  nand2 gate668(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate669(.a(s_17), .b(gate168inter3), .O(gate168inter10));
  nor2  gate670(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate671(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate672(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2507(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2508(.a(gate169inter0), .b(s_280), .O(gate169inter1));
  and2  gate2509(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2510(.a(s_280), .O(gate169inter3));
  inv1  gate2511(.a(s_281), .O(gate169inter4));
  nand2 gate2512(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2513(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2514(.a(G474), .O(gate169inter7));
  inv1  gate2515(.a(G546), .O(gate169inter8));
  nand2 gate2516(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2517(.a(s_281), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2518(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2519(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2520(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2773(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2774(.a(gate172inter0), .b(s_318), .O(gate172inter1));
  and2  gate2775(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2776(.a(s_318), .O(gate172inter3));
  inv1  gate2777(.a(s_319), .O(gate172inter4));
  nand2 gate2778(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2779(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2780(.a(G483), .O(gate172inter7));
  inv1  gate2781(.a(G549), .O(gate172inter8));
  nand2 gate2782(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2783(.a(s_319), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2784(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2785(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2786(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1639(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1640(.a(gate173inter0), .b(s_156), .O(gate173inter1));
  and2  gate1641(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1642(.a(s_156), .O(gate173inter3));
  inv1  gate1643(.a(s_157), .O(gate173inter4));
  nand2 gate1644(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1645(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1646(.a(G486), .O(gate173inter7));
  inv1  gate1647(.a(G552), .O(gate173inter8));
  nand2 gate1648(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1649(.a(s_157), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1650(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1651(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1652(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2353(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2354(.a(gate179inter0), .b(s_258), .O(gate179inter1));
  and2  gate2355(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2356(.a(s_258), .O(gate179inter3));
  inv1  gate2357(.a(s_259), .O(gate179inter4));
  nand2 gate2358(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2359(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2360(.a(G504), .O(gate179inter7));
  inv1  gate2361(.a(G561), .O(gate179inter8));
  nand2 gate2362(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2363(.a(s_259), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2364(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2365(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2366(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate2199(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2200(.a(gate180inter0), .b(s_236), .O(gate180inter1));
  and2  gate2201(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2202(.a(s_236), .O(gate180inter3));
  inv1  gate2203(.a(s_237), .O(gate180inter4));
  nand2 gate2204(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2205(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2206(.a(G507), .O(gate180inter7));
  inv1  gate2207(.a(G561), .O(gate180inter8));
  nand2 gate2208(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2209(.a(s_237), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2210(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2211(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2212(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2619(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2620(.a(gate182inter0), .b(s_296), .O(gate182inter1));
  and2  gate2621(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2622(.a(s_296), .O(gate182inter3));
  inv1  gate2623(.a(s_297), .O(gate182inter4));
  nand2 gate2624(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2625(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2626(.a(G513), .O(gate182inter7));
  inv1  gate2627(.a(G564), .O(gate182inter8));
  nand2 gate2628(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2629(.a(s_297), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2630(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2631(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2632(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1877(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1878(.a(gate183inter0), .b(s_190), .O(gate183inter1));
  and2  gate1879(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1880(.a(s_190), .O(gate183inter3));
  inv1  gate1881(.a(s_191), .O(gate183inter4));
  nand2 gate1882(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1883(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1884(.a(G516), .O(gate183inter7));
  inv1  gate1885(.a(G567), .O(gate183inter8));
  nand2 gate1886(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1887(.a(s_191), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1888(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1889(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1890(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate3193(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate3194(.a(gate184inter0), .b(s_378), .O(gate184inter1));
  and2  gate3195(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate3196(.a(s_378), .O(gate184inter3));
  inv1  gate3197(.a(s_379), .O(gate184inter4));
  nand2 gate3198(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate3199(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate3200(.a(G519), .O(gate184inter7));
  inv1  gate3201(.a(G567), .O(gate184inter8));
  nand2 gate3202(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate3203(.a(s_379), .b(gate184inter3), .O(gate184inter10));
  nor2  gate3204(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate3205(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate3206(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate827(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate828(.a(gate187inter0), .b(s_40), .O(gate187inter1));
  and2  gate829(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate830(.a(s_40), .O(gate187inter3));
  inv1  gate831(.a(s_41), .O(gate187inter4));
  nand2 gate832(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate833(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate834(.a(G574), .O(gate187inter7));
  inv1  gate835(.a(G575), .O(gate187inter8));
  nand2 gate836(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate837(.a(s_41), .b(gate187inter3), .O(gate187inter10));
  nor2  gate838(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate839(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate840(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate701(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate702(.a(gate190inter0), .b(s_22), .O(gate190inter1));
  and2  gate703(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate704(.a(s_22), .O(gate190inter3));
  inv1  gate705(.a(s_23), .O(gate190inter4));
  nand2 gate706(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate707(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate708(.a(G580), .O(gate190inter7));
  inv1  gate709(.a(G581), .O(gate190inter8));
  nand2 gate710(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate711(.a(s_23), .b(gate190inter3), .O(gate190inter10));
  nor2  gate712(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate713(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate714(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2647(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2648(.a(gate195inter0), .b(s_300), .O(gate195inter1));
  and2  gate2649(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2650(.a(s_300), .O(gate195inter3));
  inv1  gate2651(.a(s_301), .O(gate195inter4));
  nand2 gate2652(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2653(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2654(.a(G590), .O(gate195inter7));
  inv1  gate2655(.a(G591), .O(gate195inter8));
  nand2 gate2656(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2657(.a(s_301), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2658(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2659(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2660(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate3165(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate3166(.a(gate197inter0), .b(s_374), .O(gate197inter1));
  and2  gate3167(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate3168(.a(s_374), .O(gate197inter3));
  inv1  gate3169(.a(s_375), .O(gate197inter4));
  nand2 gate3170(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate3171(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate3172(.a(G594), .O(gate197inter7));
  inv1  gate3173(.a(G595), .O(gate197inter8));
  nand2 gate3174(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate3175(.a(s_375), .b(gate197inter3), .O(gate197inter10));
  nor2  gate3176(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate3177(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate3178(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2689(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2690(.a(gate201inter0), .b(s_306), .O(gate201inter1));
  and2  gate2691(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2692(.a(s_306), .O(gate201inter3));
  inv1  gate2693(.a(s_307), .O(gate201inter4));
  nand2 gate2694(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2695(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2696(.a(G602), .O(gate201inter7));
  inv1  gate2697(.a(G607), .O(gate201inter8));
  nand2 gate2698(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2699(.a(s_307), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2700(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2701(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2702(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2367(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2368(.a(gate205inter0), .b(s_260), .O(gate205inter1));
  and2  gate2369(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2370(.a(s_260), .O(gate205inter3));
  inv1  gate2371(.a(s_261), .O(gate205inter4));
  nand2 gate2372(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2373(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2374(.a(G622), .O(gate205inter7));
  inv1  gate2375(.a(G627), .O(gate205inter8));
  nand2 gate2376(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2377(.a(s_261), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2378(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2379(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2380(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1835(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1836(.a(gate206inter0), .b(s_184), .O(gate206inter1));
  and2  gate1837(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1838(.a(s_184), .O(gate206inter3));
  inv1  gate1839(.a(s_185), .O(gate206inter4));
  nand2 gate1840(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1841(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1842(.a(G632), .O(gate206inter7));
  inv1  gate1843(.a(G637), .O(gate206inter8));
  nand2 gate1844(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1845(.a(s_185), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1846(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1847(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1848(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1947(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1948(.a(gate208inter0), .b(s_200), .O(gate208inter1));
  and2  gate1949(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1950(.a(s_200), .O(gate208inter3));
  inv1  gate1951(.a(s_201), .O(gate208inter4));
  nand2 gate1952(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1953(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1954(.a(G627), .O(gate208inter7));
  inv1  gate1955(.a(G637), .O(gate208inter8));
  nand2 gate1956(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1957(.a(s_201), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1958(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1959(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1960(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1065(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1066(.a(gate209inter0), .b(s_74), .O(gate209inter1));
  and2  gate1067(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1068(.a(s_74), .O(gate209inter3));
  inv1  gate1069(.a(s_75), .O(gate209inter4));
  nand2 gate1070(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1071(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1072(.a(G602), .O(gate209inter7));
  inv1  gate1073(.a(G666), .O(gate209inter8));
  nand2 gate1074(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1075(.a(s_75), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1076(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1077(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1078(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1121(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1122(.a(gate210inter0), .b(s_82), .O(gate210inter1));
  and2  gate1123(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1124(.a(s_82), .O(gate210inter3));
  inv1  gate1125(.a(s_83), .O(gate210inter4));
  nand2 gate1126(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1127(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1128(.a(G607), .O(gate210inter7));
  inv1  gate1129(.a(G666), .O(gate210inter8));
  nand2 gate1130(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1131(.a(s_83), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1132(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1133(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1134(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1555(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1556(.a(gate211inter0), .b(s_144), .O(gate211inter1));
  and2  gate1557(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1558(.a(s_144), .O(gate211inter3));
  inv1  gate1559(.a(s_145), .O(gate211inter4));
  nand2 gate1560(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1561(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1562(.a(G612), .O(gate211inter7));
  inv1  gate1563(.a(G669), .O(gate211inter8));
  nand2 gate1564(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1565(.a(s_145), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1566(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1567(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1568(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2395(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2396(.a(gate214inter0), .b(s_264), .O(gate214inter1));
  and2  gate2397(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2398(.a(s_264), .O(gate214inter3));
  inv1  gate2399(.a(s_265), .O(gate214inter4));
  nand2 gate2400(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2401(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2402(.a(G612), .O(gate214inter7));
  inv1  gate2403(.a(G672), .O(gate214inter8));
  nand2 gate2404(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2405(.a(s_265), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2406(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2407(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2408(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2997(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2998(.a(gate217inter0), .b(s_350), .O(gate217inter1));
  and2  gate2999(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate3000(.a(s_350), .O(gate217inter3));
  inv1  gate3001(.a(s_351), .O(gate217inter4));
  nand2 gate3002(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate3003(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate3004(.a(G622), .O(gate217inter7));
  inv1  gate3005(.a(G678), .O(gate217inter8));
  nand2 gate3006(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate3007(.a(s_351), .b(gate217inter3), .O(gate217inter10));
  nor2  gate3008(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate3009(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate3010(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate3025(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate3026(.a(gate218inter0), .b(s_354), .O(gate218inter1));
  and2  gate3027(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate3028(.a(s_354), .O(gate218inter3));
  inv1  gate3029(.a(s_355), .O(gate218inter4));
  nand2 gate3030(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate3031(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate3032(.a(G627), .O(gate218inter7));
  inv1  gate3033(.a(G678), .O(gate218inter8));
  nand2 gate3034(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate3035(.a(s_355), .b(gate218inter3), .O(gate218inter10));
  nor2  gate3036(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate3037(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate3038(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2731(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2732(.a(gate219inter0), .b(s_312), .O(gate219inter1));
  and2  gate2733(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2734(.a(s_312), .O(gate219inter3));
  inv1  gate2735(.a(s_313), .O(gate219inter4));
  nand2 gate2736(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2737(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2738(.a(G632), .O(gate219inter7));
  inv1  gate2739(.a(G681), .O(gate219inter8));
  nand2 gate2740(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2741(.a(s_313), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2742(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2743(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2744(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate2465(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2466(.a(gate220inter0), .b(s_274), .O(gate220inter1));
  and2  gate2467(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2468(.a(s_274), .O(gate220inter3));
  inv1  gate2469(.a(s_275), .O(gate220inter4));
  nand2 gate2470(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2471(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2472(.a(G637), .O(gate220inter7));
  inv1  gate2473(.a(G681), .O(gate220inter8));
  nand2 gate2474(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2475(.a(s_275), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2476(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2477(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2478(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate3081(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate3082(.a(gate222inter0), .b(s_362), .O(gate222inter1));
  and2  gate3083(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate3084(.a(s_362), .O(gate222inter3));
  inv1  gate3085(.a(s_363), .O(gate222inter4));
  nand2 gate3086(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate3087(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate3088(.a(G632), .O(gate222inter7));
  inv1  gate3089(.a(G684), .O(gate222inter8));
  nand2 gate3090(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate3091(.a(s_363), .b(gate222inter3), .O(gate222inter10));
  nor2  gate3092(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate3093(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate3094(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2409(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2410(.a(gate223inter0), .b(s_266), .O(gate223inter1));
  and2  gate2411(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2412(.a(s_266), .O(gate223inter3));
  inv1  gate2413(.a(s_267), .O(gate223inter4));
  nand2 gate2414(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2415(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2416(.a(G627), .O(gate223inter7));
  inv1  gate2417(.a(G687), .O(gate223inter8));
  nand2 gate2418(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2419(.a(s_267), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2420(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2421(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2422(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1401(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1402(.a(gate226inter0), .b(s_122), .O(gate226inter1));
  and2  gate1403(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1404(.a(s_122), .O(gate226inter3));
  inv1  gate1405(.a(s_123), .O(gate226inter4));
  nand2 gate1406(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1407(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1408(.a(G692), .O(gate226inter7));
  inv1  gate1409(.a(G693), .O(gate226inter8));
  nand2 gate1410(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1411(.a(s_123), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1412(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1413(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1414(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate645(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate646(.a(gate227inter0), .b(s_14), .O(gate227inter1));
  and2  gate647(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate648(.a(s_14), .O(gate227inter3));
  inv1  gate649(.a(s_15), .O(gate227inter4));
  nand2 gate650(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate651(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate652(.a(G694), .O(gate227inter7));
  inv1  gate653(.a(G695), .O(gate227inter8));
  nand2 gate654(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate655(.a(s_15), .b(gate227inter3), .O(gate227inter10));
  nor2  gate656(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate657(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate658(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1499(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1500(.a(gate234inter0), .b(s_136), .O(gate234inter1));
  and2  gate1501(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1502(.a(s_136), .O(gate234inter3));
  inv1  gate1503(.a(s_137), .O(gate234inter4));
  nand2 gate1504(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1505(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1506(.a(G245), .O(gate234inter7));
  inv1  gate1507(.a(G721), .O(gate234inter8));
  nand2 gate1508(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1509(.a(s_137), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1510(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1511(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1512(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2045(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2046(.a(gate236inter0), .b(s_214), .O(gate236inter1));
  and2  gate2047(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2048(.a(s_214), .O(gate236inter3));
  inv1  gate2049(.a(s_215), .O(gate236inter4));
  nand2 gate2050(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2051(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2052(.a(G251), .O(gate236inter7));
  inv1  gate2053(.a(G727), .O(gate236inter8));
  nand2 gate2054(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2055(.a(s_215), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2056(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2057(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2058(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate2087(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2088(.a(gate237inter0), .b(s_220), .O(gate237inter1));
  and2  gate2089(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2090(.a(s_220), .O(gate237inter3));
  inv1  gate2091(.a(s_221), .O(gate237inter4));
  nand2 gate2092(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2093(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2094(.a(G254), .O(gate237inter7));
  inv1  gate2095(.a(G706), .O(gate237inter8));
  nand2 gate2096(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2097(.a(s_221), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2098(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2099(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2100(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate673(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate674(.a(gate240inter0), .b(s_18), .O(gate240inter1));
  and2  gate675(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate676(.a(s_18), .O(gate240inter3));
  inv1  gate677(.a(s_19), .O(gate240inter4));
  nand2 gate678(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate679(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate680(.a(G263), .O(gate240inter7));
  inv1  gate681(.a(G715), .O(gate240inter8));
  nand2 gate682(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate683(.a(s_19), .b(gate240inter3), .O(gate240inter10));
  nor2  gate684(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate685(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate686(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1849(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1850(.a(gate241inter0), .b(s_186), .O(gate241inter1));
  and2  gate1851(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1852(.a(s_186), .O(gate241inter3));
  inv1  gate1853(.a(s_187), .O(gate241inter4));
  nand2 gate1854(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1855(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1856(.a(G242), .O(gate241inter7));
  inv1  gate1857(.a(G730), .O(gate241inter8));
  nand2 gate1858(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1859(.a(s_187), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1860(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1861(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1862(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate771(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate772(.a(gate242inter0), .b(s_32), .O(gate242inter1));
  and2  gate773(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate774(.a(s_32), .O(gate242inter3));
  inv1  gate775(.a(s_33), .O(gate242inter4));
  nand2 gate776(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate777(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate778(.a(G718), .O(gate242inter7));
  inv1  gate779(.a(G730), .O(gate242inter8));
  nand2 gate780(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate781(.a(s_33), .b(gate242inter3), .O(gate242inter10));
  nor2  gate782(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate783(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate784(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1345(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1346(.a(gate244inter0), .b(s_114), .O(gate244inter1));
  and2  gate1347(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1348(.a(s_114), .O(gate244inter3));
  inv1  gate1349(.a(s_115), .O(gate244inter4));
  nand2 gate1350(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1351(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1352(.a(G721), .O(gate244inter7));
  inv1  gate1353(.a(G733), .O(gate244inter8));
  nand2 gate1354(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1355(.a(s_115), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1356(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1357(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1358(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2493(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2494(.a(gate246inter0), .b(s_278), .O(gate246inter1));
  and2  gate2495(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2496(.a(s_278), .O(gate246inter3));
  inv1  gate2497(.a(s_279), .O(gate246inter4));
  nand2 gate2498(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2499(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2500(.a(G724), .O(gate246inter7));
  inv1  gate2501(.a(G736), .O(gate246inter8));
  nand2 gate2502(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2503(.a(s_279), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2504(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2505(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2506(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate897(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate898(.a(gate248inter0), .b(s_50), .O(gate248inter1));
  and2  gate899(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate900(.a(s_50), .O(gate248inter3));
  inv1  gate901(.a(s_51), .O(gate248inter4));
  nand2 gate902(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate903(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate904(.a(G727), .O(gate248inter7));
  inv1  gate905(.a(G739), .O(gate248inter8));
  nand2 gate906(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate907(.a(s_51), .b(gate248inter3), .O(gate248inter10));
  nor2  gate908(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate909(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate910(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2815(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2816(.a(gate249inter0), .b(s_324), .O(gate249inter1));
  and2  gate2817(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2818(.a(s_324), .O(gate249inter3));
  inv1  gate2819(.a(s_325), .O(gate249inter4));
  nand2 gate2820(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2821(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2822(.a(G254), .O(gate249inter7));
  inv1  gate2823(.a(G742), .O(gate249inter8));
  nand2 gate2824(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2825(.a(s_325), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2826(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2827(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2828(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2283(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2284(.a(gate250inter0), .b(s_248), .O(gate250inter1));
  and2  gate2285(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2286(.a(s_248), .O(gate250inter3));
  inv1  gate2287(.a(s_249), .O(gate250inter4));
  nand2 gate2288(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2289(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2290(.a(G706), .O(gate250inter7));
  inv1  gate2291(.a(G742), .O(gate250inter8));
  nand2 gate2292(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2293(.a(s_249), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2294(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2295(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2296(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate995(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate996(.a(gate252inter0), .b(s_64), .O(gate252inter1));
  and2  gate997(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate998(.a(s_64), .O(gate252inter3));
  inv1  gate999(.a(s_65), .O(gate252inter4));
  nand2 gate1000(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1001(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1002(.a(G709), .O(gate252inter7));
  inv1  gate1003(.a(G745), .O(gate252inter8));
  nand2 gate1004(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1005(.a(s_65), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1006(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1007(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1008(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate1093(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1094(.a(gate253inter0), .b(s_78), .O(gate253inter1));
  and2  gate1095(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1096(.a(s_78), .O(gate253inter3));
  inv1  gate1097(.a(s_79), .O(gate253inter4));
  nand2 gate1098(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1099(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1100(.a(G260), .O(gate253inter7));
  inv1  gate1101(.a(G748), .O(gate253inter8));
  nand2 gate1102(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1103(.a(s_79), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1104(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1105(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1106(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2913(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2914(.a(gate256inter0), .b(s_338), .O(gate256inter1));
  and2  gate2915(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2916(.a(s_338), .O(gate256inter3));
  inv1  gate2917(.a(s_339), .O(gate256inter4));
  nand2 gate2918(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2919(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2920(.a(G715), .O(gate256inter7));
  inv1  gate2921(.a(G751), .O(gate256inter8));
  nand2 gate2922(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2923(.a(s_339), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2924(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2925(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2926(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate561(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate562(.a(gate258inter0), .b(s_2), .O(gate258inter1));
  and2  gate563(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate564(.a(s_2), .O(gate258inter3));
  inv1  gate565(.a(s_3), .O(gate258inter4));
  nand2 gate566(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate567(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate568(.a(G756), .O(gate258inter7));
  inv1  gate569(.a(G757), .O(gate258inter8));
  nand2 gate570(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate571(.a(s_3), .b(gate258inter3), .O(gate258inter10));
  nor2  gate572(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate573(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate574(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate2745(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2746(.a(gate259inter0), .b(s_314), .O(gate259inter1));
  and2  gate2747(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2748(.a(s_314), .O(gate259inter3));
  inv1  gate2749(.a(s_315), .O(gate259inter4));
  nand2 gate2750(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2751(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2752(.a(G758), .O(gate259inter7));
  inv1  gate2753(.a(G759), .O(gate259inter8));
  nand2 gate2754(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2755(.a(s_315), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2756(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2757(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2758(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate3123(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate3124(.a(gate260inter0), .b(s_368), .O(gate260inter1));
  and2  gate3125(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate3126(.a(s_368), .O(gate260inter3));
  inv1  gate3127(.a(s_369), .O(gate260inter4));
  nand2 gate3128(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate3129(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate3130(.a(G760), .O(gate260inter7));
  inv1  gate3131(.a(G761), .O(gate260inter8));
  nand2 gate3132(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate3133(.a(s_369), .b(gate260inter3), .O(gate260inter10));
  nor2  gate3134(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate3135(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate3136(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2633(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2634(.a(gate261inter0), .b(s_298), .O(gate261inter1));
  and2  gate2635(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2636(.a(s_298), .O(gate261inter3));
  inv1  gate2637(.a(s_299), .O(gate261inter4));
  nand2 gate2638(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2639(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2640(.a(G762), .O(gate261inter7));
  inv1  gate2641(.a(G763), .O(gate261inter8));
  nand2 gate2642(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2643(.a(s_299), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2644(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2645(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2646(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1597(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1598(.a(gate262inter0), .b(s_150), .O(gate262inter1));
  and2  gate1599(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1600(.a(s_150), .O(gate262inter3));
  inv1  gate1601(.a(s_151), .O(gate262inter4));
  nand2 gate1602(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1603(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1604(.a(G764), .O(gate262inter7));
  inv1  gate1605(.a(G765), .O(gate262inter8));
  nand2 gate1606(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1607(.a(s_151), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1608(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1609(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1610(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1205(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1206(.a(gate270inter0), .b(s_94), .O(gate270inter1));
  and2  gate1207(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1208(.a(s_94), .O(gate270inter3));
  inv1  gate1209(.a(s_95), .O(gate270inter4));
  nand2 gate1210(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1211(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1212(.a(G657), .O(gate270inter7));
  inv1  gate1213(.a(G785), .O(gate270inter8));
  nand2 gate1214(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1215(.a(s_95), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1216(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1217(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1218(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate547(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate548(.a(gate271inter0), .b(s_0), .O(gate271inter1));
  and2  gate549(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate550(.a(s_0), .O(gate271inter3));
  inv1  gate551(.a(s_1), .O(gate271inter4));
  nand2 gate552(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate553(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate554(.a(G660), .O(gate271inter7));
  inv1  gate555(.a(G788), .O(gate271inter8));
  nand2 gate556(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate557(.a(s_1), .b(gate271inter3), .O(gate271inter10));
  nor2  gate558(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate559(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate560(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1331(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1332(.a(gate272inter0), .b(s_112), .O(gate272inter1));
  and2  gate1333(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1334(.a(s_112), .O(gate272inter3));
  inv1  gate1335(.a(s_113), .O(gate272inter4));
  nand2 gate1336(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1337(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1338(.a(G663), .O(gate272inter7));
  inv1  gate1339(.a(G791), .O(gate272inter8));
  nand2 gate1340(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1341(.a(s_113), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1342(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1343(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1344(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate631(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate632(.a(gate273inter0), .b(s_12), .O(gate273inter1));
  and2  gate633(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate634(.a(s_12), .O(gate273inter3));
  inv1  gate635(.a(s_13), .O(gate273inter4));
  nand2 gate636(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate637(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate638(.a(G642), .O(gate273inter7));
  inv1  gate639(.a(G794), .O(gate273inter8));
  nand2 gate640(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate641(.a(s_13), .b(gate273inter3), .O(gate273inter10));
  nor2  gate642(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate643(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate644(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2059(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2060(.a(gate274inter0), .b(s_216), .O(gate274inter1));
  and2  gate2061(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2062(.a(s_216), .O(gate274inter3));
  inv1  gate2063(.a(s_217), .O(gate274inter4));
  nand2 gate2064(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2065(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2066(.a(G770), .O(gate274inter7));
  inv1  gate2067(.a(G794), .O(gate274inter8));
  nand2 gate2068(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2069(.a(s_217), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2070(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2071(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2072(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1051(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1052(.a(gate276inter0), .b(s_72), .O(gate276inter1));
  and2  gate1053(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1054(.a(s_72), .O(gate276inter3));
  inv1  gate1055(.a(s_73), .O(gate276inter4));
  nand2 gate1056(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1057(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1058(.a(G773), .O(gate276inter7));
  inv1  gate1059(.a(G797), .O(gate276inter8));
  nand2 gate1060(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1061(.a(s_73), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1062(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1063(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1064(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate2311(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2312(.a(gate277inter0), .b(s_252), .O(gate277inter1));
  and2  gate2313(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2314(.a(s_252), .O(gate277inter3));
  inv1  gate2315(.a(s_253), .O(gate277inter4));
  nand2 gate2316(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2317(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2318(.a(G648), .O(gate277inter7));
  inv1  gate2319(.a(G800), .O(gate277inter8));
  nand2 gate2320(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2321(.a(s_253), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2322(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2323(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2324(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1359(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1360(.a(gate281inter0), .b(s_116), .O(gate281inter1));
  and2  gate1361(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1362(.a(s_116), .O(gate281inter3));
  inv1  gate1363(.a(s_117), .O(gate281inter4));
  nand2 gate1364(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1365(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1366(.a(G654), .O(gate281inter7));
  inv1  gate1367(.a(G806), .O(gate281inter8));
  nand2 gate1368(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1369(.a(s_117), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1370(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1371(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1372(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1373(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1374(.a(gate283inter0), .b(s_118), .O(gate283inter1));
  and2  gate1375(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1376(.a(s_118), .O(gate283inter3));
  inv1  gate1377(.a(s_119), .O(gate283inter4));
  nand2 gate1378(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1379(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1380(.a(G657), .O(gate283inter7));
  inv1  gate1381(.a(G809), .O(gate283inter8));
  nand2 gate1382(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1383(.a(s_119), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1384(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1385(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1386(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2899(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2900(.a(gate285inter0), .b(s_336), .O(gate285inter1));
  and2  gate2901(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2902(.a(s_336), .O(gate285inter3));
  inv1  gate2903(.a(s_337), .O(gate285inter4));
  nand2 gate2904(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2905(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2906(.a(G660), .O(gate285inter7));
  inv1  gate2907(.a(G812), .O(gate285inter8));
  nand2 gate2908(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2909(.a(s_337), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2910(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2911(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2912(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1443(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1444(.a(gate287inter0), .b(s_128), .O(gate287inter1));
  and2  gate1445(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1446(.a(s_128), .O(gate287inter3));
  inv1  gate1447(.a(s_129), .O(gate287inter4));
  nand2 gate1448(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1449(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1450(.a(G663), .O(gate287inter7));
  inv1  gate1451(.a(G815), .O(gate287inter8));
  nand2 gate1452(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1453(.a(s_129), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1454(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1455(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1456(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate981(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate982(.a(gate289inter0), .b(s_62), .O(gate289inter1));
  and2  gate983(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate984(.a(s_62), .O(gate289inter3));
  inv1  gate985(.a(s_63), .O(gate289inter4));
  nand2 gate986(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate987(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate988(.a(G818), .O(gate289inter7));
  inv1  gate989(.a(G819), .O(gate289inter8));
  nand2 gate990(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate991(.a(s_63), .b(gate289inter3), .O(gate289inter10));
  nor2  gate992(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate993(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate994(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate2325(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2326(.a(gate290inter0), .b(s_254), .O(gate290inter1));
  and2  gate2327(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2328(.a(s_254), .O(gate290inter3));
  inv1  gate2329(.a(s_255), .O(gate290inter4));
  nand2 gate2330(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2331(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2332(.a(G820), .O(gate290inter7));
  inv1  gate2333(.a(G821), .O(gate290inter8));
  nand2 gate2334(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2335(.a(s_255), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2336(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2337(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2338(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1737(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1738(.a(gate292inter0), .b(s_170), .O(gate292inter1));
  and2  gate1739(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1740(.a(s_170), .O(gate292inter3));
  inv1  gate1741(.a(s_171), .O(gate292inter4));
  nand2 gate1742(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1743(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1744(.a(G824), .O(gate292inter7));
  inv1  gate1745(.a(G825), .O(gate292inter8));
  nand2 gate1746(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1747(.a(s_171), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1748(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1749(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1750(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1177(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1178(.a(gate294inter0), .b(s_90), .O(gate294inter1));
  and2  gate1179(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1180(.a(s_90), .O(gate294inter3));
  inv1  gate1181(.a(s_91), .O(gate294inter4));
  nand2 gate1182(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1183(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1184(.a(G832), .O(gate294inter7));
  inv1  gate1185(.a(G833), .O(gate294inter8));
  nand2 gate1186(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1187(.a(s_91), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1188(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1189(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1190(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate2703(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2704(.a(gate295inter0), .b(s_308), .O(gate295inter1));
  and2  gate2705(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2706(.a(s_308), .O(gate295inter3));
  inv1  gate2707(.a(s_309), .O(gate295inter4));
  nand2 gate2708(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2709(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2710(.a(G830), .O(gate295inter7));
  inv1  gate2711(.a(G831), .O(gate295inter8));
  nand2 gate2712(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2713(.a(s_309), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2714(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2715(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2716(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate715(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate716(.a(gate296inter0), .b(s_24), .O(gate296inter1));
  and2  gate717(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate718(.a(s_24), .O(gate296inter3));
  inv1  gate719(.a(s_25), .O(gate296inter4));
  nand2 gate720(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate721(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate722(.a(G826), .O(gate296inter7));
  inv1  gate723(.a(G827), .O(gate296inter8));
  nand2 gate724(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate725(.a(s_25), .b(gate296inter3), .O(gate296inter10));
  nor2  gate726(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate727(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate728(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1415(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1416(.a(gate389inter0), .b(s_124), .O(gate389inter1));
  and2  gate1417(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1418(.a(s_124), .O(gate389inter3));
  inv1  gate1419(.a(s_125), .O(gate389inter4));
  nand2 gate1420(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1421(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1422(.a(G3), .O(gate389inter7));
  inv1  gate1423(.a(G1042), .O(gate389inter8));
  nand2 gate1424(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1425(.a(s_125), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1426(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1427(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1428(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate2185(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2186(.a(gate390inter0), .b(s_234), .O(gate390inter1));
  and2  gate2187(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2188(.a(s_234), .O(gate390inter3));
  inv1  gate2189(.a(s_235), .O(gate390inter4));
  nand2 gate2190(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2191(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2192(.a(G4), .O(gate390inter7));
  inv1  gate2193(.a(G1045), .O(gate390inter8));
  nand2 gate2194(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2195(.a(s_235), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2196(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2197(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2198(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate3095(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate3096(.a(gate391inter0), .b(s_364), .O(gate391inter1));
  and2  gate3097(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate3098(.a(s_364), .O(gate391inter3));
  inv1  gate3099(.a(s_365), .O(gate391inter4));
  nand2 gate3100(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate3101(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate3102(.a(G5), .O(gate391inter7));
  inv1  gate3103(.a(G1048), .O(gate391inter8));
  nand2 gate3104(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate3105(.a(s_365), .b(gate391inter3), .O(gate391inter10));
  nor2  gate3106(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate3107(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate3108(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1933(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1934(.a(gate392inter0), .b(s_198), .O(gate392inter1));
  and2  gate1935(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1936(.a(s_198), .O(gate392inter3));
  inv1  gate1937(.a(s_199), .O(gate392inter4));
  nand2 gate1938(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1939(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1940(.a(G6), .O(gate392inter7));
  inv1  gate1941(.a(G1051), .O(gate392inter8));
  nand2 gate1942(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1943(.a(s_199), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1944(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1945(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1946(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1303(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1304(.a(gate393inter0), .b(s_108), .O(gate393inter1));
  and2  gate1305(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1306(.a(s_108), .O(gate393inter3));
  inv1  gate1307(.a(s_109), .O(gate393inter4));
  nand2 gate1308(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1309(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1310(.a(G7), .O(gate393inter7));
  inv1  gate1311(.a(G1054), .O(gate393inter8));
  nand2 gate1312(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1313(.a(s_109), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1314(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1315(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1316(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2129(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2130(.a(gate394inter0), .b(s_226), .O(gate394inter1));
  and2  gate2131(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2132(.a(s_226), .O(gate394inter3));
  inv1  gate2133(.a(s_227), .O(gate394inter4));
  nand2 gate2134(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2135(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2136(.a(G8), .O(gate394inter7));
  inv1  gate2137(.a(G1057), .O(gate394inter8));
  nand2 gate2138(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2139(.a(s_227), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2140(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2141(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2142(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1765(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1766(.a(gate398inter0), .b(s_174), .O(gate398inter1));
  and2  gate1767(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1768(.a(s_174), .O(gate398inter3));
  inv1  gate1769(.a(s_175), .O(gate398inter4));
  nand2 gate1770(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1771(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1772(.a(G12), .O(gate398inter7));
  inv1  gate1773(.a(G1069), .O(gate398inter8));
  nand2 gate1774(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1775(.a(s_175), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1776(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1777(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1778(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2451(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2452(.a(gate401inter0), .b(s_272), .O(gate401inter1));
  and2  gate2453(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2454(.a(s_272), .O(gate401inter3));
  inv1  gate2455(.a(s_273), .O(gate401inter4));
  nand2 gate2456(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2457(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2458(.a(G15), .O(gate401inter7));
  inv1  gate2459(.a(G1078), .O(gate401inter8));
  nand2 gate2460(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2461(.a(s_273), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2462(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2463(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2464(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1317(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1318(.a(gate404inter0), .b(s_110), .O(gate404inter1));
  and2  gate1319(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1320(.a(s_110), .O(gate404inter3));
  inv1  gate1321(.a(s_111), .O(gate404inter4));
  nand2 gate1322(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1323(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1324(.a(G18), .O(gate404inter7));
  inv1  gate1325(.a(G1087), .O(gate404inter8));
  nand2 gate1326(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1327(.a(s_111), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1328(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1329(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1330(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate2213(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2214(.a(gate405inter0), .b(s_238), .O(gate405inter1));
  and2  gate2215(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2216(.a(s_238), .O(gate405inter3));
  inv1  gate2217(.a(s_239), .O(gate405inter4));
  nand2 gate2218(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2219(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2220(.a(G19), .O(gate405inter7));
  inv1  gate2221(.a(G1090), .O(gate405inter8));
  nand2 gate2222(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2223(.a(s_239), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2224(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2225(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2226(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1989(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1990(.a(gate407inter0), .b(s_206), .O(gate407inter1));
  and2  gate1991(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1992(.a(s_206), .O(gate407inter3));
  inv1  gate1993(.a(s_207), .O(gate407inter4));
  nand2 gate1994(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1995(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1996(.a(G21), .O(gate407inter7));
  inv1  gate1997(.a(G1096), .O(gate407inter8));
  nand2 gate1998(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1999(.a(s_207), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2000(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2001(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2002(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1569(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1570(.a(gate410inter0), .b(s_146), .O(gate410inter1));
  and2  gate1571(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1572(.a(s_146), .O(gate410inter3));
  inv1  gate1573(.a(s_147), .O(gate410inter4));
  nand2 gate1574(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1575(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1576(.a(G24), .O(gate410inter7));
  inv1  gate1577(.a(G1105), .O(gate410inter8));
  nand2 gate1578(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1579(.a(s_147), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1580(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1581(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1582(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1135(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1136(.a(gate413inter0), .b(s_84), .O(gate413inter1));
  and2  gate1137(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1138(.a(s_84), .O(gate413inter3));
  inv1  gate1139(.a(s_85), .O(gate413inter4));
  nand2 gate1140(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1141(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1142(.a(G27), .O(gate413inter7));
  inv1  gate1143(.a(G1114), .O(gate413inter8));
  nand2 gate1144(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1145(.a(s_85), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1146(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1147(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1148(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1023(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1024(.a(gate414inter0), .b(s_68), .O(gate414inter1));
  and2  gate1025(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1026(.a(s_68), .O(gate414inter3));
  inv1  gate1027(.a(s_69), .O(gate414inter4));
  nand2 gate1028(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1029(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1030(.a(G28), .O(gate414inter7));
  inv1  gate1031(.a(G1117), .O(gate414inter8));
  nand2 gate1032(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1033(.a(s_69), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1034(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1035(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1036(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2591(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2592(.a(gate418inter0), .b(s_292), .O(gate418inter1));
  and2  gate2593(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2594(.a(s_292), .O(gate418inter3));
  inv1  gate2595(.a(s_293), .O(gate418inter4));
  nand2 gate2596(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2597(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2598(.a(G32), .O(gate418inter7));
  inv1  gate2599(.a(G1129), .O(gate418inter8));
  nand2 gate2600(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2601(.a(s_293), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2602(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2603(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2604(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1625(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1626(.a(gate420inter0), .b(s_154), .O(gate420inter1));
  and2  gate1627(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1628(.a(s_154), .O(gate420inter3));
  inv1  gate1629(.a(s_155), .O(gate420inter4));
  nand2 gate1630(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1631(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1632(.a(G1036), .O(gate420inter7));
  inv1  gate1633(.a(G1132), .O(gate420inter8));
  nand2 gate1634(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1635(.a(s_155), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1636(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1637(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1638(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2983(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2984(.a(gate421inter0), .b(s_348), .O(gate421inter1));
  and2  gate2985(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2986(.a(s_348), .O(gate421inter3));
  inv1  gate2987(.a(s_349), .O(gate421inter4));
  nand2 gate2988(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2989(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2990(.a(G2), .O(gate421inter7));
  inv1  gate2991(.a(G1135), .O(gate421inter8));
  nand2 gate2992(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2993(.a(s_349), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2994(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2995(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2996(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate799(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate800(.a(gate422inter0), .b(s_36), .O(gate422inter1));
  and2  gate801(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate802(.a(s_36), .O(gate422inter3));
  inv1  gate803(.a(s_37), .O(gate422inter4));
  nand2 gate804(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate805(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate806(.a(G1039), .O(gate422inter7));
  inv1  gate807(.a(G1135), .O(gate422inter8));
  nand2 gate808(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate809(.a(s_37), .b(gate422inter3), .O(gate422inter10));
  nor2  gate810(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate811(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate812(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1611(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1612(.a(gate423inter0), .b(s_152), .O(gate423inter1));
  and2  gate1613(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1614(.a(s_152), .O(gate423inter3));
  inv1  gate1615(.a(s_153), .O(gate423inter4));
  nand2 gate1616(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1617(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1618(.a(G3), .O(gate423inter7));
  inv1  gate1619(.a(G1138), .O(gate423inter8));
  nand2 gate1620(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1621(.a(s_153), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1622(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1623(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1624(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2829(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2830(.a(gate424inter0), .b(s_326), .O(gate424inter1));
  and2  gate2831(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2832(.a(s_326), .O(gate424inter3));
  inv1  gate2833(.a(s_327), .O(gate424inter4));
  nand2 gate2834(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2835(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2836(.a(G1042), .O(gate424inter7));
  inv1  gate2837(.a(G1138), .O(gate424inter8));
  nand2 gate2838(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2839(.a(s_327), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2840(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2841(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2842(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1779(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1780(.a(gate426inter0), .b(s_176), .O(gate426inter1));
  and2  gate1781(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1782(.a(s_176), .O(gate426inter3));
  inv1  gate1783(.a(s_177), .O(gate426inter4));
  nand2 gate1784(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1785(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1786(.a(G1045), .O(gate426inter7));
  inv1  gate1787(.a(G1141), .O(gate426inter8));
  nand2 gate1788(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1789(.a(s_177), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1790(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1791(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1792(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2157(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2158(.a(gate427inter0), .b(s_230), .O(gate427inter1));
  and2  gate2159(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2160(.a(s_230), .O(gate427inter3));
  inv1  gate2161(.a(s_231), .O(gate427inter4));
  nand2 gate2162(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2163(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2164(.a(G5), .O(gate427inter7));
  inv1  gate2165(.a(G1144), .O(gate427inter8));
  nand2 gate2166(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2167(.a(s_231), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2168(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2169(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2170(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1975(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1976(.a(gate430inter0), .b(s_204), .O(gate430inter1));
  and2  gate1977(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1978(.a(s_204), .O(gate430inter3));
  inv1  gate1979(.a(s_205), .O(gate430inter4));
  nand2 gate1980(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1981(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1982(.a(G1051), .O(gate430inter7));
  inv1  gate1983(.a(G1147), .O(gate430inter8));
  nand2 gate1984(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1985(.a(s_205), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1986(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1987(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1988(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate785(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate786(.a(gate438inter0), .b(s_34), .O(gate438inter1));
  and2  gate787(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate788(.a(s_34), .O(gate438inter3));
  inv1  gate789(.a(s_35), .O(gate438inter4));
  nand2 gate790(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate791(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate792(.a(G1063), .O(gate438inter7));
  inv1  gate793(.a(G1159), .O(gate438inter8));
  nand2 gate794(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate795(.a(s_35), .b(gate438inter3), .O(gate438inter10));
  nor2  gate796(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate797(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate798(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1527(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1528(.a(gate439inter0), .b(s_140), .O(gate439inter1));
  and2  gate1529(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1530(.a(s_140), .O(gate439inter3));
  inv1  gate1531(.a(s_141), .O(gate439inter4));
  nand2 gate1532(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1533(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1534(.a(G11), .O(gate439inter7));
  inv1  gate1535(.a(G1162), .O(gate439inter8));
  nand2 gate1536(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1537(.a(s_141), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1538(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1539(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1540(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2423(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2424(.a(gate441inter0), .b(s_268), .O(gate441inter1));
  and2  gate2425(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2426(.a(s_268), .O(gate441inter3));
  inv1  gate2427(.a(s_269), .O(gate441inter4));
  nand2 gate2428(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2429(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2430(.a(G12), .O(gate441inter7));
  inv1  gate2431(.a(G1165), .O(gate441inter8));
  nand2 gate2432(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2433(.a(s_269), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2434(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2435(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2436(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2563(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2564(.a(gate442inter0), .b(s_288), .O(gate442inter1));
  and2  gate2565(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2566(.a(s_288), .O(gate442inter3));
  inv1  gate2567(.a(s_289), .O(gate442inter4));
  nand2 gate2568(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2569(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2570(.a(G1069), .O(gate442inter7));
  inv1  gate2571(.a(G1165), .O(gate442inter8));
  nand2 gate2572(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2573(.a(s_289), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2574(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2575(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2576(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate3039(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate3040(.a(gate444inter0), .b(s_356), .O(gate444inter1));
  and2  gate3041(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate3042(.a(s_356), .O(gate444inter3));
  inv1  gate3043(.a(s_357), .O(gate444inter4));
  nand2 gate3044(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate3045(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate3046(.a(G1072), .O(gate444inter7));
  inv1  gate3047(.a(G1168), .O(gate444inter8));
  nand2 gate3048(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate3049(.a(s_357), .b(gate444inter3), .O(gate444inter10));
  nor2  gate3050(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate3051(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate3052(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1261(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1262(.a(gate449inter0), .b(s_102), .O(gate449inter1));
  and2  gate1263(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1264(.a(s_102), .O(gate449inter3));
  inv1  gate1265(.a(s_103), .O(gate449inter4));
  nand2 gate1266(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1267(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1268(.a(G16), .O(gate449inter7));
  inv1  gate1269(.a(G1177), .O(gate449inter8));
  nand2 gate1270(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1271(.a(s_103), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1272(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1273(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1274(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate687(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate688(.a(gate450inter0), .b(s_20), .O(gate450inter1));
  and2  gate689(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate690(.a(s_20), .O(gate450inter3));
  inv1  gate691(.a(s_21), .O(gate450inter4));
  nand2 gate692(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate693(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate694(.a(G1081), .O(gate450inter7));
  inv1  gate695(.a(G1177), .O(gate450inter8));
  nand2 gate696(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate697(.a(s_21), .b(gate450inter3), .O(gate450inter10));
  nor2  gate698(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate699(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate700(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1149(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1150(.a(gate462inter0), .b(s_86), .O(gate462inter1));
  and2  gate1151(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1152(.a(s_86), .O(gate462inter3));
  inv1  gate1153(.a(s_87), .O(gate462inter4));
  nand2 gate1154(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1155(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1156(.a(G1099), .O(gate462inter7));
  inv1  gate1157(.a(G1195), .O(gate462inter8));
  nand2 gate1158(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1159(.a(s_87), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1160(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1161(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1162(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2521(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2522(.a(gate463inter0), .b(s_282), .O(gate463inter1));
  and2  gate2523(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2524(.a(s_282), .O(gate463inter3));
  inv1  gate2525(.a(s_283), .O(gate463inter4));
  nand2 gate2526(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2527(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2528(.a(G23), .O(gate463inter7));
  inv1  gate2529(.a(G1198), .O(gate463inter8));
  nand2 gate2530(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2531(.a(s_283), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2532(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2533(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2534(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1667(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1668(.a(gate464inter0), .b(s_160), .O(gate464inter1));
  and2  gate1669(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1670(.a(s_160), .O(gate464inter3));
  inv1  gate1671(.a(s_161), .O(gate464inter4));
  nand2 gate1672(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1673(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1674(.a(G1102), .O(gate464inter7));
  inv1  gate1675(.a(G1198), .O(gate464inter8));
  nand2 gate1676(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1677(.a(s_161), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1678(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1679(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1680(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2269(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2270(.a(gate465inter0), .b(s_246), .O(gate465inter1));
  and2  gate2271(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2272(.a(s_246), .O(gate465inter3));
  inv1  gate2273(.a(s_247), .O(gate465inter4));
  nand2 gate2274(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2275(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2276(.a(G24), .O(gate465inter7));
  inv1  gate2277(.a(G1201), .O(gate465inter8));
  nand2 gate2278(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2279(.a(s_247), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2280(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2281(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2282(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1961(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1962(.a(gate468inter0), .b(s_202), .O(gate468inter1));
  and2  gate1963(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1964(.a(s_202), .O(gate468inter3));
  inv1  gate1965(.a(s_203), .O(gate468inter4));
  nand2 gate1966(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1967(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1968(.a(G1108), .O(gate468inter7));
  inv1  gate1969(.a(G1204), .O(gate468inter8));
  nand2 gate1970(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1971(.a(s_203), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1972(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1973(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1974(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate3137(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate3138(.a(gate469inter0), .b(s_370), .O(gate469inter1));
  and2  gate3139(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate3140(.a(s_370), .O(gate469inter3));
  inv1  gate3141(.a(s_371), .O(gate469inter4));
  nand2 gate3142(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate3143(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate3144(.a(G26), .O(gate469inter7));
  inv1  gate3145(.a(G1207), .O(gate469inter8));
  nand2 gate3146(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate3147(.a(s_371), .b(gate469inter3), .O(gate469inter10));
  nor2  gate3148(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate3149(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate3150(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate589(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate590(.a(gate470inter0), .b(s_6), .O(gate470inter1));
  and2  gate591(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate592(.a(s_6), .O(gate470inter3));
  inv1  gate593(.a(s_7), .O(gate470inter4));
  nand2 gate594(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate595(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate596(.a(G1111), .O(gate470inter7));
  inv1  gate597(.a(G1207), .O(gate470inter8));
  nand2 gate598(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate599(.a(s_7), .b(gate470inter3), .O(gate470inter10));
  nor2  gate600(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate601(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate602(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2381(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2382(.a(gate472inter0), .b(s_262), .O(gate472inter1));
  and2  gate2383(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2384(.a(s_262), .O(gate472inter3));
  inv1  gate2385(.a(s_263), .O(gate472inter4));
  nand2 gate2386(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2387(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2388(.a(G1114), .O(gate472inter7));
  inv1  gate2389(.a(G1210), .O(gate472inter8));
  nand2 gate2390(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2391(.a(s_263), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2392(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2393(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2394(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate2605(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2606(.a(gate473inter0), .b(s_294), .O(gate473inter1));
  and2  gate2607(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2608(.a(s_294), .O(gate473inter3));
  inv1  gate2609(.a(s_295), .O(gate473inter4));
  nand2 gate2610(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2611(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2612(.a(G28), .O(gate473inter7));
  inv1  gate2613(.a(G1213), .O(gate473inter8));
  nand2 gate2614(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2615(.a(s_295), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2616(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2617(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2618(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2255(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2256(.a(gate475inter0), .b(s_244), .O(gate475inter1));
  and2  gate2257(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2258(.a(s_244), .O(gate475inter3));
  inv1  gate2259(.a(s_245), .O(gate475inter4));
  nand2 gate2260(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2261(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2262(.a(G29), .O(gate475inter7));
  inv1  gate2263(.a(G1216), .O(gate475inter8));
  nand2 gate2264(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2265(.a(s_245), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2266(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2267(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2268(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1429(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1430(.a(gate483inter0), .b(s_126), .O(gate483inter1));
  and2  gate1431(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1432(.a(s_126), .O(gate483inter3));
  inv1  gate1433(.a(s_127), .O(gate483inter4));
  nand2 gate1434(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1435(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1436(.a(G1228), .O(gate483inter7));
  inv1  gate1437(.a(G1229), .O(gate483inter8));
  nand2 gate1438(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1439(.a(s_127), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1440(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1441(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1442(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2871(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2872(.a(gate485inter0), .b(s_332), .O(gate485inter1));
  and2  gate2873(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2874(.a(s_332), .O(gate485inter3));
  inv1  gate2875(.a(s_333), .O(gate485inter4));
  nand2 gate2876(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2877(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2878(.a(G1232), .O(gate485inter7));
  inv1  gate2879(.a(G1233), .O(gate485inter8));
  nand2 gate2880(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2881(.a(s_333), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2882(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2883(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2884(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate2437(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2438(.a(gate486inter0), .b(s_270), .O(gate486inter1));
  and2  gate2439(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2440(.a(s_270), .O(gate486inter3));
  inv1  gate2441(.a(s_271), .O(gate486inter4));
  nand2 gate2442(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2443(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2444(.a(G1234), .O(gate486inter7));
  inv1  gate2445(.a(G1235), .O(gate486inter8));
  nand2 gate2446(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2447(.a(s_271), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2448(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2449(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2450(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2941(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2942(.a(gate488inter0), .b(s_342), .O(gate488inter1));
  and2  gate2943(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2944(.a(s_342), .O(gate488inter3));
  inv1  gate2945(.a(s_343), .O(gate488inter4));
  nand2 gate2946(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2947(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2948(.a(G1238), .O(gate488inter7));
  inv1  gate2949(.a(G1239), .O(gate488inter8));
  nand2 gate2950(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2951(.a(s_343), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2952(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2953(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2954(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate2017(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2018(.a(gate489inter0), .b(s_210), .O(gate489inter1));
  and2  gate2019(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2020(.a(s_210), .O(gate489inter3));
  inv1  gate2021(.a(s_211), .O(gate489inter4));
  nand2 gate2022(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2023(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2024(.a(G1240), .O(gate489inter7));
  inv1  gate2025(.a(G1241), .O(gate489inter8));
  nand2 gate2026(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2027(.a(s_211), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2028(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2029(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2030(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1723(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1724(.a(gate490inter0), .b(s_168), .O(gate490inter1));
  and2  gate1725(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1726(.a(s_168), .O(gate490inter3));
  inv1  gate1727(.a(s_169), .O(gate490inter4));
  nand2 gate1728(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1729(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1730(.a(G1242), .O(gate490inter7));
  inv1  gate1731(.a(G1243), .O(gate490inter8));
  nand2 gate1732(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1733(.a(s_169), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1734(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1735(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1736(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate2115(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2116(.a(gate491inter0), .b(s_224), .O(gate491inter1));
  and2  gate2117(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2118(.a(s_224), .O(gate491inter3));
  inv1  gate2119(.a(s_225), .O(gate491inter4));
  nand2 gate2120(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2121(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2122(.a(G1244), .O(gate491inter7));
  inv1  gate2123(.a(G1245), .O(gate491inter8));
  nand2 gate2124(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2125(.a(s_225), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2126(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2127(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2128(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1681(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1682(.a(gate492inter0), .b(s_162), .O(gate492inter1));
  and2  gate1683(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1684(.a(s_162), .O(gate492inter3));
  inv1  gate1685(.a(s_163), .O(gate492inter4));
  nand2 gate1686(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1687(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1688(.a(G1246), .O(gate492inter7));
  inv1  gate1689(.a(G1247), .O(gate492inter8));
  nand2 gate1690(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1691(.a(s_163), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1692(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1693(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1694(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1107(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1108(.a(gate493inter0), .b(s_80), .O(gate493inter1));
  and2  gate1109(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1110(.a(s_80), .O(gate493inter3));
  inv1  gate1111(.a(s_81), .O(gate493inter4));
  nand2 gate1112(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1113(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1114(.a(G1248), .O(gate493inter7));
  inv1  gate1115(.a(G1249), .O(gate493inter8));
  nand2 gate1116(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1117(.a(s_81), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1118(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1119(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1120(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1695(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1696(.a(gate494inter0), .b(s_164), .O(gate494inter1));
  and2  gate1697(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1698(.a(s_164), .O(gate494inter3));
  inv1  gate1699(.a(s_165), .O(gate494inter4));
  nand2 gate1700(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1701(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1702(.a(G1250), .O(gate494inter7));
  inv1  gate1703(.a(G1251), .O(gate494inter8));
  nand2 gate1704(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1705(.a(s_165), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1706(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1707(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1708(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2857(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2858(.a(gate495inter0), .b(s_330), .O(gate495inter1));
  and2  gate2859(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2860(.a(s_330), .O(gate495inter3));
  inv1  gate2861(.a(s_331), .O(gate495inter4));
  nand2 gate2862(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2863(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2864(.a(G1252), .O(gate495inter7));
  inv1  gate2865(.a(G1253), .O(gate495inter8));
  nand2 gate2866(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2867(.a(s_331), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2868(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2869(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2870(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate953(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate954(.a(gate498inter0), .b(s_58), .O(gate498inter1));
  and2  gate955(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate956(.a(s_58), .O(gate498inter3));
  inv1  gate957(.a(s_59), .O(gate498inter4));
  nand2 gate958(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate959(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate960(.a(G1258), .O(gate498inter7));
  inv1  gate961(.a(G1259), .O(gate498inter8));
  nand2 gate962(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate963(.a(s_59), .b(gate498inter3), .O(gate498inter10));
  nor2  gate964(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate965(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate966(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate743(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate744(.a(gate505inter0), .b(s_28), .O(gate505inter1));
  and2  gate745(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate746(.a(s_28), .O(gate505inter3));
  inv1  gate747(.a(s_29), .O(gate505inter4));
  nand2 gate748(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate749(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate750(.a(G1272), .O(gate505inter7));
  inv1  gate751(.a(G1273), .O(gate505inter8));
  nand2 gate752(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate753(.a(s_29), .b(gate505inter3), .O(gate505inter10));
  nor2  gate754(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate755(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate756(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate2955(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2956(.a(gate506inter0), .b(s_344), .O(gate506inter1));
  and2  gate2957(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2958(.a(s_344), .O(gate506inter3));
  inv1  gate2959(.a(s_345), .O(gate506inter4));
  nand2 gate2960(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2961(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2962(.a(G1274), .O(gate506inter7));
  inv1  gate2963(.a(G1275), .O(gate506inter8));
  nand2 gate2964(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2965(.a(s_345), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2966(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2967(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2968(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate757(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate758(.a(gate507inter0), .b(s_30), .O(gate507inter1));
  and2  gate759(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate760(.a(s_30), .O(gate507inter3));
  inv1  gate761(.a(s_31), .O(gate507inter4));
  nand2 gate762(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate763(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate764(.a(G1276), .O(gate507inter7));
  inv1  gate765(.a(G1277), .O(gate507inter8));
  nand2 gate766(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate767(.a(s_31), .b(gate507inter3), .O(gate507inter10));
  nor2  gate768(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate769(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate770(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate967(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate968(.a(gate508inter0), .b(s_60), .O(gate508inter1));
  and2  gate969(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate970(.a(s_60), .O(gate508inter3));
  inv1  gate971(.a(s_61), .O(gate508inter4));
  nand2 gate972(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate973(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate974(.a(G1278), .O(gate508inter7));
  inv1  gate975(.a(G1279), .O(gate508inter8));
  nand2 gate976(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate977(.a(s_61), .b(gate508inter3), .O(gate508inter10));
  nor2  gate978(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate979(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate980(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1163(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1164(.a(gate509inter0), .b(s_88), .O(gate509inter1));
  and2  gate1165(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1166(.a(s_88), .O(gate509inter3));
  inv1  gate1167(.a(s_89), .O(gate509inter4));
  nand2 gate1168(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1169(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1170(.a(G1280), .O(gate509inter7));
  inv1  gate1171(.a(G1281), .O(gate509inter8));
  nand2 gate1172(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1173(.a(s_89), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1174(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1175(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1176(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate2031(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2032(.a(gate510inter0), .b(s_212), .O(gate510inter1));
  and2  gate2033(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2034(.a(s_212), .O(gate510inter3));
  inv1  gate2035(.a(s_213), .O(gate510inter4));
  nand2 gate2036(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2037(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2038(.a(G1282), .O(gate510inter7));
  inv1  gate2039(.a(G1283), .O(gate510inter8));
  nand2 gate2040(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2041(.a(s_213), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2042(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2043(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2044(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate617(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate618(.a(gate511inter0), .b(s_10), .O(gate511inter1));
  and2  gate619(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate620(.a(s_10), .O(gate511inter3));
  inv1  gate621(.a(s_11), .O(gate511inter4));
  nand2 gate622(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate623(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate624(.a(G1284), .O(gate511inter7));
  inv1  gate625(.a(G1285), .O(gate511inter8));
  nand2 gate626(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate627(.a(s_11), .b(gate511inter3), .O(gate511inter10));
  nor2  gate628(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate629(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate630(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule