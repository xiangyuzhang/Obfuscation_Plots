module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate673(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate674(.a(gate9inter0), .b(s_18), .O(gate9inter1));
  and2  gate675(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate676(.a(s_18), .O(gate9inter3));
  inv1  gate677(.a(s_19), .O(gate9inter4));
  nand2 gate678(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate679(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate680(.a(G1), .O(gate9inter7));
  inv1  gate681(.a(G2), .O(gate9inter8));
  nand2 gate682(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate683(.a(s_19), .b(gate9inter3), .O(gate9inter10));
  nor2  gate684(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate685(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate686(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1065(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1066(.a(gate23inter0), .b(s_74), .O(gate23inter1));
  and2  gate1067(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1068(.a(s_74), .O(gate23inter3));
  inv1  gate1069(.a(s_75), .O(gate23inter4));
  nand2 gate1070(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1071(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1072(.a(G29), .O(gate23inter7));
  inv1  gate1073(.a(G30), .O(gate23inter8));
  nand2 gate1074(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1075(.a(s_75), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1076(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1077(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1078(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2143(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2144(.a(gate34inter0), .b(s_228), .O(gate34inter1));
  and2  gate2145(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2146(.a(s_228), .O(gate34inter3));
  inv1  gate2147(.a(s_229), .O(gate34inter4));
  nand2 gate2148(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2149(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2150(.a(G25), .O(gate34inter7));
  inv1  gate2151(.a(G29), .O(gate34inter8));
  nand2 gate2152(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2153(.a(s_229), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2154(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2155(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2156(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1471(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1472(.a(gate37inter0), .b(s_132), .O(gate37inter1));
  and2  gate1473(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1474(.a(s_132), .O(gate37inter3));
  inv1  gate1475(.a(s_133), .O(gate37inter4));
  nand2 gate1476(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1477(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1478(.a(G19), .O(gate37inter7));
  inv1  gate1479(.a(G23), .O(gate37inter8));
  nand2 gate1480(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1481(.a(s_133), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1482(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1483(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1484(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1135(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1136(.a(gate42inter0), .b(s_84), .O(gate42inter1));
  and2  gate1137(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1138(.a(s_84), .O(gate42inter3));
  inv1  gate1139(.a(s_85), .O(gate42inter4));
  nand2 gate1140(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1141(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1142(.a(G2), .O(gate42inter7));
  inv1  gate1143(.a(G266), .O(gate42inter8));
  nand2 gate1144(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1145(.a(s_85), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1146(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1147(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1148(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1275(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1276(.a(gate44inter0), .b(s_104), .O(gate44inter1));
  and2  gate1277(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1278(.a(s_104), .O(gate44inter3));
  inv1  gate1279(.a(s_105), .O(gate44inter4));
  nand2 gate1280(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1281(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1282(.a(G4), .O(gate44inter7));
  inv1  gate1283(.a(G269), .O(gate44inter8));
  nand2 gate1284(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1285(.a(s_105), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1286(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1287(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1288(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1317(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1318(.a(gate54inter0), .b(s_110), .O(gate54inter1));
  and2  gate1319(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1320(.a(s_110), .O(gate54inter3));
  inv1  gate1321(.a(s_111), .O(gate54inter4));
  nand2 gate1322(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1323(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1324(.a(G14), .O(gate54inter7));
  inv1  gate1325(.a(G284), .O(gate54inter8));
  nand2 gate1326(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1327(.a(s_111), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1328(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1329(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1330(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate617(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate618(.a(gate58inter0), .b(s_10), .O(gate58inter1));
  and2  gate619(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate620(.a(s_10), .O(gate58inter3));
  inv1  gate621(.a(s_11), .O(gate58inter4));
  nand2 gate622(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate623(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate624(.a(G18), .O(gate58inter7));
  inv1  gate625(.a(G290), .O(gate58inter8));
  nand2 gate626(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate627(.a(s_11), .b(gate58inter3), .O(gate58inter10));
  nor2  gate628(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate629(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate630(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1415(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1416(.a(gate60inter0), .b(s_124), .O(gate60inter1));
  and2  gate1417(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1418(.a(s_124), .O(gate60inter3));
  inv1  gate1419(.a(s_125), .O(gate60inter4));
  nand2 gate1420(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1421(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1422(.a(G20), .O(gate60inter7));
  inv1  gate1423(.a(G293), .O(gate60inter8));
  nand2 gate1424(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1425(.a(s_125), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1426(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1427(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1428(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1863(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1864(.a(gate62inter0), .b(s_188), .O(gate62inter1));
  and2  gate1865(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1866(.a(s_188), .O(gate62inter3));
  inv1  gate1867(.a(s_189), .O(gate62inter4));
  nand2 gate1868(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1869(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1870(.a(G22), .O(gate62inter7));
  inv1  gate1871(.a(G296), .O(gate62inter8));
  nand2 gate1872(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1873(.a(s_189), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1874(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1875(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1876(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1765(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1766(.a(gate63inter0), .b(s_174), .O(gate63inter1));
  and2  gate1767(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1768(.a(s_174), .O(gate63inter3));
  inv1  gate1769(.a(s_175), .O(gate63inter4));
  nand2 gate1770(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1771(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1772(.a(G23), .O(gate63inter7));
  inv1  gate1773(.a(G299), .O(gate63inter8));
  nand2 gate1774(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1775(.a(s_175), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1776(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1777(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1778(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1905(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1906(.a(gate73inter0), .b(s_194), .O(gate73inter1));
  and2  gate1907(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1908(.a(s_194), .O(gate73inter3));
  inv1  gate1909(.a(s_195), .O(gate73inter4));
  nand2 gate1910(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1911(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1912(.a(G1), .O(gate73inter7));
  inv1  gate1913(.a(G314), .O(gate73inter8));
  nand2 gate1914(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1915(.a(s_195), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1916(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1917(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1918(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1331(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1332(.a(gate74inter0), .b(s_112), .O(gate74inter1));
  and2  gate1333(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1334(.a(s_112), .O(gate74inter3));
  inv1  gate1335(.a(s_113), .O(gate74inter4));
  nand2 gate1336(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1337(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1338(.a(G5), .O(gate74inter7));
  inv1  gate1339(.a(G314), .O(gate74inter8));
  nand2 gate1340(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1341(.a(s_113), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1342(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1343(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1344(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate841(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate842(.a(gate75inter0), .b(s_42), .O(gate75inter1));
  and2  gate843(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate844(.a(s_42), .O(gate75inter3));
  inv1  gate845(.a(s_43), .O(gate75inter4));
  nand2 gate846(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate847(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate848(.a(G9), .O(gate75inter7));
  inv1  gate849(.a(G317), .O(gate75inter8));
  nand2 gate850(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate851(.a(s_43), .b(gate75inter3), .O(gate75inter10));
  nor2  gate852(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate853(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate854(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2283(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2284(.a(gate80inter0), .b(s_248), .O(gate80inter1));
  and2  gate2285(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2286(.a(s_248), .O(gate80inter3));
  inv1  gate2287(.a(s_249), .O(gate80inter4));
  nand2 gate2288(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2289(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2290(.a(G14), .O(gate80inter7));
  inv1  gate2291(.a(G323), .O(gate80inter8));
  nand2 gate2292(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2293(.a(s_249), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2294(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2295(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2296(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2129(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2130(.a(gate82inter0), .b(s_226), .O(gate82inter1));
  and2  gate2131(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2132(.a(s_226), .O(gate82inter3));
  inv1  gate2133(.a(s_227), .O(gate82inter4));
  nand2 gate2134(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2135(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2136(.a(G7), .O(gate82inter7));
  inv1  gate2137(.a(G326), .O(gate82inter8));
  nand2 gate2138(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2139(.a(s_227), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2140(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2141(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2142(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1345(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1346(.a(gate84inter0), .b(s_114), .O(gate84inter1));
  and2  gate1347(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1348(.a(s_114), .O(gate84inter3));
  inv1  gate1349(.a(s_115), .O(gate84inter4));
  nand2 gate1350(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1351(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1352(.a(G15), .O(gate84inter7));
  inv1  gate1353(.a(G329), .O(gate84inter8));
  nand2 gate1354(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1355(.a(s_115), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1356(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1357(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1358(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate631(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate632(.a(gate87inter0), .b(s_12), .O(gate87inter1));
  and2  gate633(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate634(.a(s_12), .O(gate87inter3));
  inv1  gate635(.a(s_13), .O(gate87inter4));
  nand2 gate636(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate637(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate638(.a(G12), .O(gate87inter7));
  inv1  gate639(.a(G335), .O(gate87inter8));
  nand2 gate640(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate641(.a(s_13), .b(gate87inter3), .O(gate87inter10));
  nor2  gate642(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate643(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate644(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1625(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1626(.a(gate92inter0), .b(s_154), .O(gate92inter1));
  and2  gate1627(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1628(.a(s_154), .O(gate92inter3));
  inv1  gate1629(.a(s_155), .O(gate92inter4));
  nand2 gate1630(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1631(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1632(.a(G29), .O(gate92inter7));
  inv1  gate1633(.a(G341), .O(gate92inter8));
  nand2 gate1634(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1635(.a(s_155), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1636(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1637(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1638(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1835(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1836(.a(gate96inter0), .b(s_184), .O(gate96inter1));
  and2  gate1837(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1838(.a(s_184), .O(gate96inter3));
  inv1  gate1839(.a(s_185), .O(gate96inter4));
  nand2 gate1840(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1841(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1842(.a(G30), .O(gate96inter7));
  inv1  gate1843(.a(G347), .O(gate96inter8));
  nand2 gate1844(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1845(.a(s_185), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1846(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1847(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1848(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate981(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate982(.a(gate99inter0), .b(s_62), .O(gate99inter1));
  and2  gate983(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate984(.a(s_62), .O(gate99inter3));
  inv1  gate985(.a(s_63), .O(gate99inter4));
  nand2 gate986(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate987(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate988(.a(G27), .O(gate99inter7));
  inv1  gate989(.a(G353), .O(gate99inter8));
  nand2 gate990(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate991(.a(s_63), .b(gate99inter3), .O(gate99inter10));
  nor2  gate992(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate993(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate994(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1499(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1500(.a(gate100inter0), .b(s_136), .O(gate100inter1));
  and2  gate1501(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1502(.a(s_136), .O(gate100inter3));
  inv1  gate1503(.a(s_137), .O(gate100inter4));
  nand2 gate1504(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1505(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1506(.a(G31), .O(gate100inter7));
  inv1  gate1507(.a(G353), .O(gate100inter8));
  nand2 gate1508(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1509(.a(s_137), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1510(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1511(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1512(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1821(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1822(.a(gate109inter0), .b(s_182), .O(gate109inter1));
  and2  gate1823(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1824(.a(s_182), .O(gate109inter3));
  inv1  gate1825(.a(s_183), .O(gate109inter4));
  nand2 gate1826(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1827(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1828(.a(G370), .O(gate109inter7));
  inv1  gate1829(.a(G371), .O(gate109inter8));
  nand2 gate1830(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1831(.a(s_183), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1832(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1833(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1834(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate939(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate940(.a(gate110inter0), .b(s_56), .O(gate110inter1));
  and2  gate941(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate942(.a(s_56), .O(gate110inter3));
  inv1  gate943(.a(s_57), .O(gate110inter4));
  nand2 gate944(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate945(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate946(.a(G372), .O(gate110inter7));
  inv1  gate947(.a(G373), .O(gate110inter8));
  nand2 gate948(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate949(.a(s_57), .b(gate110inter3), .O(gate110inter10));
  nor2  gate950(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate951(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate952(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate869(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate870(.a(gate112inter0), .b(s_46), .O(gate112inter1));
  and2  gate871(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate872(.a(s_46), .O(gate112inter3));
  inv1  gate873(.a(s_47), .O(gate112inter4));
  nand2 gate874(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate875(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate876(.a(G376), .O(gate112inter7));
  inv1  gate877(.a(G377), .O(gate112inter8));
  nand2 gate878(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate879(.a(s_47), .b(gate112inter3), .O(gate112inter10));
  nor2  gate880(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate881(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate882(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate897(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate898(.a(gate122inter0), .b(s_50), .O(gate122inter1));
  and2  gate899(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate900(.a(s_50), .O(gate122inter3));
  inv1  gate901(.a(s_51), .O(gate122inter4));
  nand2 gate902(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate903(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate904(.a(G396), .O(gate122inter7));
  inv1  gate905(.a(G397), .O(gate122inter8));
  nand2 gate906(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate907(.a(s_51), .b(gate122inter3), .O(gate122inter10));
  nor2  gate908(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate909(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate910(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1933(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1934(.a(gate123inter0), .b(s_198), .O(gate123inter1));
  and2  gate1935(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1936(.a(s_198), .O(gate123inter3));
  inv1  gate1937(.a(s_199), .O(gate123inter4));
  nand2 gate1938(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1939(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1940(.a(G398), .O(gate123inter7));
  inv1  gate1941(.a(G399), .O(gate123inter8));
  nand2 gate1942(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1943(.a(s_199), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1944(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1945(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1946(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate813(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate814(.a(gate126inter0), .b(s_38), .O(gate126inter1));
  and2  gate815(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate816(.a(s_38), .O(gate126inter3));
  inv1  gate817(.a(s_39), .O(gate126inter4));
  nand2 gate818(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate819(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate820(.a(G404), .O(gate126inter7));
  inv1  gate821(.a(G405), .O(gate126inter8));
  nand2 gate822(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate823(.a(s_39), .b(gate126inter3), .O(gate126inter10));
  nor2  gate824(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate825(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate826(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1709(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1710(.a(gate128inter0), .b(s_166), .O(gate128inter1));
  and2  gate1711(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1712(.a(s_166), .O(gate128inter3));
  inv1  gate1713(.a(s_167), .O(gate128inter4));
  nand2 gate1714(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1715(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1716(.a(G408), .O(gate128inter7));
  inv1  gate1717(.a(G409), .O(gate128inter8));
  nand2 gate1718(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1719(.a(s_167), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1720(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1721(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1722(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate2255(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2256(.a(gate130inter0), .b(s_244), .O(gate130inter1));
  and2  gate2257(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2258(.a(s_244), .O(gate130inter3));
  inv1  gate2259(.a(s_245), .O(gate130inter4));
  nand2 gate2260(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2261(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2262(.a(G412), .O(gate130inter7));
  inv1  gate2263(.a(G413), .O(gate130inter8));
  nand2 gate2264(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2265(.a(s_245), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2266(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2267(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2268(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate589(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate590(.a(gate134inter0), .b(s_6), .O(gate134inter1));
  and2  gate591(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate592(.a(s_6), .O(gate134inter3));
  inv1  gate593(.a(s_7), .O(gate134inter4));
  nand2 gate594(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate595(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate596(.a(G420), .O(gate134inter7));
  inv1  gate597(.a(G421), .O(gate134inter8));
  nand2 gate598(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate599(.a(s_7), .b(gate134inter3), .O(gate134inter10));
  nor2  gate600(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate601(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate602(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2269(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2270(.a(gate135inter0), .b(s_246), .O(gate135inter1));
  and2  gate2271(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2272(.a(s_246), .O(gate135inter3));
  inv1  gate2273(.a(s_247), .O(gate135inter4));
  nand2 gate2274(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2275(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2276(.a(G422), .O(gate135inter7));
  inv1  gate2277(.a(G423), .O(gate135inter8));
  nand2 gate2278(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2279(.a(s_247), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2280(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2281(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2282(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1891(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1892(.a(gate136inter0), .b(s_192), .O(gate136inter1));
  and2  gate1893(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1894(.a(s_192), .O(gate136inter3));
  inv1  gate1895(.a(s_193), .O(gate136inter4));
  nand2 gate1896(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1897(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1898(.a(G424), .O(gate136inter7));
  inv1  gate1899(.a(G425), .O(gate136inter8));
  nand2 gate1900(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1901(.a(s_193), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1902(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1903(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1904(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1121(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1122(.a(gate141inter0), .b(s_82), .O(gate141inter1));
  and2  gate1123(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1124(.a(s_82), .O(gate141inter3));
  inv1  gate1125(.a(s_83), .O(gate141inter4));
  nand2 gate1126(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1127(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1128(.a(G450), .O(gate141inter7));
  inv1  gate1129(.a(G453), .O(gate141inter8));
  nand2 gate1130(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1131(.a(s_83), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1132(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1133(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1134(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1877(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1878(.a(gate145inter0), .b(s_190), .O(gate145inter1));
  and2  gate1879(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1880(.a(s_190), .O(gate145inter3));
  inv1  gate1881(.a(s_191), .O(gate145inter4));
  nand2 gate1882(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1883(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1884(.a(G474), .O(gate145inter7));
  inv1  gate1885(.a(G477), .O(gate145inter8));
  nand2 gate1886(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1887(.a(s_191), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1888(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1889(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1890(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1359(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1360(.a(gate149inter0), .b(s_116), .O(gate149inter1));
  and2  gate1361(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1362(.a(s_116), .O(gate149inter3));
  inv1  gate1363(.a(s_117), .O(gate149inter4));
  nand2 gate1364(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1365(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1366(.a(G498), .O(gate149inter7));
  inv1  gate1367(.a(G501), .O(gate149inter8));
  nand2 gate1368(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1369(.a(s_117), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1370(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1371(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1372(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1793(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1794(.a(gate150inter0), .b(s_178), .O(gate150inter1));
  and2  gate1795(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1796(.a(s_178), .O(gate150inter3));
  inv1  gate1797(.a(s_179), .O(gate150inter4));
  nand2 gate1798(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1799(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1800(.a(G504), .O(gate150inter7));
  inv1  gate1801(.a(G507), .O(gate150inter8));
  nand2 gate1802(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1803(.a(s_179), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1804(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1805(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1806(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1443(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1444(.a(gate153inter0), .b(s_128), .O(gate153inter1));
  and2  gate1445(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1446(.a(s_128), .O(gate153inter3));
  inv1  gate1447(.a(s_129), .O(gate153inter4));
  nand2 gate1448(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1449(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1450(.a(G426), .O(gate153inter7));
  inv1  gate1451(.a(G522), .O(gate153inter8));
  nand2 gate1452(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1453(.a(s_129), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1454(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1455(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1456(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1009(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1010(.a(gate156inter0), .b(s_66), .O(gate156inter1));
  and2  gate1011(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1012(.a(s_66), .O(gate156inter3));
  inv1  gate1013(.a(s_67), .O(gate156inter4));
  nand2 gate1014(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1015(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1016(.a(G435), .O(gate156inter7));
  inv1  gate1017(.a(G525), .O(gate156inter8));
  nand2 gate1018(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1019(.a(s_67), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1020(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1021(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1022(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2017(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2018(.a(gate157inter0), .b(s_210), .O(gate157inter1));
  and2  gate2019(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2020(.a(s_210), .O(gate157inter3));
  inv1  gate2021(.a(s_211), .O(gate157inter4));
  nand2 gate2022(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2023(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2024(.a(G438), .O(gate157inter7));
  inv1  gate2025(.a(G528), .O(gate157inter8));
  nand2 gate2026(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2027(.a(s_211), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2028(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2029(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2030(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1751(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1752(.a(gate159inter0), .b(s_172), .O(gate159inter1));
  and2  gate1753(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1754(.a(s_172), .O(gate159inter3));
  inv1  gate1755(.a(s_173), .O(gate159inter4));
  nand2 gate1756(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1757(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1758(.a(G444), .O(gate159inter7));
  inv1  gate1759(.a(G531), .O(gate159inter8));
  nand2 gate1760(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1761(.a(s_173), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1762(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1763(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1764(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate799(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate800(.a(gate166inter0), .b(s_36), .O(gate166inter1));
  and2  gate801(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate802(.a(s_36), .O(gate166inter3));
  inv1  gate803(.a(s_37), .O(gate166inter4));
  nand2 gate804(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate805(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate806(.a(G465), .O(gate166inter7));
  inv1  gate807(.a(G540), .O(gate166inter8));
  nand2 gate808(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate809(.a(s_37), .b(gate166inter3), .O(gate166inter10));
  nor2  gate810(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate811(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate812(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1233(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1234(.a(gate175inter0), .b(s_98), .O(gate175inter1));
  and2  gate1235(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1236(.a(s_98), .O(gate175inter3));
  inv1  gate1237(.a(s_99), .O(gate175inter4));
  nand2 gate1238(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1239(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1240(.a(G492), .O(gate175inter7));
  inv1  gate1241(.a(G555), .O(gate175inter8));
  nand2 gate1242(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1243(.a(s_99), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1244(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1245(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1246(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1149(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1150(.a(gate176inter0), .b(s_86), .O(gate176inter1));
  and2  gate1151(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1152(.a(s_86), .O(gate176inter3));
  inv1  gate1153(.a(s_87), .O(gate176inter4));
  nand2 gate1154(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1155(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1156(.a(G495), .O(gate176inter7));
  inv1  gate1157(.a(G555), .O(gate176inter8));
  nand2 gate1158(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1159(.a(s_87), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1160(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1161(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1162(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1975(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1976(.a(gate178inter0), .b(s_204), .O(gate178inter1));
  and2  gate1977(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1978(.a(s_204), .O(gate178inter3));
  inv1  gate1979(.a(s_205), .O(gate178inter4));
  nand2 gate1980(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1981(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1982(.a(G501), .O(gate178inter7));
  inv1  gate1983(.a(G558), .O(gate178inter8));
  nand2 gate1984(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1985(.a(s_205), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1986(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1987(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1988(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2171(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2172(.a(gate184inter0), .b(s_232), .O(gate184inter1));
  and2  gate2173(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2174(.a(s_232), .O(gate184inter3));
  inv1  gate2175(.a(s_233), .O(gate184inter4));
  nand2 gate2176(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2177(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2178(.a(G519), .O(gate184inter7));
  inv1  gate2179(.a(G567), .O(gate184inter8));
  nand2 gate2180(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2181(.a(s_233), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2182(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2183(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2184(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2227(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2228(.a(gate185inter0), .b(s_240), .O(gate185inter1));
  and2  gate2229(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2230(.a(s_240), .O(gate185inter3));
  inv1  gate2231(.a(s_241), .O(gate185inter4));
  nand2 gate2232(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2233(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2234(.a(G570), .O(gate185inter7));
  inv1  gate2235(.a(G571), .O(gate185inter8));
  nand2 gate2236(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2237(.a(s_241), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2238(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2239(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2240(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1177(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1178(.a(gate186inter0), .b(s_90), .O(gate186inter1));
  and2  gate1179(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1180(.a(s_90), .O(gate186inter3));
  inv1  gate1181(.a(s_91), .O(gate186inter4));
  nand2 gate1182(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1183(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1184(.a(G572), .O(gate186inter7));
  inv1  gate1185(.a(G573), .O(gate186inter8));
  nand2 gate1186(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1187(.a(s_91), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1188(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1189(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1190(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1261(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1262(.a(gate187inter0), .b(s_102), .O(gate187inter1));
  and2  gate1263(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1264(.a(s_102), .O(gate187inter3));
  inv1  gate1265(.a(s_103), .O(gate187inter4));
  nand2 gate1266(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1267(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1268(.a(G574), .O(gate187inter7));
  inv1  gate1269(.a(G575), .O(gate187inter8));
  nand2 gate1270(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1271(.a(s_103), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1272(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1273(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1274(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1681(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1682(.a(gate188inter0), .b(s_162), .O(gate188inter1));
  and2  gate1683(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1684(.a(s_162), .O(gate188inter3));
  inv1  gate1685(.a(s_163), .O(gate188inter4));
  nand2 gate1686(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1687(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1688(.a(G576), .O(gate188inter7));
  inv1  gate1689(.a(G577), .O(gate188inter8));
  nand2 gate1690(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1691(.a(s_163), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1692(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1693(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1694(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1583(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1584(.a(gate192inter0), .b(s_148), .O(gate192inter1));
  and2  gate1585(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1586(.a(s_148), .O(gate192inter3));
  inv1  gate1587(.a(s_149), .O(gate192inter4));
  nand2 gate1588(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1589(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1590(.a(G584), .O(gate192inter7));
  inv1  gate1591(.a(G585), .O(gate192inter8));
  nand2 gate1592(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1593(.a(s_149), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1594(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1595(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1596(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1695(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1696(.a(gate198inter0), .b(s_164), .O(gate198inter1));
  and2  gate1697(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1698(.a(s_164), .O(gate198inter3));
  inv1  gate1699(.a(s_165), .O(gate198inter4));
  nand2 gate1700(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1701(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1702(.a(G596), .O(gate198inter7));
  inv1  gate1703(.a(G597), .O(gate198inter8));
  nand2 gate1704(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1705(.a(s_165), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1706(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1707(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1708(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate729(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate730(.a(gate199inter0), .b(s_26), .O(gate199inter1));
  and2  gate731(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate732(.a(s_26), .O(gate199inter3));
  inv1  gate733(.a(s_27), .O(gate199inter4));
  nand2 gate734(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate735(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate736(.a(G598), .O(gate199inter7));
  inv1  gate737(.a(G599), .O(gate199inter8));
  nand2 gate738(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate739(.a(s_27), .b(gate199inter3), .O(gate199inter10));
  nor2  gate740(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate741(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate742(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1037(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1038(.a(gate200inter0), .b(s_70), .O(gate200inter1));
  and2  gate1039(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1040(.a(s_70), .O(gate200inter3));
  inv1  gate1041(.a(s_71), .O(gate200inter4));
  nand2 gate1042(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1043(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1044(.a(G600), .O(gate200inter7));
  inv1  gate1045(.a(G601), .O(gate200inter8));
  nand2 gate1046(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1047(.a(s_71), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1048(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1049(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1050(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1611(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1612(.a(gate204inter0), .b(s_152), .O(gate204inter1));
  and2  gate1613(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1614(.a(s_152), .O(gate204inter3));
  inv1  gate1615(.a(s_153), .O(gate204inter4));
  nand2 gate1616(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1617(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1618(.a(G607), .O(gate204inter7));
  inv1  gate1619(.a(G617), .O(gate204inter8));
  nand2 gate1620(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1621(.a(s_153), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1622(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1623(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1624(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate827(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate828(.a(gate206inter0), .b(s_40), .O(gate206inter1));
  and2  gate829(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate830(.a(s_40), .O(gate206inter3));
  inv1  gate831(.a(s_41), .O(gate206inter4));
  nand2 gate832(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate833(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate834(.a(G632), .O(gate206inter7));
  inv1  gate835(.a(G637), .O(gate206inter8));
  nand2 gate836(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate837(.a(s_41), .b(gate206inter3), .O(gate206inter10));
  nor2  gate838(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate839(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate840(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate967(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate968(.a(gate208inter0), .b(s_60), .O(gate208inter1));
  and2  gate969(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate970(.a(s_60), .O(gate208inter3));
  inv1  gate971(.a(s_61), .O(gate208inter4));
  nand2 gate972(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate973(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate974(.a(G627), .O(gate208inter7));
  inv1  gate975(.a(G637), .O(gate208inter8));
  nand2 gate976(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate977(.a(s_61), .b(gate208inter3), .O(gate208inter10));
  nor2  gate978(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate979(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate980(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate771(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate772(.a(gate210inter0), .b(s_32), .O(gate210inter1));
  and2  gate773(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate774(.a(s_32), .O(gate210inter3));
  inv1  gate775(.a(s_33), .O(gate210inter4));
  nand2 gate776(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate777(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate778(.a(G607), .O(gate210inter7));
  inv1  gate779(.a(G666), .O(gate210inter8));
  nand2 gate780(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate781(.a(s_33), .b(gate210inter3), .O(gate210inter10));
  nor2  gate782(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate783(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate784(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1779(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1780(.a(gate216inter0), .b(s_176), .O(gate216inter1));
  and2  gate1781(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1782(.a(s_176), .O(gate216inter3));
  inv1  gate1783(.a(s_177), .O(gate216inter4));
  nand2 gate1784(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1785(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1786(.a(G617), .O(gate216inter7));
  inv1  gate1787(.a(G675), .O(gate216inter8));
  nand2 gate1788(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1789(.a(s_177), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1790(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1791(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1792(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2059(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2060(.a(gate220inter0), .b(s_216), .O(gate220inter1));
  and2  gate2061(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2062(.a(s_216), .O(gate220inter3));
  inv1  gate2063(.a(s_217), .O(gate220inter4));
  nand2 gate2064(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2065(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2066(.a(G637), .O(gate220inter7));
  inv1  gate2067(.a(G681), .O(gate220inter8));
  nand2 gate2068(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2069(.a(s_217), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2070(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2071(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2072(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate743(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate744(.a(gate224inter0), .b(s_28), .O(gate224inter1));
  and2  gate745(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate746(.a(s_28), .O(gate224inter3));
  inv1  gate747(.a(s_29), .O(gate224inter4));
  nand2 gate748(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate749(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate750(.a(G637), .O(gate224inter7));
  inv1  gate751(.a(G687), .O(gate224inter8));
  nand2 gate752(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate753(.a(s_29), .b(gate224inter3), .O(gate224inter10));
  nor2  gate754(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate755(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate756(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1485(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1486(.a(gate226inter0), .b(s_134), .O(gate226inter1));
  and2  gate1487(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1488(.a(s_134), .O(gate226inter3));
  inv1  gate1489(.a(s_135), .O(gate226inter4));
  nand2 gate1490(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1491(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1492(.a(G692), .O(gate226inter7));
  inv1  gate1493(.a(G693), .O(gate226inter8));
  nand2 gate1494(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1495(.a(s_135), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1496(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1497(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1498(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1093(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1094(.a(gate227inter0), .b(s_78), .O(gate227inter1));
  and2  gate1095(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1096(.a(s_78), .O(gate227inter3));
  inv1  gate1097(.a(s_79), .O(gate227inter4));
  nand2 gate1098(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1099(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1100(.a(G694), .O(gate227inter7));
  inv1  gate1101(.a(G695), .O(gate227inter8));
  nand2 gate1102(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1103(.a(s_79), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1104(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1105(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1106(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1513(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1514(.a(gate228inter0), .b(s_138), .O(gate228inter1));
  and2  gate1515(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1516(.a(s_138), .O(gate228inter3));
  inv1  gate1517(.a(s_139), .O(gate228inter4));
  nand2 gate1518(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1519(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1520(.a(G696), .O(gate228inter7));
  inv1  gate1521(.a(G697), .O(gate228inter8));
  nand2 gate1522(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1523(.a(s_139), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1524(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1525(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1526(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1947(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1948(.a(gate231inter0), .b(s_200), .O(gate231inter1));
  and2  gate1949(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1950(.a(s_200), .O(gate231inter3));
  inv1  gate1951(.a(s_201), .O(gate231inter4));
  nand2 gate1952(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1953(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1954(.a(G702), .O(gate231inter7));
  inv1  gate1955(.a(G703), .O(gate231inter8));
  nand2 gate1956(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1957(.a(s_201), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1958(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1959(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1960(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate2031(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2032(.a(gate235inter0), .b(s_212), .O(gate235inter1));
  and2  gate2033(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2034(.a(s_212), .O(gate235inter3));
  inv1  gate2035(.a(s_213), .O(gate235inter4));
  nand2 gate2036(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2037(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2038(.a(G248), .O(gate235inter7));
  inv1  gate2039(.a(G724), .O(gate235inter8));
  nand2 gate2040(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2041(.a(s_213), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2042(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2043(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2044(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate603(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate604(.a(gate239inter0), .b(s_8), .O(gate239inter1));
  and2  gate605(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate606(.a(s_8), .O(gate239inter3));
  inv1  gate607(.a(s_9), .O(gate239inter4));
  nand2 gate608(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate609(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate610(.a(G260), .O(gate239inter7));
  inv1  gate611(.a(G712), .O(gate239inter8));
  nand2 gate612(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate613(.a(s_9), .b(gate239inter3), .O(gate239inter10));
  nor2  gate614(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate615(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate616(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1051(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1052(.a(gate244inter0), .b(s_72), .O(gate244inter1));
  and2  gate1053(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1054(.a(s_72), .O(gate244inter3));
  inv1  gate1055(.a(s_73), .O(gate244inter4));
  nand2 gate1056(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1057(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1058(.a(G721), .O(gate244inter7));
  inv1  gate1059(.a(G733), .O(gate244inter8));
  nand2 gate1060(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1061(.a(s_73), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1062(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1063(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1064(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate561(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate562(.a(gate245inter0), .b(s_2), .O(gate245inter1));
  and2  gate563(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate564(.a(s_2), .O(gate245inter3));
  inv1  gate565(.a(s_3), .O(gate245inter4));
  nand2 gate566(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate567(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate568(.a(G248), .O(gate245inter7));
  inv1  gate569(.a(G736), .O(gate245inter8));
  nand2 gate570(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate571(.a(s_3), .b(gate245inter3), .O(gate245inter10));
  nor2  gate572(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate573(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate574(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1289(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1290(.a(gate250inter0), .b(s_106), .O(gate250inter1));
  and2  gate1291(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1292(.a(s_106), .O(gate250inter3));
  inv1  gate1293(.a(s_107), .O(gate250inter4));
  nand2 gate1294(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1295(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1296(.a(G706), .O(gate250inter7));
  inv1  gate1297(.a(G742), .O(gate250inter8));
  nand2 gate1298(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1299(.a(s_107), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1300(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1301(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1302(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1849(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1850(.a(gate255inter0), .b(s_186), .O(gate255inter1));
  and2  gate1851(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1852(.a(s_186), .O(gate255inter3));
  inv1  gate1853(.a(s_187), .O(gate255inter4));
  nand2 gate1854(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1855(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1856(.a(G263), .O(gate255inter7));
  inv1  gate1857(.a(G751), .O(gate255inter8));
  nand2 gate1858(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1859(.a(s_187), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1860(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1861(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1862(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2213(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2214(.a(gate262inter0), .b(s_238), .O(gate262inter1));
  and2  gate2215(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2216(.a(s_238), .O(gate262inter3));
  inv1  gate2217(.a(s_239), .O(gate262inter4));
  nand2 gate2218(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2219(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2220(.a(G764), .O(gate262inter7));
  inv1  gate2221(.a(G765), .O(gate262inter8));
  nand2 gate2222(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2223(.a(s_239), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2224(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2225(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2226(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1541(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1542(.a(gate263inter0), .b(s_142), .O(gate263inter1));
  and2  gate1543(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1544(.a(s_142), .O(gate263inter3));
  inv1  gate1545(.a(s_143), .O(gate263inter4));
  nand2 gate1546(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1547(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1548(.a(G766), .O(gate263inter7));
  inv1  gate1549(.a(G767), .O(gate263inter8));
  nand2 gate1550(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1551(.a(s_143), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1552(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1553(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1554(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate995(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate996(.a(gate264inter0), .b(s_64), .O(gate264inter1));
  and2  gate997(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate998(.a(s_64), .O(gate264inter3));
  inv1  gate999(.a(s_65), .O(gate264inter4));
  nand2 gate1000(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1001(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1002(.a(G768), .O(gate264inter7));
  inv1  gate1003(.a(G769), .O(gate264inter8));
  nand2 gate1004(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1005(.a(s_65), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1006(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1007(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1008(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1387(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1388(.a(gate265inter0), .b(s_120), .O(gate265inter1));
  and2  gate1389(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1390(.a(s_120), .O(gate265inter3));
  inv1  gate1391(.a(s_121), .O(gate265inter4));
  nand2 gate1392(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1393(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1394(.a(G642), .O(gate265inter7));
  inv1  gate1395(.a(G770), .O(gate265inter8));
  nand2 gate1396(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1397(.a(s_121), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1398(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1399(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1400(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1163(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1164(.a(gate267inter0), .b(s_88), .O(gate267inter1));
  and2  gate1165(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1166(.a(s_88), .O(gate267inter3));
  inv1  gate1167(.a(s_89), .O(gate267inter4));
  nand2 gate1168(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1169(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1170(.a(G648), .O(gate267inter7));
  inv1  gate1171(.a(G776), .O(gate267inter8));
  nand2 gate1172(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1173(.a(s_89), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1174(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1175(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1176(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1527(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1528(.a(gate268inter0), .b(s_140), .O(gate268inter1));
  and2  gate1529(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1530(.a(s_140), .O(gate268inter3));
  inv1  gate1531(.a(s_141), .O(gate268inter4));
  nand2 gate1532(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1533(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1534(.a(G651), .O(gate268inter7));
  inv1  gate1535(.a(G779), .O(gate268inter8));
  nand2 gate1536(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1537(.a(s_141), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1538(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1539(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1540(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1023(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1024(.a(gate270inter0), .b(s_68), .O(gate270inter1));
  and2  gate1025(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1026(.a(s_68), .O(gate270inter3));
  inv1  gate1027(.a(s_69), .O(gate270inter4));
  nand2 gate1028(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1029(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1030(.a(G657), .O(gate270inter7));
  inv1  gate1031(.a(G785), .O(gate270inter8));
  nand2 gate1032(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1033(.a(s_69), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1034(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1035(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1036(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate659(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate660(.a(gate271inter0), .b(s_16), .O(gate271inter1));
  and2  gate661(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate662(.a(s_16), .O(gate271inter3));
  inv1  gate663(.a(s_17), .O(gate271inter4));
  nand2 gate664(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate665(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate666(.a(G660), .O(gate271inter7));
  inv1  gate667(.a(G788), .O(gate271inter8));
  nand2 gate668(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate669(.a(s_17), .b(gate271inter3), .O(gate271inter10));
  nor2  gate670(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate671(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate672(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate785(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate786(.a(gate274inter0), .b(s_34), .O(gate274inter1));
  and2  gate787(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate788(.a(s_34), .O(gate274inter3));
  inv1  gate789(.a(s_35), .O(gate274inter4));
  nand2 gate790(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate791(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate792(.a(G770), .O(gate274inter7));
  inv1  gate793(.a(G794), .O(gate274inter8));
  nand2 gate794(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate795(.a(s_35), .b(gate274inter3), .O(gate274inter10));
  nor2  gate796(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate797(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate798(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1667(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1668(.a(gate277inter0), .b(s_160), .O(gate277inter1));
  and2  gate1669(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1670(.a(s_160), .O(gate277inter3));
  inv1  gate1671(.a(s_161), .O(gate277inter4));
  nand2 gate1672(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1673(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1674(.a(G648), .O(gate277inter7));
  inv1  gate1675(.a(G800), .O(gate277inter8));
  nand2 gate1676(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1677(.a(s_161), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1678(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1679(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1680(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1107(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1108(.a(gate293inter0), .b(s_80), .O(gate293inter1));
  and2  gate1109(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1110(.a(s_80), .O(gate293inter3));
  inv1  gate1111(.a(s_81), .O(gate293inter4));
  nand2 gate1112(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1113(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1114(.a(G828), .O(gate293inter7));
  inv1  gate1115(.a(G829), .O(gate293inter8));
  nand2 gate1116(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1117(.a(s_81), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1118(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1119(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1120(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2297(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2298(.a(gate296inter0), .b(s_250), .O(gate296inter1));
  and2  gate2299(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2300(.a(s_250), .O(gate296inter3));
  inv1  gate2301(.a(s_251), .O(gate296inter4));
  nand2 gate2302(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2303(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2304(.a(G826), .O(gate296inter7));
  inv1  gate2305(.a(G827), .O(gate296inter8));
  nand2 gate2306(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2307(.a(s_251), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2308(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2309(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2310(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1205(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1206(.a(gate387inter0), .b(s_94), .O(gate387inter1));
  and2  gate1207(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1208(.a(s_94), .O(gate387inter3));
  inv1  gate1209(.a(s_95), .O(gate387inter4));
  nand2 gate1210(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1211(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1212(.a(G1), .O(gate387inter7));
  inv1  gate1213(.a(G1036), .O(gate387inter8));
  nand2 gate1214(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1215(.a(s_95), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1216(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1217(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1218(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate855(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate856(.a(gate389inter0), .b(s_44), .O(gate389inter1));
  and2  gate857(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate858(.a(s_44), .O(gate389inter3));
  inv1  gate859(.a(s_45), .O(gate389inter4));
  nand2 gate860(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate861(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate862(.a(G3), .O(gate389inter7));
  inv1  gate863(.a(G1042), .O(gate389inter8));
  nand2 gate864(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate865(.a(s_45), .b(gate389inter3), .O(gate389inter10));
  nor2  gate866(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate867(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate868(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2045(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2046(.a(gate393inter0), .b(s_214), .O(gate393inter1));
  and2  gate2047(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2048(.a(s_214), .O(gate393inter3));
  inv1  gate2049(.a(s_215), .O(gate393inter4));
  nand2 gate2050(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2051(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2052(.a(G7), .O(gate393inter7));
  inv1  gate2053(.a(G1054), .O(gate393inter8));
  nand2 gate2054(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2055(.a(s_215), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2056(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2057(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2058(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2241(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2242(.a(gate395inter0), .b(s_242), .O(gate395inter1));
  and2  gate2243(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2244(.a(s_242), .O(gate395inter3));
  inv1  gate2245(.a(s_243), .O(gate395inter4));
  nand2 gate2246(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2247(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2248(.a(G9), .O(gate395inter7));
  inv1  gate2249(.a(G1060), .O(gate395inter8));
  nand2 gate2250(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2251(.a(s_243), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2252(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2253(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2254(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate547(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate548(.a(gate399inter0), .b(s_0), .O(gate399inter1));
  and2  gate549(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate550(.a(s_0), .O(gate399inter3));
  inv1  gate551(.a(s_1), .O(gate399inter4));
  nand2 gate552(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate553(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate554(.a(G13), .O(gate399inter7));
  inv1  gate555(.a(G1072), .O(gate399inter8));
  nand2 gate556(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate557(.a(s_1), .b(gate399inter3), .O(gate399inter10));
  nor2  gate558(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate559(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate560(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1247(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1248(.a(gate405inter0), .b(s_100), .O(gate405inter1));
  and2  gate1249(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1250(.a(s_100), .O(gate405inter3));
  inv1  gate1251(.a(s_101), .O(gate405inter4));
  nand2 gate1252(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1253(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1254(.a(G19), .O(gate405inter7));
  inv1  gate1255(.a(G1090), .O(gate405inter8));
  nand2 gate1256(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1257(.a(s_101), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1258(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1259(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1260(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2003(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2004(.a(gate410inter0), .b(s_208), .O(gate410inter1));
  and2  gate2005(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2006(.a(s_208), .O(gate410inter3));
  inv1  gate2007(.a(s_209), .O(gate410inter4));
  nand2 gate2008(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2009(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2010(.a(G24), .O(gate410inter7));
  inv1  gate2011(.a(G1105), .O(gate410inter8));
  nand2 gate2012(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2013(.a(s_209), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2014(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2015(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2016(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1373(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1374(.a(gate413inter0), .b(s_118), .O(gate413inter1));
  and2  gate1375(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1376(.a(s_118), .O(gate413inter3));
  inv1  gate1377(.a(s_119), .O(gate413inter4));
  nand2 gate1378(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1379(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1380(.a(G27), .O(gate413inter7));
  inv1  gate1381(.a(G1114), .O(gate413inter8));
  nand2 gate1382(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1383(.a(s_119), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1384(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1385(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1386(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1079(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1080(.a(gate415inter0), .b(s_76), .O(gate415inter1));
  and2  gate1081(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1082(.a(s_76), .O(gate415inter3));
  inv1  gate1083(.a(s_77), .O(gate415inter4));
  nand2 gate1084(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1085(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1086(.a(G29), .O(gate415inter7));
  inv1  gate1087(.a(G1120), .O(gate415inter8));
  nand2 gate1088(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1089(.a(s_77), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1090(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1091(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1092(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1597(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1598(.a(gate417inter0), .b(s_150), .O(gate417inter1));
  and2  gate1599(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1600(.a(s_150), .O(gate417inter3));
  inv1  gate1601(.a(s_151), .O(gate417inter4));
  nand2 gate1602(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1603(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1604(.a(G31), .O(gate417inter7));
  inv1  gate1605(.a(G1126), .O(gate417inter8));
  nand2 gate1606(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1607(.a(s_151), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1608(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1609(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1610(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2101(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2102(.a(gate422inter0), .b(s_222), .O(gate422inter1));
  and2  gate2103(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2104(.a(s_222), .O(gate422inter3));
  inv1  gate2105(.a(s_223), .O(gate422inter4));
  nand2 gate2106(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2107(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2108(.a(G1039), .O(gate422inter7));
  inv1  gate2109(.a(G1135), .O(gate422inter8));
  nand2 gate2110(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2111(.a(s_223), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2112(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2113(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2114(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate575(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate576(.a(gate424inter0), .b(s_4), .O(gate424inter1));
  and2  gate577(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate578(.a(s_4), .O(gate424inter3));
  inv1  gate579(.a(s_5), .O(gate424inter4));
  nand2 gate580(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate581(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate582(.a(G1042), .O(gate424inter7));
  inv1  gate583(.a(G1138), .O(gate424inter8));
  nand2 gate584(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate585(.a(s_5), .b(gate424inter3), .O(gate424inter10));
  nor2  gate586(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate587(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate588(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1919(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1920(.a(gate432inter0), .b(s_196), .O(gate432inter1));
  and2  gate1921(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1922(.a(s_196), .O(gate432inter3));
  inv1  gate1923(.a(s_197), .O(gate432inter4));
  nand2 gate1924(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1925(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1926(.a(G1054), .O(gate432inter7));
  inv1  gate1927(.a(G1150), .O(gate432inter8));
  nand2 gate1928(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1929(.a(s_197), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1930(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1931(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1932(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1219(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1220(.a(gate434inter0), .b(s_96), .O(gate434inter1));
  and2  gate1221(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1222(.a(s_96), .O(gate434inter3));
  inv1  gate1223(.a(s_97), .O(gate434inter4));
  nand2 gate1224(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1225(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1226(.a(G1057), .O(gate434inter7));
  inv1  gate1227(.a(G1153), .O(gate434inter8));
  nand2 gate1228(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1229(.a(s_97), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1230(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1231(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1232(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1555(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1556(.a(gate436inter0), .b(s_144), .O(gate436inter1));
  and2  gate1557(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1558(.a(s_144), .O(gate436inter3));
  inv1  gate1559(.a(s_145), .O(gate436inter4));
  nand2 gate1560(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1561(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1562(.a(G1060), .O(gate436inter7));
  inv1  gate1563(.a(G1156), .O(gate436inter8));
  nand2 gate1564(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1565(.a(s_145), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1566(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1567(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1568(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate757(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate758(.a(gate439inter0), .b(s_30), .O(gate439inter1));
  and2  gate759(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate760(.a(s_30), .O(gate439inter3));
  inv1  gate761(.a(s_31), .O(gate439inter4));
  nand2 gate762(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate763(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate764(.a(G11), .O(gate439inter7));
  inv1  gate765(.a(G1162), .O(gate439inter8));
  nand2 gate766(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate767(.a(s_31), .b(gate439inter3), .O(gate439inter10));
  nor2  gate768(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate769(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate770(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1639(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1640(.a(gate440inter0), .b(s_156), .O(gate440inter1));
  and2  gate1641(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1642(.a(s_156), .O(gate440inter3));
  inv1  gate1643(.a(s_157), .O(gate440inter4));
  nand2 gate1644(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1645(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1646(.a(G1066), .O(gate440inter7));
  inv1  gate1647(.a(G1162), .O(gate440inter8));
  nand2 gate1648(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1649(.a(s_157), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1650(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1651(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1652(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate953(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate954(.a(gate442inter0), .b(s_58), .O(gate442inter1));
  and2  gate955(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate956(.a(s_58), .O(gate442inter3));
  inv1  gate957(.a(s_59), .O(gate442inter4));
  nand2 gate958(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate959(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate960(.a(G1069), .O(gate442inter7));
  inv1  gate961(.a(G1165), .O(gate442inter8));
  nand2 gate962(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate963(.a(s_59), .b(gate442inter3), .O(gate442inter10));
  nor2  gate964(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate965(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate966(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1989(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1990(.a(gate444inter0), .b(s_206), .O(gate444inter1));
  and2  gate1991(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1992(.a(s_206), .O(gate444inter3));
  inv1  gate1993(.a(s_207), .O(gate444inter4));
  nand2 gate1994(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1995(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1996(.a(G1072), .O(gate444inter7));
  inv1  gate1997(.a(G1168), .O(gate444inter8));
  nand2 gate1998(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1999(.a(s_207), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2000(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2001(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2002(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate883(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate884(.a(gate448inter0), .b(s_48), .O(gate448inter1));
  and2  gate885(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate886(.a(s_48), .O(gate448inter3));
  inv1  gate887(.a(s_49), .O(gate448inter4));
  nand2 gate888(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate889(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate890(.a(G1078), .O(gate448inter7));
  inv1  gate891(.a(G1174), .O(gate448inter8));
  nand2 gate892(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate893(.a(s_49), .b(gate448inter3), .O(gate448inter10));
  nor2  gate894(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate895(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate896(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1191(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1192(.a(gate450inter0), .b(s_92), .O(gate450inter1));
  and2  gate1193(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1194(.a(s_92), .O(gate450inter3));
  inv1  gate1195(.a(s_93), .O(gate450inter4));
  nand2 gate1196(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1197(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1198(.a(G1081), .O(gate450inter7));
  inv1  gate1199(.a(G1177), .O(gate450inter8));
  nand2 gate1200(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1201(.a(s_93), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1202(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1203(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1204(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate645(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate646(.a(gate451inter0), .b(s_14), .O(gate451inter1));
  and2  gate647(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate648(.a(s_14), .O(gate451inter3));
  inv1  gate649(.a(s_15), .O(gate451inter4));
  nand2 gate650(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate651(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate652(.a(G17), .O(gate451inter7));
  inv1  gate653(.a(G1180), .O(gate451inter8));
  nand2 gate654(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate655(.a(s_15), .b(gate451inter3), .O(gate451inter10));
  nor2  gate656(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate657(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate658(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2115(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2116(.a(gate463inter0), .b(s_224), .O(gate463inter1));
  and2  gate2117(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2118(.a(s_224), .O(gate463inter3));
  inv1  gate2119(.a(s_225), .O(gate463inter4));
  nand2 gate2120(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2121(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2122(.a(G23), .O(gate463inter7));
  inv1  gate2123(.a(G1198), .O(gate463inter8));
  nand2 gate2124(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2125(.a(s_225), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2126(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2127(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2128(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1737(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1738(.a(gate464inter0), .b(s_170), .O(gate464inter1));
  and2  gate1739(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1740(.a(s_170), .O(gate464inter3));
  inv1  gate1741(.a(s_171), .O(gate464inter4));
  nand2 gate1742(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1743(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1744(.a(G1102), .O(gate464inter7));
  inv1  gate1745(.a(G1198), .O(gate464inter8));
  nand2 gate1746(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1747(.a(s_171), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1748(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1749(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1750(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1429(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1430(.a(gate466inter0), .b(s_126), .O(gate466inter1));
  and2  gate1431(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1432(.a(s_126), .O(gate466inter3));
  inv1  gate1433(.a(s_127), .O(gate466inter4));
  nand2 gate1434(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1435(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1436(.a(G1105), .O(gate466inter7));
  inv1  gate1437(.a(G1201), .O(gate466inter8));
  nand2 gate1438(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1439(.a(s_127), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1440(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1441(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1442(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1807(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1808(.a(gate467inter0), .b(s_180), .O(gate467inter1));
  and2  gate1809(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1810(.a(s_180), .O(gate467inter3));
  inv1  gate1811(.a(s_181), .O(gate467inter4));
  nand2 gate1812(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1813(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1814(.a(G25), .O(gate467inter7));
  inv1  gate1815(.a(G1204), .O(gate467inter8));
  nand2 gate1816(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1817(.a(s_181), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1818(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1819(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1820(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate715(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate716(.a(gate468inter0), .b(s_24), .O(gate468inter1));
  and2  gate717(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate718(.a(s_24), .O(gate468inter3));
  inv1  gate719(.a(s_25), .O(gate468inter4));
  nand2 gate720(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate721(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate722(.a(G1108), .O(gate468inter7));
  inv1  gate723(.a(G1204), .O(gate468inter8));
  nand2 gate724(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate725(.a(s_25), .b(gate468inter3), .O(gate468inter10));
  nor2  gate726(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate727(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate728(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2199(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2200(.a(gate476inter0), .b(s_236), .O(gate476inter1));
  and2  gate2201(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2202(.a(s_236), .O(gate476inter3));
  inv1  gate2203(.a(s_237), .O(gate476inter4));
  nand2 gate2204(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2205(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2206(.a(G1120), .O(gate476inter7));
  inv1  gate2207(.a(G1216), .O(gate476inter8));
  nand2 gate2208(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2209(.a(s_237), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2210(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2211(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2212(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1961(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1962(.a(gate479inter0), .b(s_202), .O(gate479inter1));
  and2  gate1963(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1964(.a(s_202), .O(gate479inter3));
  inv1  gate1965(.a(s_203), .O(gate479inter4));
  nand2 gate1966(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1967(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1968(.a(G31), .O(gate479inter7));
  inv1  gate1969(.a(G1222), .O(gate479inter8));
  nand2 gate1970(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1971(.a(s_203), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1972(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1973(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1974(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1457(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1458(.a(gate483inter0), .b(s_130), .O(gate483inter1));
  and2  gate1459(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1460(.a(s_130), .O(gate483inter3));
  inv1  gate1461(.a(s_131), .O(gate483inter4));
  nand2 gate1462(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1463(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1464(.a(G1228), .O(gate483inter7));
  inv1  gate1465(.a(G1229), .O(gate483inter8));
  nand2 gate1466(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1467(.a(s_131), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1468(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1469(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1470(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate2157(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate2158(.a(gate484inter0), .b(s_230), .O(gate484inter1));
  and2  gate2159(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate2160(.a(s_230), .O(gate484inter3));
  inv1  gate2161(.a(s_231), .O(gate484inter4));
  nand2 gate2162(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate2163(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate2164(.a(G1230), .O(gate484inter7));
  inv1  gate2165(.a(G1231), .O(gate484inter8));
  nand2 gate2166(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate2167(.a(s_231), .b(gate484inter3), .O(gate484inter10));
  nor2  gate2168(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate2169(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate2170(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate701(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate702(.a(gate486inter0), .b(s_22), .O(gate486inter1));
  and2  gate703(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate704(.a(s_22), .O(gate486inter3));
  inv1  gate705(.a(s_23), .O(gate486inter4));
  nand2 gate706(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate707(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate708(.a(G1234), .O(gate486inter7));
  inv1  gate709(.a(G1235), .O(gate486inter8));
  nand2 gate710(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate711(.a(s_23), .b(gate486inter3), .O(gate486inter10));
  nor2  gate712(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate713(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate714(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2073(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2074(.a(gate488inter0), .b(s_218), .O(gate488inter1));
  and2  gate2075(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2076(.a(s_218), .O(gate488inter3));
  inv1  gate2077(.a(s_219), .O(gate488inter4));
  nand2 gate2078(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2079(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2080(.a(G1238), .O(gate488inter7));
  inv1  gate2081(.a(G1239), .O(gate488inter8));
  nand2 gate2082(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2083(.a(s_219), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2084(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2085(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2086(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate687(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate688(.a(gate494inter0), .b(s_20), .O(gate494inter1));
  and2  gate689(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate690(.a(s_20), .O(gate494inter3));
  inv1  gate691(.a(s_21), .O(gate494inter4));
  nand2 gate692(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate693(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate694(.a(G1250), .O(gate494inter7));
  inv1  gate695(.a(G1251), .O(gate494inter8));
  nand2 gate696(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate697(.a(s_21), .b(gate494inter3), .O(gate494inter10));
  nor2  gate698(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate699(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate700(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1401(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1402(.a(gate496inter0), .b(s_122), .O(gate496inter1));
  and2  gate1403(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1404(.a(s_122), .O(gate496inter3));
  inv1  gate1405(.a(s_123), .O(gate496inter4));
  nand2 gate1406(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1407(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1408(.a(G1254), .O(gate496inter7));
  inv1  gate1409(.a(G1255), .O(gate496inter8));
  nand2 gate1410(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1411(.a(s_123), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1412(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1413(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1414(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate911(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate912(.a(gate500inter0), .b(s_52), .O(gate500inter1));
  and2  gate913(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate914(.a(s_52), .O(gate500inter3));
  inv1  gate915(.a(s_53), .O(gate500inter4));
  nand2 gate916(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate917(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate918(.a(G1262), .O(gate500inter7));
  inv1  gate919(.a(G1263), .O(gate500inter8));
  nand2 gate920(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate921(.a(s_53), .b(gate500inter3), .O(gate500inter10));
  nor2  gate922(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate923(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate924(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1723(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1724(.a(gate502inter0), .b(s_168), .O(gate502inter1));
  and2  gate1725(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1726(.a(s_168), .O(gate502inter3));
  inv1  gate1727(.a(s_169), .O(gate502inter4));
  nand2 gate1728(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1729(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1730(.a(G1266), .O(gate502inter7));
  inv1  gate1731(.a(G1267), .O(gate502inter8));
  nand2 gate1732(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1733(.a(s_169), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1734(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1735(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1736(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate2087(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2088(.a(gate504inter0), .b(s_220), .O(gate504inter1));
  and2  gate2089(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2090(.a(s_220), .O(gate504inter3));
  inv1  gate2091(.a(s_221), .O(gate504inter4));
  nand2 gate2092(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2093(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2094(.a(G1270), .O(gate504inter7));
  inv1  gate2095(.a(G1271), .O(gate504inter8));
  nand2 gate2096(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2097(.a(s_221), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2098(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2099(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2100(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2185(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2186(.a(gate508inter0), .b(s_234), .O(gate508inter1));
  and2  gate2187(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2188(.a(s_234), .O(gate508inter3));
  inv1  gate2189(.a(s_235), .O(gate508inter4));
  nand2 gate2190(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2191(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2192(.a(G1278), .O(gate508inter7));
  inv1  gate2193(.a(G1279), .O(gate508inter8));
  nand2 gate2194(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2195(.a(s_235), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2196(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2197(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2198(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate925(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate926(.a(gate509inter0), .b(s_54), .O(gate509inter1));
  and2  gate927(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate928(.a(s_54), .O(gate509inter3));
  inv1  gate929(.a(s_55), .O(gate509inter4));
  nand2 gate930(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate931(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate932(.a(G1280), .O(gate509inter7));
  inv1  gate933(.a(G1281), .O(gate509inter8));
  nand2 gate934(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate935(.a(s_55), .b(gate509inter3), .O(gate509inter10));
  nor2  gate936(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate937(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate938(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1303(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1304(.a(gate512inter0), .b(s_108), .O(gate512inter1));
  and2  gate1305(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1306(.a(s_108), .O(gate512inter3));
  inv1  gate1307(.a(s_109), .O(gate512inter4));
  nand2 gate1308(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1309(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1310(.a(G1286), .O(gate512inter7));
  inv1  gate1311(.a(G1287), .O(gate512inter8));
  nand2 gate1312(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1313(.a(s_109), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1314(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1315(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1316(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate1653(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1654(.a(gate513inter0), .b(s_158), .O(gate513inter1));
  and2  gate1655(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1656(.a(s_158), .O(gate513inter3));
  inv1  gate1657(.a(s_159), .O(gate513inter4));
  nand2 gate1658(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1659(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1660(.a(G1288), .O(gate513inter7));
  inv1  gate1661(.a(G1289), .O(gate513inter8));
  nand2 gate1662(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1663(.a(s_159), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1664(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1665(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1666(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1569(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1570(.a(gate514inter0), .b(s_146), .O(gate514inter1));
  and2  gate1571(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1572(.a(s_146), .O(gate514inter3));
  inv1  gate1573(.a(s_147), .O(gate514inter4));
  nand2 gate1574(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1575(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1576(.a(G1290), .O(gate514inter7));
  inv1  gate1577(.a(G1291), .O(gate514inter8));
  nand2 gate1578(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1579(.a(s_147), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1580(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1581(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1582(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule