module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate855(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate856(.a(gate12inter0), .b(s_44), .O(gate12inter1));
  and2  gate857(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate858(.a(s_44), .O(gate12inter3));
  inv1  gate859(.a(s_45), .O(gate12inter4));
  nand2 gate860(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate861(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate862(.a(G7), .O(gate12inter7));
  inv1  gate863(.a(G8), .O(gate12inter8));
  nand2 gate864(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate865(.a(s_45), .b(gate12inter3), .O(gate12inter10));
  nor2  gate866(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate867(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate868(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate2773(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2774(.a(gate13inter0), .b(s_318), .O(gate13inter1));
  and2  gate2775(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2776(.a(s_318), .O(gate13inter3));
  inv1  gate2777(.a(s_319), .O(gate13inter4));
  nand2 gate2778(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2779(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2780(.a(G9), .O(gate13inter7));
  inv1  gate2781(.a(G10), .O(gate13inter8));
  nand2 gate2782(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2783(.a(s_319), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2784(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2785(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2786(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1345(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1346(.a(gate16inter0), .b(s_114), .O(gate16inter1));
  and2  gate1347(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1348(.a(s_114), .O(gate16inter3));
  inv1  gate1349(.a(s_115), .O(gate16inter4));
  nand2 gate1350(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1351(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1352(.a(G15), .O(gate16inter7));
  inv1  gate1353(.a(G16), .O(gate16inter8));
  nand2 gate1354(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1355(.a(s_115), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1356(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1357(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1358(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate561(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate562(.a(gate17inter0), .b(s_2), .O(gate17inter1));
  and2  gate563(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate564(.a(s_2), .O(gate17inter3));
  inv1  gate565(.a(s_3), .O(gate17inter4));
  nand2 gate566(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate567(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate568(.a(G17), .O(gate17inter7));
  inv1  gate569(.a(G18), .O(gate17inter8));
  nand2 gate570(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate571(.a(s_3), .b(gate17inter3), .O(gate17inter10));
  nor2  gate572(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate573(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate574(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1919(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1920(.a(gate23inter0), .b(s_196), .O(gate23inter1));
  and2  gate1921(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1922(.a(s_196), .O(gate23inter3));
  inv1  gate1923(.a(s_197), .O(gate23inter4));
  nand2 gate1924(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1925(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1926(.a(G29), .O(gate23inter7));
  inv1  gate1927(.a(G30), .O(gate23inter8));
  nand2 gate1928(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1929(.a(s_197), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1930(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1931(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1932(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2227(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2228(.a(gate24inter0), .b(s_240), .O(gate24inter1));
  and2  gate2229(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2230(.a(s_240), .O(gate24inter3));
  inv1  gate2231(.a(s_241), .O(gate24inter4));
  nand2 gate2232(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2233(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2234(.a(G31), .O(gate24inter7));
  inv1  gate2235(.a(G32), .O(gate24inter8));
  nand2 gate2236(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2237(.a(s_241), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2238(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2239(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2240(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1247(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1248(.a(gate27inter0), .b(s_100), .O(gate27inter1));
  and2  gate1249(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1250(.a(s_100), .O(gate27inter3));
  inv1  gate1251(.a(s_101), .O(gate27inter4));
  nand2 gate1252(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1253(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1254(.a(G2), .O(gate27inter7));
  inv1  gate1255(.a(G6), .O(gate27inter8));
  nand2 gate1256(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1257(.a(s_101), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1258(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1259(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1260(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2143(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2144(.a(gate29inter0), .b(s_228), .O(gate29inter1));
  and2  gate2145(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2146(.a(s_228), .O(gate29inter3));
  inv1  gate2147(.a(s_229), .O(gate29inter4));
  nand2 gate2148(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2149(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2150(.a(G3), .O(gate29inter7));
  inv1  gate2151(.a(G7), .O(gate29inter8));
  nand2 gate2152(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2153(.a(s_229), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2154(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2155(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2156(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2871(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2872(.a(gate30inter0), .b(s_332), .O(gate30inter1));
  and2  gate2873(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2874(.a(s_332), .O(gate30inter3));
  inv1  gate2875(.a(s_333), .O(gate30inter4));
  nand2 gate2876(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2877(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2878(.a(G11), .O(gate30inter7));
  inv1  gate2879(.a(G15), .O(gate30inter8));
  nand2 gate2880(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2881(.a(s_333), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2882(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2883(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2884(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1821(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1822(.a(gate31inter0), .b(s_182), .O(gate31inter1));
  and2  gate1823(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1824(.a(s_182), .O(gate31inter3));
  inv1  gate1825(.a(s_183), .O(gate31inter4));
  nand2 gate1826(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1827(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1828(.a(G4), .O(gate31inter7));
  inv1  gate1829(.a(G8), .O(gate31inter8));
  nand2 gate1830(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1831(.a(s_183), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1832(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1833(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1834(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate827(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate828(.a(gate32inter0), .b(s_40), .O(gate32inter1));
  and2  gate829(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate830(.a(s_40), .O(gate32inter3));
  inv1  gate831(.a(s_41), .O(gate32inter4));
  nand2 gate832(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate833(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate834(.a(G12), .O(gate32inter7));
  inv1  gate835(.a(G16), .O(gate32inter8));
  nand2 gate836(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate837(.a(s_41), .b(gate32inter3), .O(gate32inter10));
  nor2  gate838(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate839(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate840(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate2661(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2662(.a(gate33inter0), .b(s_302), .O(gate33inter1));
  and2  gate2663(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2664(.a(s_302), .O(gate33inter3));
  inv1  gate2665(.a(s_303), .O(gate33inter4));
  nand2 gate2666(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2667(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2668(.a(G17), .O(gate33inter7));
  inv1  gate2669(.a(G21), .O(gate33inter8));
  nand2 gate2670(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2671(.a(s_303), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2672(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2673(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2674(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2045(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2046(.a(gate36inter0), .b(s_214), .O(gate36inter1));
  and2  gate2047(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2048(.a(s_214), .O(gate36inter3));
  inv1  gate2049(.a(s_215), .O(gate36inter4));
  nand2 gate2050(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2051(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2052(.a(G26), .O(gate36inter7));
  inv1  gate2053(.a(G30), .O(gate36inter8));
  nand2 gate2054(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2055(.a(s_215), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2056(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2057(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2058(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1401(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1402(.a(gate37inter0), .b(s_122), .O(gate37inter1));
  and2  gate1403(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1404(.a(s_122), .O(gate37inter3));
  inv1  gate1405(.a(s_123), .O(gate37inter4));
  nand2 gate1406(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1407(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1408(.a(G19), .O(gate37inter7));
  inv1  gate1409(.a(G23), .O(gate37inter8));
  nand2 gate1410(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1411(.a(s_123), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1412(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1413(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1414(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate2521(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2522(.a(gate38inter0), .b(s_282), .O(gate38inter1));
  and2  gate2523(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2524(.a(s_282), .O(gate38inter3));
  inv1  gate2525(.a(s_283), .O(gate38inter4));
  nand2 gate2526(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2527(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2528(.a(G27), .O(gate38inter7));
  inv1  gate2529(.a(G31), .O(gate38inter8));
  nand2 gate2530(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2531(.a(s_283), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2532(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2533(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2534(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2563(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2564(.a(gate39inter0), .b(s_288), .O(gate39inter1));
  and2  gate2565(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2566(.a(s_288), .O(gate39inter3));
  inv1  gate2567(.a(s_289), .O(gate39inter4));
  nand2 gate2568(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2569(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2570(.a(G20), .O(gate39inter7));
  inv1  gate2571(.a(G24), .O(gate39inter8));
  nand2 gate2572(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2573(.a(s_289), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2574(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2575(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2576(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1877(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1878(.a(gate44inter0), .b(s_190), .O(gate44inter1));
  and2  gate1879(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1880(.a(s_190), .O(gate44inter3));
  inv1  gate1881(.a(s_191), .O(gate44inter4));
  nand2 gate1882(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1883(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1884(.a(G4), .O(gate44inter7));
  inv1  gate1885(.a(G269), .O(gate44inter8));
  nand2 gate1886(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1887(.a(s_191), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1888(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1889(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1890(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2745(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2746(.a(gate47inter0), .b(s_314), .O(gate47inter1));
  and2  gate2747(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2748(.a(s_314), .O(gate47inter3));
  inv1  gate2749(.a(s_315), .O(gate47inter4));
  nand2 gate2750(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2751(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2752(.a(G7), .O(gate47inter7));
  inv1  gate2753(.a(G275), .O(gate47inter8));
  nand2 gate2754(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2755(.a(s_315), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2756(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2757(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2758(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate953(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate954(.a(gate48inter0), .b(s_58), .O(gate48inter1));
  and2  gate955(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate956(.a(s_58), .O(gate48inter3));
  inv1  gate957(.a(s_59), .O(gate48inter4));
  nand2 gate958(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate959(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate960(.a(G8), .O(gate48inter7));
  inv1  gate961(.a(G275), .O(gate48inter8));
  nand2 gate962(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate963(.a(s_59), .b(gate48inter3), .O(gate48inter10));
  nor2  gate964(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate965(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate966(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2339(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2340(.a(gate49inter0), .b(s_256), .O(gate49inter1));
  and2  gate2341(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2342(.a(s_256), .O(gate49inter3));
  inv1  gate2343(.a(s_257), .O(gate49inter4));
  nand2 gate2344(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2345(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2346(.a(G9), .O(gate49inter7));
  inv1  gate2347(.a(G278), .O(gate49inter8));
  nand2 gate2348(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2349(.a(s_257), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2350(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2351(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2352(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2381(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2382(.a(gate50inter0), .b(s_262), .O(gate50inter1));
  and2  gate2383(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2384(.a(s_262), .O(gate50inter3));
  inv1  gate2385(.a(s_263), .O(gate50inter4));
  nand2 gate2386(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2387(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2388(.a(G10), .O(gate50inter7));
  inv1  gate2389(.a(G278), .O(gate50inter8));
  nand2 gate2390(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2391(.a(s_263), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2392(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2393(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2394(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate3193(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate3194(.a(gate56inter0), .b(s_378), .O(gate56inter1));
  and2  gate3195(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate3196(.a(s_378), .O(gate56inter3));
  inv1  gate3197(.a(s_379), .O(gate56inter4));
  nand2 gate3198(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate3199(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate3200(.a(G16), .O(gate56inter7));
  inv1  gate3201(.a(G287), .O(gate56inter8));
  nand2 gate3202(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate3203(.a(s_379), .b(gate56inter3), .O(gate56inter10));
  nor2  gate3204(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate3205(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate3206(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1429(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1430(.a(gate60inter0), .b(s_126), .O(gate60inter1));
  and2  gate1431(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1432(.a(s_126), .O(gate60inter3));
  inv1  gate1433(.a(s_127), .O(gate60inter4));
  nand2 gate1434(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1435(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1436(.a(G20), .O(gate60inter7));
  inv1  gate1437(.a(G293), .O(gate60inter8));
  nand2 gate1438(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1439(.a(s_127), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1440(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1441(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1442(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2171(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2172(.a(gate62inter0), .b(s_232), .O(gate62inter1));
  and2  gate2173(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2174(.a(s_232), .O(gate62inter3));
  inv1  gate2175(.a(s_233), .O(gate62inter4));
  nand2 gate2176(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2177(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2178(.a(G22), .O(gate62inter7));
  inv1  gate2179(.a(G296), .O(gate62inter8));
  nand2 gate2180(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2181(.a(s_233), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2182(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2183(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2184(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1695(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1696(.a(gate64inter0), .b(s_164), .O(gate64inter1));
  and2  gate1697(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1698(.a(s_164), .O(gate64inter3));
  inv1  gate1699(.a(s_165), .O(gate64inter4));
  nand2 gate1700(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1701(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1702(.a(G24), .O(gate64inter7));
  inv1  gate1703(.a(G299), .O(gate64inter8));
  nand2 gate1704(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1705(.a(s_165), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1706(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1707(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1708(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2241(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2242(.a(gate66inter0), .b(s_242), .O(gate66inter1));
  and2  gate2243(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2244(.a(s_242), .O(gate66inter3));
  inv1  gate2245(.a(s_243), .O(gate66inter4));
  nand2 gate2246(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2247(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2248(.a(G26), .O(gate66inter7));
  inv1  gate2249(.a(G302), .O(gate66inter8));
  nand2 gate2250(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2251(.a(s_243), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2252(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2253(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2254(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2703(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2704(.a(gate68inter0), .b(s_308), .O(gate68inter1));
  and2  gate2705(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2706(.a(s_308), .O(gate68inter3));
  inv1  gate2707(.a(s_309), .O(gate68inter4));
  nand2 gate2708(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2709(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2710(.a(G28), .O(gate68inter7));
  inv1  gate2711(.a(G305), .O(gate68inter8));
  nand2 gate2712(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2713(.a(s_309), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2714(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2715(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2716(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate2017(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2018(.a(gate69inter0), .b(s_210), .O(gate69inter1));
  and2  gate2019(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2020(.a(s_210), .O(gate69inter3));
  inv1  gate2021(.a(s_211), .O(gate69inter4));
  nand2 gate2022(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2023(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2024(.a(G29), .O(gate69inter7));
  inv1  gate2025(.a(G308), .O(gate69inter8));
  nand2 gate2026(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2027(.a(s_211), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2028(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2029(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2030(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate995(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate996(.a(gate73inter0), .b(s_64), .O(gate73inter1));
  and2  gate997(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate998(.a(s_64), .O(gate73inter3));
  inv1  gate999(.a(s_65), .O(gate73inter4));
  nand2 gate1000(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1001(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1002(.a(G1), .O(gate73inter7));
  inv1  gate1003(.a(G314), .O(gate73inter8));
  nand2 gate1004(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1005(.a(s_65), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1006(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1007(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1008(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate2507(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2508(.a(gate75inter0), .b(s_280), .O(gate75inter1));
  and2  gate2509(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2510(.a(s_280), .O(gate75inter3));
  inv1  gate2511(.a(s_281), .O(gate75inter4));
  nand2 gate2512(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2513(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2514(.a(G9), .O(gate75inter7));
  inv1  gate2515(.a(G317), .O(gate75inter8));
  nand2 gate2516(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2517(.a(s_281), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2518(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2519(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2520(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1457(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1458(.a(gate76inter0), .b(s_130), .O(gate76inter1));
  and2  gate1459(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1460(.a(s_130), .O(gate76inter3));
  inv1  gate1461(.a(s_131), .O(gate76inter4));
  nand2 gate1462(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1463(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1464(.a(G13), .O(gate76inter7));
  inv1  gate1465(.a(G317), .O(gate76inter8));
  nand2 gate1466(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1467(.a(s_131), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1468(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1469(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1470(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1261(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1262(.a(gate80inter0), .b(s_102), .O(gate80inter1));
  and2  gate1263(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1264(.a(s_102), .O(gate80inter3));
  inv1  gate1265(.a(s_103), .O(gate80inter4));
  nand2 gate1266(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1267(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1268(.a(G14), .O(gate80inter7));
  inv1  gate1269(.a(G323), .O(gate80inter8));
  nand2 gate1270(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1271(.a(s_103), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1272(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1273(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1274(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1415(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1416(.a(gate86inter0), .b(s_124), .O(gate86inter1));
  and2  gate1417(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1418(.a(s_124), .O(gate86inter3));
  inv1  gate1419(.a(s_125), .O(gate86inter4));
  nand2 gate1420(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1421(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1422(.a(G8), .O(gate86inter7));
  inv1  gate1423(.a(G332), .O(gate86inter8));
  nand2 gate1424(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1425(.a(s_125), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1426(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1427(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1428(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1793(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1794(.a(gate88inter0), .b(s_178), .O(gate88inter1));
  and2  gate1795(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1796(.a(s_178), .O(gate88inter3));
  inv1  gate1797(.a(s_179), .O(gate88inter4));
  nand2 gate1798(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1799(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1800(.a(G16), .O(gate88inter7));
  inv1  gate1801(.a(G335), .O(gate88inter8));
  nand2 gate1802(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1803(.a(s_179), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1804(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1805(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1806(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2885(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2886(.a(gate92inter0), .b(s_334), .O(gate92inter1));
  and2  gate2887(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2888(.a(s_334), .O(gate92inter3));
  inv1  gate2889(.a(s_335), .O(gate92inter4));
  nand2 gate2890(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2891(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2892(.a(G29), .O(gate92inter7));
  inv1  gate2893(.a(G341), .O(gate92inter8));
  nand2 gate2894(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2895(.a(s_335), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2896(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2897(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2898(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate2297(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2298(.a(gate93inter0), .b(s_250), .O(gate93inter1));
  and2  gate2299(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2300(.a(s_250), .O(gate93inter3));
  inv1  gate2301(.a(s_251), .O(gate93inter4));
  nand2 gate2302(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2303(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2304(.a(G18), .O(gate93inter7));
  inv1  gate2305(.a(G344), .O(gate93inter8));
  nand2 gate2306(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2307(.a(s_251), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2308(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2309(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2310(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2675(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2676(.a(gate97inter0), .b(s_304), .O(gate97inter1));
  and2  gate2677(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2678(.a(s_304), .O(gate97inter3));
  inv1  gate2679(.a(s_305), .O(gate97inter4));
  nand2 gate2680(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2681(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2682(.a(G19), .O(gate97inter7));
  inv1  gate2683(.a(G350), .O(gate97inter8));
  nand2 gate2684(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2685(.a(s_305), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2686(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2687(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2688(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate3025(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate3026(.a(gate98inter0), .b(s_354), .O(gate98inter1));
  and2  gate3027(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate3028(.a(s_354), .O(gate98inter3));
  inv1  gate3029(.a(s_355), .O(gate98inter4));
  nand2 gate3030(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate3031(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate3032(.a(G23), .O(gate98inter7));
  inv1  gate3033(.a(G350), .O(gate98inter8));
  nand2 gate3034(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate3035(.a(s_355), .b(gate98inter3), .O(gate98inter10));
  nor2  gate3036(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate3037(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate3038(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2759(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2760(.a(gate99inter0), .b(s_316), .O(gate99inter1));
  and2  gate2761(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2762(.a(s_316), .O(gate99inter3));
  inv1  gate2763(.a(s_317), .O(gate99inter4));
  nand2 gate2764(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2765(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2766(.a(G27), .O(gate99inter7));
  inv1  gate2767(.a(G353), .O(gate99inter8));
  nand2 gate2768(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2769(.a(s_317), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2770(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2771(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2772(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1723(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1724(.a(gate101inter0), .b(s_168), .O(gate101inter1));
  and2  gate1725(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1726(.a(s_168), .O(gate101inter3));
  inv1  gate1727(.a(s_169), .O(gate101inter4));
  nand2 gate1728(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1729(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1730(.a(G20), .O(gate101inter7));
  inv1  gate1731(.a(G356), .O(gate101inter8));
  nand2 gate1732(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1733(.a(s_169), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1734(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1735(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1736(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1639(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1640(.a(gate102inter0), .b(s_156), .O(gate102inter1));
  and2  gate1641(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1642(.a(s_156), .O(gate102inter3));
  inv1  gate1643(.a(s_157), .O(gate102inter4));
  nand2 gate1644(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1645(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1646(.a(G24), .O(gate102inter7));
  inv1  gate1647(.a(G356), .O(gate102inter8));
  nand2 gate1648(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1649(.a(s_157), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1650(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1651(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1652(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2185(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2186(.a(gate104inter0), .b(s_234), .O(gate104inter1));
  and2  gate2187(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2188(.a(s_234), .O(gate104inter3));
  inv1  gate2189(.a(s_235), .O(gate104inter4));
  nand2 gate2190(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2191(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2192(.a(G32), .O(gate104inter7));
  inv1  gate2193(.a(G359), .O(gate104inter8));
  nand2 gate2194(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2195(.a(s_235), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2196(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2197(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2198(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate743(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate744(.a(gate106inter0), .b(s_28), .O(gate106inter1));
  and2  gate745(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate746(.a(s_28), .O(gate106inter3));
  inv1  gate747(.a(s_29), .O(gate106inter4));
  nand2 gate748(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate749(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate750(.a(G364), .O(gate106inter7));
  inv1  gate751(.a(G365), .O(gate106inter8));
  nand2 gate752(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate753(.a(s_29), .b(gate106inter3), .O(gate106inter10));
  nor2  gate754(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate755(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate756(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate981(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate982(.a(gate110inter0), .b(s_62), .O(gate110inter1));
  and2  gate983(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate984(.a(s_62), .O(gate110inter3));
  inv1  gate985(.a(s_63), .O(gate110inter4));
  nand2 gate986(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate987(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate988(.a(G372), .O(gate110inter7));
  inv1  gate989(.a(G373), .O(gate110inter8));
  nand2 gate990(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate991(.a(s_63), .b(gate110inter3), .O(gate110inter10));
  nor2  gate992(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate993(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate994(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate3137(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate3138(.a(gate111inter0), .b(s_370), .O(gate111inter1));
  and2  gate3139(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate3140(.a(s_370), .O(gate111inter3));
  inv1  gate3141(.a(s_371), .O(gate111inter4));
  nand2 gate3142(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate3143(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate3144(.a(G374), .O(gate111inter7));
  inv1  gate3145(.a(G375), .O(gate111inter8));
  nand2 gate3146(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate3147(.a(s_371), .b(gate111inter3), .O(gate111inter10));
  nor2  gate3148(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate3149(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate3150(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1681(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1682(.a(gate114inter0), .b(s_162), .O(gate114inter1));
  and2  gate1683(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1684(.a(s_162), .O(gate114inter3));
  inv1  gate1685(.a(s_163), .O(gate114inter4));
  nand2 gate1686(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1687(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1688(.a(G380), .O(gate114inter7));
  inv1  gate1689(.a(G381), .O(gate114inter8));
  nand2 gate1690(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1691(.a(s_163), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1692(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1693(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1694(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2073(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2074(.a(gate117inter0), .b(s_218), .O(gate117inter1));
  and2  gate2075(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2076(.a(s_218), .O(gate117inter3));
  inv1  gate2077(.a(s_219), .O(gate117inter4));
  nand2 gate2078(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2079(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2080(.a(G386), .O(gate117inter7));
  inv1  gate2081(.a(G387), .O(gate117inter8));
  nand2 gate2082(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2083(.a(s_219), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2084(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2085(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2086(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2969(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2970(.a(gate119inter0), .b(s_346), .O(gate119inter1));
  and2  gate2971(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2972(.a(s_346), .O(gate119inter3));
  inv1  gate2973(.a(s_347), .O(gate119inter4));
  nand2 gate2974(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2975(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2976(.a(G390), .O(gate119inter7));
  inv1  gate2977(.a(G391), .O(gate119inter8));
  nand2 gate2978(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2979(.a(s_347), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2980(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2981(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2982(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2129(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2130(.a(gate124inter0), .b(s_226), .O(gate124inter1));
  and2  gate2131(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2132(.a(s_226), .O(gate124inter3));
  inv1  gate2133(.a(s_227), .O(gate124inter4));
  nand2 gate2134(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2135(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2136(.a(G400), .O(gate124inter7));
  inv1  gate2137(.a(G401), .O(gate124inter8));
  nand2 gate2138(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2139(.a(s_227), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2140(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2141(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2142(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1121(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1122(.a(gate125inter0), .b(s_82), .O(gate125inter1));
  and2  gate1123(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1124(.a(s_82), .O(gate125inter3));
  inv1  gate1125(.a(s_83), .O(gate125inter4));
  nand2 gate1126(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1127(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1128(.a(G402), .O(gate125inter7));
  inv1  gate1129(.a(G403), .O(gate125inter8));
  nand2 gate1130(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1131(.a(s_83), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1132(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1133(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1134(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate2549(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2550(.a(gate130inter0), .b(s_286), .O(gate130inter1));
  and2  gate2551(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2552(.a(s_286), .O(gate130inter3));
  inv1  gate2553(.a(s_287), .O(gate130inter4));
  nand2 gate2554(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2555(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2556(.a(G412), .O(gate130inter7));
  inv1  gate2557(.a(G413), .O(gate130inter8));
  nand2 gate2558(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2559(.a(s_287), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2560(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2561(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2562(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2353(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2354(.a(gate131inter0), .b(s_258), .O(gate131inter1));
  and2  gate2355(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2356(.a(s_258), .O(gate131inter3));
  inv1  gate2357(.a(s_259), .O(gate131inter4));
  nand2 gate2358(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2359(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2360(.a(G414), .O(gate131inter7));
  inv1  gate2361(.a(G415), .O(gate131inter8));
  nand2 gate2362(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2363(.a(s_259), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2364(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2365(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2366(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1485(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1486(.a(gate132inter0), .b(s_134), .O(gate132inter1));
  and2  gate1487(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1488(.a(s_134), .O(gate132inter3));
  inv1  gate1489(.a(s_135), .O(gate132inter4));
  nand2 gate1490(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1491(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1492(.a(G416), .O(gate132inter7));
  inv1  gate1493(.a(G417), .O(gate132inter8));
  nand2 gate1494(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1495(.a(s_135), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1496(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1497(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1498(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1905(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1906(.a(gate136inter0), .b(s_194), .O(gate136inter1));
  and2  gate1907(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1908(.a(s_194), .O(gate136inter3));
  inv1  gate1909(.a(s_195), .O(gate136inter4));
  nand2 gate1910(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1911(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1912(.a(G424), .O(gate136inter7));
  inv1  gate1913(.a(G425), .O(gate136inter8));
  nand2 gate1914(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1915(.a(s_195), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1916(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1917(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1918(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2927(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2928(.a(gate137inter0), .b(s_340), .O(gate137inter1));
  and2  gate2929(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2930(.a(s_340), .O(gate137inter3));
  inv1  gate2931(.a(s_341), .O(gate137inter4));
  nand2 gate2932(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2933(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2934(.a(G426), .O(gate137inter7));
  inv1  gate2935(.a(G429), .O(gate137inter8));
  nand2 gate2936(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2937(.a(s_341), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2938(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2939(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2940(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate3123(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate3124(.a(gate139inter0), .b(s_368), .O(gate139inter1));
  and2  gate3125(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate3126(.a(s_368), .O(gate139inter3));
  inv1  gate3127(.a(s_369), .O(gate139inter4));
  nand2 gate3128(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate3129(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate3130(.a(G438), .O(gate139inter7));
  inv1  gate3131(.a(G441), .O(gate139inter8));
  nand2 gate3132(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate3133(.a(s_369), .b(gate139inter3), .O(gate139inter10));
  nor2  gate3134(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate3135(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate3136(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1275(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1276(.a(gate141inter0), .b(s_104), .O(gate141inter1));
  and2  gate1277(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1278(.a(s_104), .O(gate141inter3));
  inv1  gate1279(.a(s_105), .O(gate141inter4));
  nand2 gate1280(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1281(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1282(.a(G450), .O(gate141inter7));
  inv1  gate1283(.a(G453), .O(gate141inter8));
  nand2 gate1284(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1285(.a(s_105), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1286(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1287(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1288(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate2717(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2718(.a(gate142inter0), .b(s_310), .O(gate142inter1));
  and2  gate2719(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2720(.a(s_310), .O(gate142inter3));
  inv1  gate2721(.a(s_311), .O(gate142inter4));
  nand2 gate2722(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2723(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2724(.a(G456), .O(gate142inter7));
  inv1  gate2725(.a(G459), .O(gate142inter8));
  nand2 gate2726(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2727(.a(s_311), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2728(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2729(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2730(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate785(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate786(.a(gate143inter0), .b(s_34), .O(gate143inter1));
  and2  gate787(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate788(.a(s_34), .O(gate143inter3));
  inv1  gate789(.a(s_35), .O(gate143inter4));
  nand2 gate790(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate791(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate792(.a(G462), .O(gate143inter7));
  inv1  gate793(.a(G465), .O(gate143inter8));
  nand2 gate794(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate795(.a(s_35), .b(gate143inter3), .O(gate143inter10));
  nor2  gate796(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate797(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate798(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1933(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1934(.a(gate145inter0), .b(s_198), .O(gate145inter1));
  and2  gate1935(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1936(.a(s_198), .O(gate145inter3));
  inv1  gate1937(.a(s_199), .O(gate145inter4));
  nand2 gate1938(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1939(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1940(.a(G474), .O(gate145inter7));
  inv1  gate1941(.a(G477), .O(gate145inter8));
  nand2 gate1942(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1943(.a(s_199), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1944(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1945(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1946(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1849(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1850(.a(gate146inter0), .b(s_186), .O(gate146inter1));
  and2  gate1851(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1852(.a(s_186), .O(gate146inter3));
  inv1  gate1853(.a(s_187), .O(gate146inter4));
  nand2 gate1854(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1855(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1856(.a(G480), .O(gate146inter7));
  inv1  gate1857(.a(G483), .O(gate146inter8));
  nand2 gate1858(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1859(.a(s_187), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1860(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1861(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1862(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate757(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate758(.a(gate147inter0), .b(s_30), .O(gate147inter1));
  and2  gate759(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate760(.a(s_30), .O(gate147inter3));
  inv1  gate761(.a(s_31), .O(gate147inter4));
  nand2 gate762(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate763(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate764(.a(G486), .O(gate147inter7));
  inv1  gate765(.a(G489), .O(gate147inter8));
  nand2 gate766(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate767(.a(s_31), .b(gate147inter3), .O(gate147inter10));
  nor2  gate768(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate769(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate770(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1611(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1612(.a(gate149inter0), .b(s_152), .O(gate149inter1));
  and2  gate1613(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1614(.a(s_152), .O(gate149inter3));
  inv1  gate1615(.a(s_153), .O(gate149inter4));
  nand2 gate1616(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1617(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1618(.a(G498), .O(gate149inter7));
  inv1  gate1619(.a(G501), .O(gate149inter8));
  nand2 gate1620(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1621(.a(s_153), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1622(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1623(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1624(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2899(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2900(.a(gate151inter0), .b(s_336), .O(gate151inter1));
  and2  gate2901(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2902(.a(s_336), .O(gate151inter3));
  inv1  gate2903(.a(s_337), .O(gate151inter4));
  nand2 gate2904(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2905(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2906(.a(G510), .O(gate151inter7));
  inv1  gate2907(.a(G513), .O(gate151inter8));
  nand2 gate2908(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2909(.a(s_337), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2910(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2911(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2912(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1863(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1864(.a(gate153inter0), .b(s_188), .O(gate153inter1));
  and2  gate1865(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1866(.a(s_188), .O(gate153inter3));
  inv1  gate1867(.a(s_189), .O(gate153inter4));
  nand2 gate1868(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1869(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1870(.a(G426), .O(gate153inter7));
  inv1  gate1871(.a(G522), .O(gate153inter8));
  nand2 gate1872(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1873(.a(s_189), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1874(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1875(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1876(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2409(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2410(.a(gate154inter0), .b(s_266), .O(gate154inter1));
  and2  gate2411(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2412(.a(s_266), .O(gate154inter3));
  inv1  gate2413(.a(s_267), .O(gate154inter4));
  nand2 gate2414(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2415(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2416(.a(G429), .O(gate154inter7));
  inv1  gate2417(.a(G522), .O(gate154inter8));
  nand2 gate2418(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2419(.a(s_267), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2420(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2421(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2422(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1737(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1738(.a(gate155inter0), .b(s_170), .O(gate155inter1));
  and2  gate1739(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1740(.a(s_170), .O(gate155inter3));
  inv1  gate1741(.a(s_171), .O(gate155inter4));
  nand2 gate1742(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1743(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1744(.a(G432), .O(gate155inter7));
  inv1  gate1745(.a(G525), .O(gate155inter8));
  nand2 gate1746(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1747(.a(s_171), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1748(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1749(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1750(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2997(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2998(.a(gate156inter0), .b(s_350), .O(gate156inter1));
  and2  gate2999(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate3000(.a(s_350), .O(gate156inter3));
  inv1  gate3001(.a(s_351), .O(gate156inter4));
  nand2 gate3002(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate3003(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate3004(.a(G435), .O(gate156inter7));
  inv1  gate3005(.a(G525), .O(gate156inter8));
  nand2 gate3006(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate3007(.a(s_351), .b(gate156inter3), .O(gate156inter10));
  nor2  gate3008(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate3009(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate3010(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1807(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1808(.a(gate163inter0), .b(s_180), .O(gate163inter1));
  and2  gate1809(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1810(.a(s_180), .O(gate163inter3));
  inv1  gate1811(.a(s_181), .O(gate163inter4));
  nand2 gate1812(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1813(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1814(.a(G456), .O(gate163inter7));
  inv1  gate1815(.a(G537), .O(gate163inter8));
  nand2 gate1816(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1817(.a(s_181), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1818(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1819(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1820(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1303(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1304(.a(gate164inter0), .b(s_108), .O(gate164inter1));
  and2  gate1305(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1306(.a(s_108), .O(gate164inter3));
  inv1  gate1307(.a(s_109), .O(gate164inter4));
  nand2 gate1308(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1309(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1310(.a(G459), .O(gate164inter7));
  inv1  gate1311(.a(G537), .O(gate164inter8));
  nand2 gate1312(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1313(.a(s_109), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1314(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1315(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1316(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate2857(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2858(.a(gate165inter0), .b(s_330), .O(gate165inter1));
  and2  gate2859(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2860(.a(s_330), .O(gate165inter3));
  inv1  gate2861(.a(s_331), .O(gate165inter4));
  nand2 gate2862(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2863(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2864(.a(G462), .O(gate165inter7));
  inv1  gate2865(.a(G540), .O(gate165inter8));
  nand2 gate2866(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2867(.a(s_331), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2868(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2869(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2870(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate659(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate660(.a(gate166inter0), .b(s_16), .O(gate166inter1));
  and2  gate661(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate662(.a(s_16), .O(gate166inter3));
  inv1  gate663(.a(s_17), .O(gate166inter4));
  nand2 gate664(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate665(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate666(.a(G465), .O(gate166inter7));
  inv1  gate667(.a(G540), .O(gate166inter8));
  nand2 gate668(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate669(.a(s_17), .b(gate166inter3), .O(gate166inter10));
  nor2  gate670(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate671(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate672(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2591(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2592(.a(gate168inter0), .b(s_292), .O(gate168inter1));
  and2  gate2593(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2594(.a(s_292), .O(gate168inter3));
  inv1  gate2595(.a(s_293), .O(gate168inter4));
  nand2 gate2596(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2597(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2598(.a(G471), .O(gate168inter7));
  inv1  gate2599(.a(G543), .O(gate168inter8));
  nand2 gate2600(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2601(.a(s_293), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2602(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2603(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2604(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1065(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1066(.a(gate170inter0), .b(s_74), .O(gate170inter1));
  and2  gate1067(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1068(.a(s_74), .O(gate170inter3));
  inv1  gate1069(.a(s_75), .O(gate170inter4));
  nand2 gate1070(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1071(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1072(.a(G477), .O(gate170inter7));
  inv1  gate1073(.a(G546), .O(gate170inter8));
  nand2 gate1074(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1075(.a(s_75), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1076(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1077(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1078(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1961(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1962(.a(gate171inter0), .b(s_202), .O(gate171inter1));
  and2  gate1963(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1964(.a(s_202), .O(gate171inter3));
  inv1  gate1965(.a(s_203), .O(gate171inter4));
  nand2 gate1966(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1967(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1968(.a(G480), .O(gate171inter7));
  inv1  gate1969(.a(G549), .O(gate171inter8));
  nand2 gate1970(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1971(.a(s_203), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1972(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1973(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1974(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1359(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1360(.a(gate172inter0), .b(s_116), .O(gate172inter1));
  and2  gate1361(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1362(.a(s_116), .O(gate172inter3));
  inv1  gate1363(.a(s_117), .O(gate172inter4));
  nand2 gate1364(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1365(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1366(.a(G483), .O(gate172inter7));
  inv1  gate1367(.a(G549), .O(gate172inter8));
  nand2 gate1368(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1369(.a(s_117), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1370(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1371(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1372(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1205(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1206(.a(gate173inter0), .b(s_94), .O(gate173inter1));
  and2  gate1207(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1208(.a(s_94), .O(gate173inter3));
  inv1  gate1209(.a(s_95), .O(gate173inter4));
  nand2 gate1210(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1211(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1212(.a(G486), .O(gate173inter7));
  inv1  gate1213(.a(G552), .O(gate173inter8));
  nand2 gate1214(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1215(.a(s_95), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1216(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1217(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1218(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1471(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1472(.a(gate176inter0), .b(s_132), .O(gate176inter1));
  and2  gate1473(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1474(.a(s_132), .O(gate176inter3));
  inv1  gate1475(.a(s_133), .O(gate176inter4));
  nand2 gate1476(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1477(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1478(.a(G495), .O(gate176inter7));
  inv1  gate1479(.a(G555), .O(gate176inter8));
  nand2 gate1480(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1481(.a(s_133), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1482(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1483(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1484(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1149(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1150(.a(gate180inter0), .b(s_86), .O(gate180inter1));
  and2  gate1151(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1152(.a(s_86), .O(gate180inter3));
  inv1  gate1153(.a(s_87), .O(gate180inter4));
  nand2 gate1154(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1155(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1156(.a(G507), .O(gate180inter7));
  inv1  gate1157(.a(G561), .O(gate180inter8));
  nand2 gate1158(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1159(.a(s_87), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1160(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1161(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1162(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate771(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate772(.a(gate181inter0), .b(s_32), .O(gate181inter1));
  and2  gate773(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate774(.a(s_32), .O(gate181inter3));
  inv1  gate775(.a(s_33), .O(gate181inter4));
  nand2 gate776(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate777(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate778(.a(G510), .O(gate181inter7));
  inv1  gate779(.a(G564), .O(gate181inter8));
  nand2 gate780(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate781(.a(s_33), .b(gate181inter3), .O(gate181inter10));
  nor2  gate782(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate783(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate784(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1373(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1374(.a(gate184inter0), .b(s_118), .O(gate184inter1));
  and2  gate1375(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1376(.a(s_118), .O(gate184inter3));
  inv1  gate1377(.a(s_119), .O(gate184inter4));
  nand2 gate1378(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1379(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1380(.a(G519), .O(gate184inter7));
  inv1  gate1381(.a(G567), .O(gate184inter8));
  nand2 gate1382(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1383(.a(s_119), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1384(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1385(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1386(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2955(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2956(.a(gate185inter0), .b(s_344), .O(gate185inter1));
  and2  gate2957(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2958(.a(s_344), .O(gate185inter3));
  inv1  gate2959(.a(s_345), .O(gate185inter4));
  nand2 gate2960(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2961(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2962(.a(G570), .O(gate185inter7));
  inv1  gate2963(.a(G571), .O(gate185inter8));
  nand2 gate2964(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2965(.a(s_345), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2966(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2967(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2968(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate3081(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate3082(.a(gate186inter0), .b(s_362), .O(gate186inter1));
  and2  gate3083(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate3084(.a(s_362), .O(gate186inter3));
  inv1  gate3085(.a(s_363), .O(gate186inter4));
  nand2 gate3086(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate3087(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate3088(.a(G572), .O(gate186inter7));
  inv1  gate3089(.a(G573), .O(gate186inter8));
  nand2 gate3090(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate3091(.a(s_363), .b(gate186inter3), .O(gate186inter10));
  nor2  gate3092(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate3093(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate3094(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1555(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1556(.a(gate188inter0), .b(s_144), .O(gate188inter1));
  and2  gate1557(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1558(.a(s_144), .O(gate188inter3));
  inv1  gate1559(.a(s_145), .O(gate188inter4));
  nand2 gate1560(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1561(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1562(.a(G576), .O(gate188inter7));
  inv1  gate1563(.a(G577), .O(gate188inter8));
  nand2 gate1564(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1565(.a(s_145), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1566(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1567(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1568(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate2787(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2788(.a(gate192inter0), .b(s_320), .O(gate192inter1));
  and2  gate2789(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2790(.a(s_320), .O(gate192inter3));
  inv1  gate2791(.a(s_321), .O(gate192inter4));
  nand2 gate2792(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2793(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2794(.a(G584), .O(gate192inter7));
  inv1  gate2795(.a(G585), .O(gate192inter8));
  nand2 gate2796(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2797(.a(s_321), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2798(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2799(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2800(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1765(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1766(.a(gate193inter0), .b(s_174), .O(gate193inter1));
  and2  gate1767(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1768(.a(s_174), .O(gate193inter3));
  inv1  gate1769(.a(s_175), .O(gate193inter4));
  nand2 gate1770(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1771(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1772(.a(G586), .O(gate193inter7));
  inv1  gate1773(.a(G587), .O(gate193inter8));
  nand2 gate1774(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1775(.a(s_175), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1776(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1777(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1778(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1135(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1136(.a(gate195inter0), .b(s_84), .O(gate195inter1));
  and2  gate1137(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1138(.a(s_84), .O(gate195inter3));
  inv1  gate1139(.a(s_85), .O(gate195inter4));
  nand2 gate1140(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1141(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1142(.a(G590), .O(gate195inter7));
  inv1  gate1143(.a(G591), .O(gate195inter8));
  nand2 gate1144(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1145(.a(s_85), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1146(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1147(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1148(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate3179(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate3180(.a(gate197inter0), .b(s_376), .O(gate197inter1));
  and2  gate3181(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate3182(.a(s_376), .O(gate197inter3));
  inv1  gate3183(.a(s_377), .O(gate197inter4));
  nand2 gate3184(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate3185(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate3186(.a(G594), .O(gate197inter7));
  inv1  gate3187(.a(G595), .O(gate197inter8));
  nand2 gate3188(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate3189(.a(s_377), .b(gate197inter3), .O(gate197inter10));
  nor2  gate3190(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate3191(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate3192(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate3039(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate3040(.a(gate201inter0), .b(s_356), .O(gate201inter1));
  and2  gate3041(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate3042(.a(s_356), .O(gate201inter3));
  inv1  gate3043(.a(s_357), .O(gate201inter4));
  nand2 gate3044(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate3045(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate3046(.a(G602), .O(gate201inter7));
  inv1  gate3047(.a(G607), .O(gate201inter8));
  nand2 gate3048(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate3049(.a(s_357), .b(gate201inter3), .O(gate201inter10));
  nor2  gate3050(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate3051(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate3052(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate897(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate898(.a(gate206inter0), .b(s_50), .O(gate206inter1));
  and2  gate899(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate900(.a(s_50), .O(gate206inter3));
  inv1  gate901(.a(s_51), .O(gate206inter4));
  nand2 gate902(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate903(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate904(.a(G632), .O(gate206inter7));
  inv1  gate905(.a(G637), .O(gate206inter8));
  nand2 gate906(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate907(.a(s_51), .b(gate206inter3), .O(gate206inter10));
  nor2  gate908(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate909(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate910(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1387(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1388(.a(gate209inter0), .b(s_120), .O(gate209inter1));
  and2  gate1389(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1390(.a(s_120), .O(gate209inter3));
  inv1  gate1391(.a(s_121), .O(gate209inter4));
  nand2 gate1392(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1393(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1394(.a(G602), .O(gate209inter7));
  inv1  gate1395(.a(G666), .O(gate209inter8));
  nand2 gate1396(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1397(.a(s_121), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1398(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1399(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1400(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1779(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1780(.a(gate210inter0), .b(s_176), .O(gate210inter1));
  and2  gate1781(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1782(.a(s_176), .O(gate210inter3));
  inv1  gate1783(.a(s_177), .O(gate210inter4));
  nand2 gate1784(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1785(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1786(.a(G607), .O(gate210inter7));
  inv1  gate1787(.a(G666), .O(gate210inter8));
  nand2 gate1788(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1789(.a(s_177), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1790(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1791(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1792(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate701(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate702(.a(gate212inter0), .b(s_22), .O(gate212inter1));
  and2  gate703(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate704(.a(s_22), .O(gate212inter3));
  inv1  gate705(.a(s_23), .O(gate212inter4));
  nand2 gate706(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate707(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate708(.a(G617), .O(gate212inter7));
  inv1  gate709(.a(G669), .O(gate212inter8));
  nand2 gate710(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate711(.a(s_23), .b(gate212inter3), .O(gate212inter10));
  nor2  gate712(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate713(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate714(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1751(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1752(.a(gate213inter0), .b(s_172), .O(gate213inter1));
  and2  gate1753(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1754(.a(s_172), .O(gate213inter3));
  inv1  gate1755(.a(s_173), .O(gate213inter4));
  nand2 gate1756(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1757(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1758(.a(G602), .O(gate213inter7));
  inv1  gate1759(.a(G672), .O(gate213inter8));
  nand2 gate1760(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1761(.a(s_173), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1762(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1763(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1764(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1023(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1024(.a(gate214inter0), .b(s_68), .O(gate214inter1));
  and2  gate1025(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1026(.a(s_68), .O(gate214inter3));
  inv1  gate1027(.a(s_69), .O(gate214inter4));
  nand2 gate1028(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1029(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1030(.a(G612), .O(gate214inter7));
  inv1  gate1031(.a(G672), .O(gate214inter8));
  nand2 gate1032(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1033(.a(s_69), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1034(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1035(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1036(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1709(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1710(.a(gate215inter0), .b(s_166), .O(gate215inter1));
  and2  gate1711(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1712(.a(s_166), .O(gate215inter3));
  inv1  gate1713(.a(s_167), .O(gate215inter4));
  nand2 gate1714(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1715(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1716(.a(G607), .O(gate215inter7));
  inv1  gate1717(.a(G675), .O(gate215inter8));
  nand2 gate1718(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1719(.a(s_167), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1720(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1721(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1722(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1975(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1976(.a(gate216inter0), .b(s_204), .O(gate216inter1));
  and2  gate1977(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1978(.a(s_204), .O(gate216inter3));
  inv1  gate1979(.a(s_205), .O(gate216inter4));
  nand2 gate1980(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1981(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1982(.a(G617), .O(gate216inter7));
  inv1  gate1983(.a(G675), .O(gate216inter8));
  nand2 gate1984(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1985(.a(s_205), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1986(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1987(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1988(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2689(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2690(.a(gate220inter0), .b(s_306), .O(gate220inter1));
  and2  gate2691(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2692(.a(s_306), .O(gate220inter3));
  inv1  gate2693(.a(s_307), .O(gate220inter4));
  nand2 gate2694(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2695(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2696(.a(G637), .O(gate220inter7));
  inv1  gate2697(.a(G681), .O(gate220inter8));
  nand2 gate2698(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2699(.a(s_307), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2700(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2701(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2702(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1331(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1332(.a(gate221inter0), .b(s_112), .O(gate221inter1));
  and2  gate1333(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1334(.a(s_112), .O(gate221inter3));
  inv1  gate1335(.a(s_113), .O(gate221inter4));
  nand2 gate1336(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1337(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1338(.a(G622), .O(gate221inter7));
  inv1  gate1339(.a(G684), .O(gate221inter8));
  nand2 gate1340(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1341(.a(s_113), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1342(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1343(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1344(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate687(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate688(.a(gate225inter0), .b(s_20), .O(gate225inter1));
  and2  gate689(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate690(.a(s_20), .O(gate225inter3));
  inv1  gate691(.a(s_21), .O(gate225inter4));
  nand2 gate692(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate693(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate694(.a(G690), .O(gate225inter7));
  inv1  gate695(.a(G691), .O(gate225inter8));
  nand2 gate696(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate697(.a(s_21), .b(gate225inter3), .O(gate225inter10));
  nor2  gate698(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate699(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate700(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate729(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate730(.a(gate226inter0), .b(s_26), .O(gate226inter1));
  and2  gate731(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate732(.a(s_26), .O(gate226inter3));
  inv1  gate733(.a(s_27), .O(gate226inter4));
  nand2 gate734(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate735(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate736(.a(G692), .O(gate226inter7));
  inv1  gate737(.a(G693), .O(gate226inter8));
  nand2 gate738(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate739(.a(s_27), .b(gate226inter3), .O(gate226inter10));
  nor2  gate740(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate741(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate742(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2815(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2816(.a(gate229inter0), .b(s_324), .O(gate229inter1));
  and2  gate2817(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2818(.a(s_324), .O(gate229inter3));
  inv1  gate2819(.a(s_325), .O(gate229inter4));
  nand2 gate2820(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2821(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2822(.a(G698), .O(gate229inter7));
  inv1  gate2823(.a(G699), .O(gate229inter8));
  nand2 gate2824(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2825(.a(s_325), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2826(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2827(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2828(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1191(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1192(.a(gate233inter0), .b(s_92), .O(gate233inter1));
  and2  gate1193(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1194(.a(s_92), .O(gate233inter3));
  inv1  gate1195(.a(s_93), .O(gate233inter4));
  nand2 gate1196(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1197(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1198(.a(G242), .O(gate233inter7));
  inv1  gate1199(.a(G718), .O(gate233inter8));
  nand2 gate1200(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1201(.a(s_93), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1202(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1203(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1204(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate3067(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate3068(.a(gate234inter0), .b(s_360), .O(gate234inter1));
  and2  gate3069(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate3070(.a(s_360), .O(gate234inter3));
  inv1  gate3071(.a(s_361), .O(gate234inter4));
  nand2 gate3072(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate3073(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate3074(.a(G245), .O(gate234inter7));
  inv1  gate3075(.a(G721), .O(gate234inter8));
  nand2 gate3076(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate3077(.a(s_361), .b(gate234inter3), .O(gate234inter10));
  nor2  gate3078(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate3079(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate3080(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2619(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2620(.a(gate235inter0), .b(s_296), .O(gate235inter1));
  and2  gate2621(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2622(.a(s_296), .O(gate235inter3));
  inv1  gate2623(.a(s_297), .O(gate235inter4));
  nand2 gate2624(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2625(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2626(.a(G248), .O(gate235inter7));
  inv1  gate2627(.a(G724), .O(gate235inter8));
  nand2 gate2628(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2629(.a(s_297), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2630(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2631(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2632(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2913(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2914(.a(gate240inter0), .b(s_338), .O(gate240inter1));
  and2  gate2915(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2916(.a(s_338), .O(gate240inter3));
  inv1  gate2917(.a(s_339), .O(gate240inter4));
  nand2 gate2918(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2919(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2920(.a(G263), .O(gate240inter7));
  inv1  gate2921(.a(G715), .O(gate240inter8));
  nand2 gate2922(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2923(.a(s_339), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2924(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2925(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2926(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate2199(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2200(.a(gate241inter0), .b(s_236), .O(gate241inter1));
  and2  gate2201(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2202(.a(s_236), .O(gate241inter3));
  inv1  gate2203(.a(s_237), .O(gate241inter4));
  nand2 gate2204(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2205(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2206(.a(G242), .O(gate241inter7));
  inv1  gate2207(.a(G730), .O(gate241inter8));
  nand2 gate2208(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2209(.a(s_237), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2210(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2211(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2212(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1443(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1444(.a(gate251inter0), .b(s_128), .O(gate251inter1));
  and2  gate1445(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1446(.a(s_128), .O(gate251inter3));
  inv1  gate1447(.a(s_129), .O(gate251inter4));
  nand2 gate1448(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1449(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1450(.a(G257), .O(gate251inter7));
  inv1  gate1451(.a(G745), .O(gate251inter8));
  nand2 gate1452(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1453(.a(s_129), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1454(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1455(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1456(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2647(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2648(.a(gate255inter0), .b(s_300), .O(gate255inter1));
  and2  gate2649(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2650(.a(s_300), .O(gate255inter3));
  inv1  gate2651(.a(s_301), .O(gate255inter4));
  nand2 gate2652(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2653(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2654(.a(G263), .O(gate255inter7));
  inv1  gate2655(.a(G751), .O(gate255inter8));
  nand2 gate2656(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2657(.a(s_301), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2658(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2659(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2660(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1947(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1948(.a(gate256inter0), .b(s_200), .O(gate256inter1));
  and2  gate1949(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1950(.a(s_200), .O(gate256inter3));
  inv1  gate1951(.a(s_201), .O(gate256inter4));
  nand2 gate1952(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1953(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1954(.a(G715), .O(gate256inter7));
  inv1  gate1955(.a(G751), .O(gate256inter8));
  nand2 gate1956(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1957(.a(s_201), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1958(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1959(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1960(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate2437(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2438(.a(gate260inter0), .b(s_270), .O(gate260inter1));
  and2  gate2439(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2440(.a(s_270), .O(gate260inter3));
  inv1  gate2441(.a(s_271), .O(gate260inter4));
  nand2 gate2442(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2443(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2444(.a(G760), .O(gate260inter7));
  inv1  gate2445(.a(G761), .O(gate260inter8));
  nand2 gate2446(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2447(.a(s_271), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2448(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2449(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2450(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1009(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1010(.a(gate262inter0), .b(s_66), .O(gate262inter1));
  and2  gate1011(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1012(.a(s_66), .O(gate262inter3));
  inv1  gate1013(.a(s_67), .O(gate262inter4));
  nand2 gate1014(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1015(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1016(.a(G764), .O(gate262inter7));
  inv1  gate1017(.a(G765), .O(gate262inter8));
  nand2 gate1018(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1019(.a(s_67), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1020(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1021(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1022(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2213(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2214(.a(gate263inter0), .b(s_238), .O(gate263inter1));
  and2  gate2215(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2216(.a(s_238), .O(gate263inter3));
  inv1  gate2217(.a(s_239), .O(gate263inter4));
  nand2 gate2218(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2219(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2220(.a(G766), .O(gate263inter7));
  inv1  gate2221(.a(G767), .O(gate263inter8));
  nand2 gate2222(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2223(.a(s_239), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2224(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2225(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2226(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2731(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2732(.a(gate264inter0), .b(s_312), .O(gate264inter1));
  and2  gate2733(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2734(.a(s_312), .O(gate264inter3));
  inv1  gate2735(.a(s_313), .O(gate264inter4));
  nand2 gate2736(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2737(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2738(.a(G768), .O(gate264inter7));
  inv1  gate2739(.a(G769), .O(gate264inter8));
  nand2 gate2740(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2741(.a(s_313), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2742(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2743(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2744(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate3165(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate3166(.a(gate266inter0), .b(s_374), .O(gate266inter1));
  and2  gate3167(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate3168(.a(s_374), .O(gate266inter3));
  inv1  gate3169(.a(s_375), .O(gate266inter4));
  nand2 gate3170(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate3171(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate3172(.a(G645), .O(gate266inter7));
  inv1  gate3173(.a(G773), .O(gate266inter8));
  nand2 gate3174(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate3175(.a(s_375), .b(gate266inter3), .O(gate266inter10));
  nor2  gate3176(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate3177(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate3178(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2255(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2256(.a(gate268inter0), .b(s_244), .O(gate268inter1));
  and2  gate2257(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2258(.a(s_244), .O(gate268inter3));
  inv1  gate2259(.a(s_245), .O(gate268inter4));
  nand2 gate2260(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2261(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2262(.a(G651), .O(gate268inter7));
  inv1  gate2263(.a(G779), .O(gate268inter8));
  nand2 gate2264(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2265(.a(s_245), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2266(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2267(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2268(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2605(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2606(.a(gate270inter0), .b(s_294), .O(gate270inter1));
  and2  gate2607(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2608(.a(s_294), .O(gate270inter3));
  inv1  gate2609(.a(s_295), .O(gate270inter4));
  nand2 gate2610(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2611(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2612(.a(G657), .O(gate270inter7));
  inv1  gate2613(.a(G785), .O(gate270inter8));
  nand2 gate2614(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2615(.a(s_295), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2616(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2617(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2618(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1289(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1290(.a(gate271inter0), .b(s_106), .O(gate271inter1));
  and2  gate1291(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1292(.a(s_106), .O(gate271inter3));
  inv1  gate1293(.a(s_107), .O(gate271inter4));
  nand2 gate1294(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1295(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1296(.a(G660), .O(gate271inter7));
  inv1  gate1297(.a(G788), .O(gate271inter8));
  nand2 gate1298(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1299(.a(s_107), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1300(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1301(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1302(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2423(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2424(.a(gate272inter0), .b(s_268), .O(gate272inter1));
  and2  gate2425(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2426(.a(s_268), .O(gate272inter3));
  inv1  gate2427(.a(s_269), .O(gate272inter4));
  nand2 gate2428(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2429(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2430(.a(G663), .O(gate272inter7));
  inv1  gate2431(.a(G791), .O(gate272inter8));
  nand2 gate2432(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2433(.a(s_269), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2434(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2435(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2436(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate631(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate632(.a(gate276inter0), .b(s_12), .O(gate276inter1));
  and2  gate633(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate634(.a(s_12), .O(gate276inter3));
  inv1  gate635(.a(s_13), .O(gate276inter4));
  nand2 gate636(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate637(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate638(.a(G773), .O(gate276inter7));
  inv1  gate639(.a(G797), .O(gate276inter8));
  nand2 gate640(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate641(.a(s_13), .b(gate276inter3), .O(gate276inter10));
  nor2  gate642(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate643(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate644(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1499(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1500(.a(gate279inter0), .b(s_136), .O(gate279inter1));
  and2  gate1501(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1502(.a(s_136), .O(gate279inter3));
  inv1  gate1503(.a(s_137), .O(gate279inter4));
  nand2 gate1504(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1505(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1506(.a(G651), .O(gate279inter7));
  inv1  gate1507(.a(G803), .O(gate279inter8));
  nand2 gate1508(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1509(.a(s_137), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1510(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1511(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1512(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1093(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1094(.a(gate283inter0), .b(s_78), .O(gate283inter1));
  and2  gate1095(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1096(.a(s_78), .O(gate283inter3));
  inv1  gate1097(.a(s_79), .O(gate283inter4));
  nand2 gate1098(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1099(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1100(.a(G657), .O(gate283inter7));
  inv1  gate1101(.a(G809), .O(gate283inter8));
  nand2 gate1102(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1103(.a(s_79), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1104(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1105(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1106(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate2395(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2396(.a(gate284inter0), .b(s_264), .O(gate284inter1));
  and2  gate2397(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2398(.a(s_264), .O(gate284inter3));
  inv1  gate2399(.a(s_265), .O(gate284inter4));
  nand2 gate2400(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2401(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2402(.a(G785), .O(gate284inter7));
  inv1  gate2403(.a(G809), .O(gate284inter8));
  nand2 gate2404(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2405(.a(s_265), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2406(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2407(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2408(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1177(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1178(.a(gate287inter0), .b(s_90), .O(gate287inter1));
  and2  gate1179(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1180(.a(s_90), .O(gate287inter3));
  inv1  gate1181(.a(s_91), .O(gate287inter4));
  nand2 gate1182(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1183(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1184(.a(G663), .O(gate287inter7));
  inv1  gate1185(.a(G815), .O(gate287inter8));
  nand2 gate1186(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1187(.a(s_91), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1188(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1189(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1190(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate575(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate576(.a(gate288inter0), .b(s_4), .O(gate288inter1));
  and2  gate577(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate578(.a(s_4), .O(gate288inter3));
  inv1  gate579(.a(s_5), .O(gate288inter4));
  nand2 gate580(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate581(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate582(.a(G791), .O(gate288inter7));
  inv1  gate583(.a(G815), .O(gate288inter8));
  nand2 gate584(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate585(.a(s_5), .b(gate288inter3), .O(gate288inter10));
  nor2  gate586(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate587(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate588(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1527(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1528(.a(gate289inter0), .b(s_140), .O(gate289inter1));
  and2  gate1529(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1530(.a(s_140), .O(gate289inter3));
  inv1  gate1531(.a(s_141), .O(gate289inter4));
  nand2 gate1532(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1533(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1534(.a(G818), .O(gate289inter7));
  inv1  gate1535(.a(G819), .O(gate289inter8));
  nand2 gate1536(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1537(.a(s_141), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1538(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1539(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1540(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate3053(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate3054(.a(gate291inter0), .b(s_358), .O(gate291inter1));
  and2  gate3055(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate3056(.a(s_358), .O(gate291inter3));
  inv1  gate3057(.a(s_359), .O(gate291inter4));
  nand2 gate3058(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate3059(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate3060(.a(G822), .O(gate291inter7));
  inv1  gate3061(.a(G823), .O(gate291inter8));
  nand2 gate3062(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate3063(.a(s_359), .b(gate291inter3), .O(gate291inter10));
  nor2  gate3064(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate3065(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate3066(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate869(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate870(.a(gate293inter0), .b(s_46), .O(gate293inter1));
  and2  gate871(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate872(.a(s_46), .O(gate293inter3));
  inv1  gate873(.a(s_47), .O(gate293inter4));
  nand2 gate874(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate875(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate876(.a(G828), .O(gate293inter7));
  inv1  gate877(.a(G829), .O(gate293inter8));
  nand2 gate878(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate879(.a(s_47), .b(gate293inter3), .O(gate293inter10));
  nor2  gate880(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate881(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate882(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2311(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2312(.a(gate295inter0), .b(s_252), .O(gate295inter1));
  and2  gate2313(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2314(.a(s_252), .O(gate295inter3));
  inv1  gate2315(.a(s_253), .O(gate295inter4));
  nand2 gate2316(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2317(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2318(.a(G830), .O(gate295inter7));
  inv1  gate2319(.a(G831), .O(gate295inter8));
  nand2 gate2320(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2321(.a(s_253), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2322(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2323(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2324(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate2801(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2802(.a(gate296inter0), .b(s_322), .O(gate296inter1));
  and2  gate2803(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2804(.a(s_322), .O(gate296inter3));
  inv1  gate2805(.a(s_323), .O(gate296inter4));
  nand2 gate2806(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2807(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2808(.a(G826), .O(gate296inter7));
  inv1  gate2809(.a(G827), .O(gate296inter8));
  nand2 gate2810(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2811(.a(s_323), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2812(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2813(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2814(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2269(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2270(.a(gate388inter0), .b(s_246), .O(gate388inter1));
  and2  gate2271(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2272(.a(s_246), .O(gate388inter3));
  inv1  gate2273(.a(s_247), .O(gate388inter4));
  nand2 gate2274(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2275(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2276(.a(G2), .O(gate388inter7));
  inv1  gate2277(.a(G1039), .O(gate388inter8));
  nand2 gate2278(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2279(.a(s_247), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2280(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2281(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2282(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate3109(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate3110(.a(gate389inter0), .b(s_366), .O(gate389inter1));
  and2  gate3111(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate3112(.a(s_366), .O(gate389inter3));
  inv1  gate3113(.a(s_367), .O(gate389inter4));
  nand2 gate3114(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate3115(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate3116(.a(G3), .O(gate389inter7));
  inv1  gate3117(.a(G1042), .O(gate389inter8));
  nand2 gate3118(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate3119(.a(s_367), .b(gate389inter3), .O(gate389inter10));
  nor2  gate3120(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate3121(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate3122(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate925(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate926(.a(gate390inter0), .b(s_54), .O(gate390inter1));
  and2  gate927(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate928(.a(s_54), .O(gate390inter3));
  inv1  gate929(.a(s_55), .O(gate390inter4));
  nand2 gate930(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate931(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate932(.a(G4), .O(gate390inter7));
  inv1  gate933(.a(G1045), .O(gate390inter8));
  nand2 gate934(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate935(.a(s_55), .b(gate390inter3), .O(gate390inter10));
  nor2  gate936(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate937(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate938(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2829(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2830(.a(gate392inter0), .b(s_326), .O(gate392inter1));
  and2  gate2831(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2832(.a(s_326), .O(gate392inter3));
  inv1  gate2833(.a(s_327), .O(gate392inter4));
  nand2 gate2834(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2835(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2836(.a(G6), .O(gate392inter7));
  inv1  gate2837(.a(G1051), .O(gate392inter8));
  nand2 gate2838(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2839(.a(s_327), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2840(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2841(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2842(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2157(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2158(.a(gate395inter0), .b(s_230), .O(gate395inter1));
  and2  gate2159(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2160(.a(s_230), .O(gate395inter3));
  inv1  gate2161(.a(s_231), .O(gate395inter4));
  nand2 gate2162(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2163(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2164(.a(G9), .O(gate395inter7));
  inv1  gate2165(.a(G1060), .O(gate395inter8));
  nand2 gate2166(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2167(.a(s_231), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2168(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2169(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2170(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate3207(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate3208(.a(gate397inter0), .b(s_380), .O(gate397inter1));
  and2  gate3209(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate3210(.a(s_380), .O(gate397inter3));
  inv1  gate3211(.a(s_381), .O(gate397inter4));
  nand2 gate3212(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate3213(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate3214(.a(G11), .O(gate397inter7));
  inv1  gate3215(.a(G1066), .O(gate397inter8));
  nand2 gate3216(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate3217(.a(s_381), .b(gate397inter3), .O(gate397inter10));
  nor2  gate3218(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate3219(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate3220(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1163(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1164(.a(gate398inter0), .b(s_88), .O(gate398inter1));
  and2  gate1165(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1166(.a(s_88), .O(gate398inter3));
  inv1  gate1167(.a(s_89), .O(gate398inter4));
  nand2 gate1168(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1169(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1170(.a(G12), .O(gate398inter7));
  inv1  gate1171(.a(G1069), .O(gate398inter8));
  nand2 gate1172(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1173(.a(s_89), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1174(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1175(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1176(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1233(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1234(.a(gate400inter0), .b(s_98), .O(gate400inter1));
  and2  gate1235(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1236(.a(s_98), .O(gate400inter3));
  inv1  gate1237(.a(s_99), .O(gate400inter4));
  nand2 gate1238(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1239(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1240(.a(G14), .O(gate400inter7));
  inv1  gate1241(.a(G1075), .O(gate400inter8));
  nand2 gate1242(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1243(.a(s_99), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1244(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1245(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1246(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2479(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2480(.a(gate404inter0), .b(s_276), .O(gate404inter1));
  and2  gate2481(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2482(.a(s_276), .O(gate404inter3));
  inv1  gate2483(.a(s_277), .O(gate404inter4));
  nand2 gate2484(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2485(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2486(.a(G18), .O(gate404inter7));
  inv1  gate2487(.a(G1087), .O(gate404inter8));
  nand2 gate2488(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2489(.a(s_277), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2490(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2491(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2492(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate911(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate912(.a(gate406inter0), .b(s_52), .O(gate406inter1));
  and2  gate913(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate914(.a(s_52), .O(gate406inter3));
  inv1  gate915(.a(s_53), .O(gate406inter4));
  nand2 gate916(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate917(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate918(.a(G20), .O(gate406inter7));
  inv1  gate919(.a(G1093), .O(gate406inter8));
  nand2 gate920(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate921(.a(s_53), .b(gate406inter3), .O(gate406inter10));
  nor2  gate922(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate923(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate924(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2633(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2634(.a(gate410inter0), .b(s_298), .O(gate410inter1));
  and2  gate2635(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2636(.a(s_298), .O(gate410inter3));
  inv1  gate2637(.a(s_299), .O(gate410inter4));
  nand2 gate2638(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2639(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2640(.a(G24), .O(gate410inter7));
  inv1  gate2641(.a(G1105), .O(gate410inter8));
  nand2 gate2642(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2643(.a(s_299), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2644(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2645(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2646(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate3095(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate3096(.a(gate411inter0), .b(s_364), .O(gate411inter1));
  and2  gate3097(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate3098(.a(s_364), .O(gate411inter3));
  inv1  gate3099(.a(s_365), .O(gate411inter4));
  nand2 gate3100(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate3101(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate3102(.a(G25), .O(gate411inter7));
  inv1  gate3103(.a(G1108), .O(gate411inter8));
  nand2 gate3104(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate3105(.a(s_365), .b(gate411inter3), .O(gate411inter10));
  nor2  gate3106(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate3107(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate3108(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2843(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2844(.a(gate412inter0), .b(s_328), .O(gate412inter1));
  and2  gate2845(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2846(.a(s_328), .O(gate412inter3));
  inv1  gate2847(.a(s_329), .O(gate412inter4));
  nand2 gate2848(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2849(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2850(.a(G26), .O(gate412inter7));
  inv1  gate2851(.a(G1111), .O(gate412inter8));
  nand2 gate2852(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2853(.a(s_329), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2854(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2855(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2856(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate2003(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2004(.a(gate413inter0), .b(s_208), .O(gate413inter1));
  and2  gate2005(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2006(.a(s_208), .O(gate413inter3));
  inv1  gate2007(.a(s_209), .O(gate413inter4));
  nand2 gate2008(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2009(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2010(.a(G27), .O(gate413inter7));
  inv1  gate2011(.a(G1114), .O(gate413inter8));
  nand2 gate2012(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2013(.a(s_209), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2014(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2015(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2016(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate715(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate716(.a(gate416inter0), .b(s_24), .O(gate416inter1));
  and2  gate717(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate718(.a(s_24), .O(gate416inter3));
  inv1  gate719(.a(s_25), .O(gate416inter4));
  nand2 gate720(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate721(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate722(.a(G30), .O(gate416inter7));
  inv1  gate723(.a(G1123), .O(gate416inter8));
  nand2 gate724(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate725(.a(s_25), .b(gate416inter3), .O(gate416inter10));
  nor2  gate726(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate727(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate728(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2367(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2368(.a(gate418inter0), .b(s_260), .O(gate418inter1));
  and2  gate2369(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2370(.a(s_260), .O(gate418inter3));
  inv1  gate2371(.a(s_261), .O(gate418inter4));
  nand2 gate2372(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2373(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2374(.a(G32), .O(gate418inter7));
  inv1  gate2375(.a(G1129), .O(gate418inter8));
  nand2 gate2376(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2377(.a(s_261), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2378(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2379(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2380(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2535(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2536(.a(gate421inter0), .b(s_284), .O(gate421inter1));
  and2  gate2537(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2538(.a(s_284), .O(gate421inter3));
  inv1  gate2539(.a(s_285), .O(gate421inter4));
  nand2 gate2540(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2541(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2542(.a(G2), .O(gate421inter7));
  inv1  gate2543(.a(G1135), .O(gate421inter8));
  nand2 gate2544(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2545(.a(s_285), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2546(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2547(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2548(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2983(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2984(.a(gate423inter0), .b(s_348), .O(gate423inter1));
  and2  gate2985(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2986(.a(s_348), .O(gate423inter3));
  inv1  gate2987(.a(s_349), .O(gate423inter4));
  nand2 gate2988(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2989(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2990(.a(G3), .O(gate423inter7));
  inv1  gate2991(.a(G1138), .O(gate423inter8));
  nand2 gate2992(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2993(.a(s_349), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2994(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2995(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2996(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate967(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate968(.a(gate424inter0), .b(s_60), .O(gate424inter1));
  and2  gate969(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate970(.a(s_60), .O(gate424inter3));
  inv1  gate971(.a(s_61), .O(gate424inter4));
  nand2 gate972(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate973(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate974(.a(G1042), .O(gate424inter7));
  inv1  gate975(.a(G1138), .O(gate424inter8));
  nand2 gate976(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate977(.a(s_61), .b(gate424inter3), .O(gate424inter10));
  nor2  gate978(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate979(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate980(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate2465(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2466(.a(gate427inter0), .b(s_274), .O(gate427inter1));
  and2  gate2467(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2468(.a(s_274), .O(gate427inter3));
  inv1  gate2469(.a(s_275), .O(gate427inter4));
  nand2 gate2470(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2471(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2472(.a(G5), .O(gate427inter7));
  inv1  gate2473(.a(G1144), .O(gate427inter8));
  nand2 gate2474(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2475(.a(s_275), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2476(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2477(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2478(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate547(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate548(.a(gate430inter0), .b(s_0), .O(gate430inter1));
  and2  gate549(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate550(.a(s_0), .O(gate430inter3));
  inv1  gate551(.a(s_1), .O(gate430inter4));
  nand2 gate552(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate553(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate554(.a(G1051), .O(gate430inter7));
  inv1  gate555(.a(G1147), .O(gate430inter8));
  nand2 gate556(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate557(.a(s_1), .b(gate430inter3), .O(gate430inter10));
  nor2  gate558(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate559(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate560(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2031(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2032(.a(gate431inter0), .b(s_212), .O(gate431inter1));
  and2  gate2033(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2034(.a(s_212), .O(gate431inter3));
  inv1  gate2035(.a(s_213), .O(gate431inter4));
  nand2 gate2036(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2037(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2038(.a(G7), .O(gate431inter7));
  inv1  gate2039(.a(G1150), .O(gate431inter8));
  nand2 gate2040(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2041(.a(s_213), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2042(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2043(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2044(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2059(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2060(.a(gate432inter0), .b(s_216), .O(gate432inter1));
  and2  gate2061(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2062(.a(s_216), .O(gate432inter3));
  inv1  gate2063(.a(s_217), .O(gate432inter4));
  nand2 gate2064(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2065(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2066(.a(G1054), .O(gate432inter7));
  inv1  gate2067(.a(G1150), .O(gate432inter8));
  nand2 gate2068(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2069(.a(s_217), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2070(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2071(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2072(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2115(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2116(.a(gate434inter0), .b(s_224), .O(gate434inter1));
  and2  gate2117(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2118(.a(s_224), .O(gate434inter3));
  inv1  gate2119(.a(s_225), .O(gate434inter4));
  nand2 gate2120(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2121(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2122(.a(G1057), .O(gate434inter7));
  inv1  gate2123(.a(G1153), .O(gate434inter8));
  nand2 gate2124(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2125(.a(s_225), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2126(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2127(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2128(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate2101(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2102(.a(gate436inter0), .b(s_222), .O(gate436inter1));
  and2  gate2103(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2104(.a(s_222), .O(gate436inter3));
  inv1  gate2105(.a(s_223), .O(gate436inter4));
  nand2 gate2106(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2107(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2108(.a(G1060), .O(gate436inter7));
  inv1  gate2109(.a(G1156), .O(gate436inter8));
  nand2 gate2110(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2111(.a(s_223), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2112(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2113(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2114(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1989(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1990(.a(gate437inter0), .b(s_206), .O(gate437inter1));
  and2  gate1991(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1992(.a(s_206), .O(gate437inter3));
  inv1  gate1993(.a(s_207), .O(gate437inter4));
  nand2 gate1994(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1995(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1996(.a(G10), .O(gate437inter7));
  inv1  gate1997(.a(G1159), .O(gate437inter8));
  nand2 gate1998(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1999(.a(s_207), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2000(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2001(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2002(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2087(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2088(.a(gate438inter0), .b(s_220), .O(gate438inter1));
  and2  gate2089(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2090(.a(s_220), .O(gate438inter3));
  inv1  gate2091(.a(s_221), .O(gate438inter4));
  nand2 gate2092(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2093(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2094(.a(G1063), .O(gate438inter7));
  inv1  gate2095(.a(G1159), .O(gate438inter8));
  nand2 gate2096(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2097(.a(s_221), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2098(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2099(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2100(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate617(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate618(.a(gate439inter0), .b(s_10), .O(gate439inter1));
  and2  gate619(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate620(.a(s_10), .O(gate439inter3));
  inv1  gate621(.a(s_11), .O(gate439inter4));
  nand2 gate622(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate623(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate624(.a(G11), .O(gate439inter7));
  inv1  gate625(.a(G1162), .O(gate439inter8));
  nand2 gate626(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate627(.a(s_11), .b(gate439inter3), .O(gate439inter10));
  nor2  gate628(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate629(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate630(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate589(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate590(.a(gate440inter0), .b(s_6), .O(gate440inter1));
  and2  gate591(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate592(.a(s_6), .O(gate440inter3));
  inv1  gate593(.a(s_7), .O(gate440inter4));
  nand2 gate594(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate595(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate596(.a(G1066), .O(gate440inter7));
  inv1  gate597(.a(G1162), .O(gate440inter8));
  nand2 gate598(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate599(.a(s_7), .b(gate440inter3), .O(gate440inter10));
  nor2  gate600(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate601(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate602(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1051(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1052(.a(gate442inter0), .b(s_72), .O(gate442inter1));
  and2  gate1053(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1054(.a(s_72), .O(gate442inter3));
  inv1  gate1055(.a(s_73), .O(gate442inter4));
  nand2 gate1056(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1057(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1058(.a(G1069), .O(gate442inter7));
  inv1  gate1059(.a(G1165), .O(gate442inter8));
  nand2 gate1060(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1061(.a(s_73), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1062(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1063(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1064(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1891(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1892(.a(gate443inter0), .b(s_192), .O(gate443inter1));
  and2  gate1893(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1894(.a(s_192), .O(gate443inter3));
  inv1  gate1895(.a(s_193), .O(gate443inter4));
  nand2 gate1896(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1897(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1898(.a(G13), .O(gate443inter7));
  inv1  gate1899(.a(G1168), .O(gate443inter8));
  nand2 gate1900(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1901(.a(s_193), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1902(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1903(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1904(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1107(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1108(.a(gate444inter0), .b(s_80), .O(gate444inter1));
  and2  gate1109(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1110(.a(s_80), .O(gate444inter3));
  inv1  gate1111(.a(s_81), .O(gate444inter4));
  nand2 gate1112(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1113(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1114(.a(G1072), .O(gate444inter7));
  inv1  gate1115(.a(G1168), .O(gate444inter8));
  nand2 gate1116(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1117(.a(s_81), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1118(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1119(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1120(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate2941(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2942(.a(gate445inter0), .b(s_342), .O(gate445inter1));
  and2  gate2943(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2944(.a(s_342), .O(gate445inter3));
  inv1  gate2945(.a(s_343), .O(gate445inter4));
  nand2 gate2946(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2947(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2948(.a(G14), .O(gate445inter7));
  inv1  gate2949(.a(G1171), .O(gate445inter8));
  nand2 gate2950(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2951(.a(s_343), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2952(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2953(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2954(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1569(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1570(.a(gate446inter0), .b(s_146), .O(gate446inter1));
  and2  gate1571(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1572(.a(s_146), .O(gate446inter3));
  inv1  gate1573(.a(s_147), .O(gate446inter4));
  nand2 gate1574(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1575(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1576(.a(G1075), .O(gate446inter7));
  inv1  gate1577(.a(G1171), .O(gate446inter8));
  nand2 gate1578(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1579(.a(s_147), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1580(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1581(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1582(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate3151(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate3152(.a(gate451inter0), .b(s_372), .O(gate451inter1));
  and2  gate3153(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate3154(.a(s_372), .O(gate451inter3));
  inv1  gate3155(.a(s_373), .O(gate451inter4));
  nand2 gate3156(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate3157(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate3158(.a(G17), .O(gate451inter7));
  inv1  gate3159(.a(G1180), .O(gate451inter8));
  nand2 gate3160(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate3161(.a(s_373), .b(gate451inter3), .O(gate451inter10));
  nor2  gate3162(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate3163(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate3164(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate841(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate842(.a(gate453inter0), .b(s_42), .O(gate453inter1));
  and2  gate843(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate844(.a(s_42), .O(gate453inter3));
  inv1  gate845(.a(s_43), .O(gate453inter4));
  nand2 gate846(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate847(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate848(.a(G18), .O(gate453inter7));
  inv1  gate849(.a(G1183), .O(gate453inter8));
  nand2 gate850(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate851(.a(s_43), .b(gate453inter3), .O(gate453inter10));
  nor2  gate852(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate853(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate854(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate813(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate814(.a(gate456inter0), .b(s_38), .O(gate456inter1));
  and2  gate815(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate816(.a(s_38), .O(gate456inter3));
  inv1  gate817(.a(s_39), .O(gate456inter4));
  nand2 gate818(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate819(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate820(.a(G1090), .O(gate456inter7));
  inv1  gate821(.a(G1186), .O(gate456inter8));
  nand2 gate822(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate823(.a(s_39), .b(gate456inter3), .O(gate456inter10));
  nor2  gate824(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate825(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate826(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1653(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1654(.a(gate457inter0), .b(s_158), .O(gate457inter1));
  and2  gate1655(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1656(.a(s_158), .O(gate457inter3));
  inv1  gate1657(.a(s_159), .O(gate457inter4));
  nand2 gate1658(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1659(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1660(.a(G20), .O(gate457inter7));
  inv1  gate1661(.a(G1189), .O(gate457inter8));
  nand2 gate1662(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1663(.a(s_159), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1664(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1665(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1666(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1625(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1626(.a(gate460inter0), .b(s_154), .O(gate460inter1));
  and2  gate1627(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1628(.a(s_154), .O(gate460inter3));
  inv1  gate1629(.a(s_155), .O(gate460inter4));
  nand2 gate1630(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1631(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1632(.a(G1096), .O(gate460inter7));
  inv1  gate1633(.a(G1192), .O(gate460inter8));
  nand2 gate1634(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1635(.a(s_155), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1636(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1637(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1638(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1583(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1584(.a(gate462inter0), .b(s_148), .O(gate462inter1));
  and2  gate1585(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1586(.a(s_148), .O(gate462inter3));
  inv1  gate1587(.a(s_149), .O(gate462inter4));
  nand2 gate1588(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1589(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1590(.a(G1099), .O(gate462inter7));
  inv1  gate1591(.a(G1195), .O(gate462inter8));
  nand2 gate1592(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1593(.a(s_149), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1594(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1595(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1596(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate799(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate800(.a(gate463inter0), .b(s_36), .O(gate463inter1));
  and2  gate801(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate802(.a(s_36), .O(gate463inter3));
  inv1  gate803(.a(s_37), .O(gate463inter4));
  nand2 gate804(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate805(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate806(.a(G23), .O(gate463inter7));
  inv1  gate807(.a(G1198), .O(gate463inter8));
  nand2 gate808(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate809(.a(s_37), .b(gate463inter3), .O(gate463inter10));
  nor2  gate810(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate811(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate812(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1219(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1220(.a(gate466inter0), .b(s_96), .O(gate466inter1));
  and2  gate1221(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1222(.a(s_96), .O(gate466inter3));
  inv1  gate1223(.a(s_97), .O(gate466inter4));
  nand2 gate1224(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1225(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1226(.a(G1105), .O(gate466inter7));
  inv1  gate1227(.a(G1201), .O(gate466inter8));
  nand2 gate1228(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1229(.a(s_97), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1230(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1231(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1232(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1079(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1080(.a(gate468inter0), .b(s_76), .O(gate468inter1));
  and2  gate1081(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1082(.a(s_76), .O(gate468inter3));
  inv1  gate1083(.a(s_77), .O(gate468inter4));
  nand2 gate1084(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1085(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1086(.a(G1108), .O(gate468inter7));
  inv1  gate1087(.a(G1204), .O(gate468inter8));
  nand2 gate1088(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1089(.a(s_77), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1090(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1091(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1092(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate645(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate646(.a(gate469inter0), .b(s_14), .O(gate469inter1));
  and2  gate647(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate648(.a(s_14), .O(gate469inter3));
  inv1  gate649(.a(s_15), .O(gate469inter4));
  nand2 gate650(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate651(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate652(.a(G26), .O(gate469inter7));
  inv1  gate653(.a(G1207), .O(gate469inter8));
  nand2 gate654(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate655(.a(s_15), .b(gate469inter3), .O(gate469inter10));
  nor2  gate656(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate657(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate658(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1317(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1318(.a(gate474inter0), .b(s_110), .O(gate474inter1));
  and2  gate1319(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1320(.a(s_110), .O(gate474inter3));
  inv1  gate1321(.a(s_111), .O(gate474inter4));
  nand2 gate1322(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1323(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1324(.a(G1117), .O(gate474inter7));
  inv1  gate1325(.a(G1213), .O(gate474inter8));
  nand2 gate1326(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1327(.a(s_111), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1328(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1329(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1330(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate673(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate674(.a(gate476inter0), .b(s_18), .O(gate476inter1));
  and2  gate675(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate676(.a(s_18), .O(gate476inter3));
  inv1  gate677(.a(s_19), .O(gate476inter4));
  nand2 gate678(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate679(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate680(.a(G1120), .O(gate476inter7));
  inv1  gate681(.a(G1216), .O(gate476inter8));
  nand2 gate682(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate683(.a(s_19), .b(gate476inter3), .O(gate476inter10));
  nor2  gate684(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate685(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate686(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1513(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1514(.a(gate479inter0), .b(s_138), .O(gate479inter1));
  and2  gate1515(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1516(.a(s_138), .O(gate479inter3));
  inv1  gate1517(.a(s_139), .O(gate479inter4));
  nand2 gate1518(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1519(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1520(.a(G31), .O(gate479inter7));
  inv1  gate1521(.a(G1222), .O(gate479inter8));
  nand2 gate1522(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1523(.a(s_139), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1524(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1525(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1526(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2493(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2494(.a(gate483inter0), .b(s_278), .O(gate483inter1));
  and2  gate2495(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2496(.a(s_278), .O(gate483inter3));
  inv1  gate2497(.a(s_279), .O(gate483inter4));
  nand2 gate2498(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2499(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2500(.a(G1228), .O(gate483inter7));
  inv1  gate2501(.a(G1229), .O(gate483inter8));
  nand2 gate2502(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2503(.a(s_279), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2504(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2505(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2506(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate3011(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate3012(.a(gate484inter0), .b(s_352), .O(gate484inter1));
  and2  gate3013(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate3014(.a(s_352), .O(gate484inter3));
  inv1  gate3015(.a(s_353), .O(gate484inter4));
  nand2 gate3016(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate3017(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate3018(.a(G1230), .O(gate484inter7));
  inv1  gate3019(.a(G1231), .O(gate484inter8));
  nand2 gate3020(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate3021(.a(s_353), .b(gate484inter3), .O(gate484inter10));
  nor2  gate3022(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate3023(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate3024(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2451(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2452(.a(gate485inter0), .b(s_272), .O(gate485inter1));
  and2  gate2453(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2454(.a(s_272), .O(gate485inter3));
  inv1  gate2455(.a(s_273), .O(gate485inter4));
  nand2 gate2456(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2457(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2458(.a(G1232), .O(gate485inter7));
  inv1  gate2459(.a(G1233), .O(gate485inter8));
  nand2 gate2460(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2461(.a(s_273), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2462(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2463(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2464(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1597(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1598(.a(gate487inter0), .b(s_150), .O(gate487inter1));
  and2  gate1599(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1600(.a(s_150), .O(gate487inter3));
  inv1  gate1601(.a(s_151), .O(gate487inter4));
  nand2 gate1602(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1603(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1604(.a(G1236), .O(gate487inter7));
  inv1  gate1605(.a(G1237), .O(gate487inter8));
  nand2 gate1606(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1607(.a(s_151), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1608(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1609(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1610(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate883(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate884(.a(gate491inter0), .b(s_48), .O(gate491inter1));
  and2  gate885(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate886(.a(s_48), .O(gate491inter3));
  inv1  gate887(.a(s_49), .O(gate491inter4));
  nand2 gate888(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate889(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate890(.a(G1244), .O(gate491inter7));
  inv1  gate891(.a(G1245), .O(gate491inter8));
  nand2 gate892(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate893(.a(s_49), .b(gate491inter3), .O(gate491inter10));
  nor2  gate894(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate895(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate896(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1835(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1836(.a(gate494inter0), .b(s_184), .O(gate494inter1));
  and2  gate1837(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1838(.a(s_184), .O(gate494inter3));
  inv1  gate1839(.a(s_185), .O(gate494inter4));
  nand2 gate1840(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1841(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1842(.a(G1250), .O(gate494inter7));
  inv1  gate1843(.a(G1251), .O(gate494inter8));
  nand2 gate1844(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1845(.a(s_185), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1846(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1847(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1848(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2577(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2578(.a(gate495inter0), .b(s_290), .O(gate495inter1));
  and2  gate2579(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2580(.a(s_290), .O(gate495inter3));
  inv1  gate2581(.a(s_291), .O(gate495inter4));
  nand2 gate2582(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2583(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2584(.a(G1252), .O(gate495inter7));
  inv1  gate2585(.a(G1253), .O(gate495inter8));
  nand2 gate2586(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2587(.a(s_291), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2588(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2589(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2590(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2325(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2326(.a(gate500inter0), .b(s_254), .O(gate500inter1));
  and2  gate2327(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2328(.a(s_254), .O(gate500inter3));
  inv1  gate2329(.a(s_255), .O(gate500inter4));
  nand2 gate2330(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2331(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2332(.a(G1262), .O(gate500inter7));
  inv1  gate2333(.a(G1263), .O(gate500inter8));
  nand2 gate2334(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2335(.a(s_255), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2336(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2337(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2338(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2283(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2284(.a(gate502inter0), .b(s_248), .O(gate502inter1));
  and2  gate2285(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2286(.a(s_248), .O(gate502inter3));
  inv1  gate2287(.a(s_249), .O(gate502inter4));
  nand2 gate2288(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2289(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2290(.a(G1266), .O(gate502inter7));
  inv1  gate2291(.a(G1267), .O(gate502inter8));
  nand2 gate2292(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2293(.a(s_249), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2294(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2295(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2296(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate603(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate604(.a(gate504inter0), .b(s_8), .O(gate504inter1));
  and2  gate605(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate606(.a(s_8), .O(gate504inter3));
  inv1  gate607(.a(s_9), .O(gate504inter4));
  nand2 gate608(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate609(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate610(.a(G1270), .O(gate504inter7));
  inv1  gate611(.a(G1271), .O(gate504inter8));
  nand2 gate612(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate613(.a(s_9), .b(gate504inter3), .O(gate504inter10));
  nor2  gate614(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate615(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate616(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1541(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1542(.a(gate506inter0), .b(s_142), .O(gate506inter1));
  and2  gate1543(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1544(.a(s_142), .O(gate506inter3));
  inv1  gate1545(.a(s_143), .O(gate506inter4));
  nand2 gate1546(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1547(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1548(.a(G1274), .O(gate506inter7));
  inv1  gate1549(.a(G1275), .O(gate506inter8));
  nand2 gate1550(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1551(.a(s_143), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1552(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1553(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1554(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1667(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1668(.a(gate507inter0), .b(s_160), .O(gate507inter1));
  and2  gate1669(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1670(.a(s_160), .O(gate507inter3));
  inv1  gate1671(.a(s_161), .O(gate507inter4));
  nand2 gate1672(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1673(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1674(.a(G1276), .O(gate507inter7));
  inv1  gate1675(.a(G1277), .O(gate507inter8));
  nand2 gate1676(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1677(.a(s_161), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1678(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1679(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1680(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1037(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1038(.a(gate511inter0), .b(s_70), .O(gate511inter1));
  and2  gate1039(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1040(.a(s_70), .O(gate511inter3));
  inv1  gate1041(.a(s_71), .O(gate511inter4));
  nand2 gate1042(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1043(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1044(.a(G1284), .O(gate511inter7));
  inv1  gate1045(.a(G1285), .O(gate511inter8));
  nand2 gate1046(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1047(.a(s_71), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1048(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1049(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1050(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate939(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate940(.a(gate513inter0), .b(s_56), .O(gate513inter1));
  and2  gate941(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate942(.a(s_56), .O(gate513inter3));
  inv1  gate943(.a(s_57), .O(gate513inter4));
  nand2 gate944(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate945(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate946(.a(G1288), .O(gate513inter7));
  inv1  gate947(.a(G1289), .O(gate513inter8));
  nand2 gate948(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate949(.a(s_57), .b(gate513inter3), .O(gate513inter10));
  nor2  gate950(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate951(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate952(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule