module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate329(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate330(.a(gate22inter0), .b(s_24), .O(gate22inter1));
  and2  gate331(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate332(.a(s_24), .O(gate22inter3));
  inv1  gate333(.a(s_25), .O(gate22inter4));
  nand2 gate334(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate335(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate336(.a(N122), .O(gate22inter7));
  inv1  gate337(.a(N17), .O(gate22inter8));
  nand2 gate338(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate339(.a(s_25), .b(gate22inter3), .O(gate22inter10));
  nor2  gate340(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate341(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate342(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate161(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate162(.a(gate24inter0), .b(s_0), .O(gate24inter1));
  and2  gate163(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate164(.a(s_0), .O(gate24inter3));
  inv1  gate165(.a(s_1), .O(gate24inter4));
  nand2 gate166(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate167(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate168(.a(N130), .O(gate24inter7));
  inv1  gate169(.a(N43), .O(gate24inter8));
  nand2 gate170(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate171(.a(s_1), .b(gate24inter3), .O(gate24inter10));
  nor2  gate172(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate173(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate174(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate189(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate190(.a(gate27inter0), .b(s_4), .O(gate27inter1));
  and2  gate191(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate192(.a(s_4), .O(gate27inter3));
  inv1  gate193(.a(s_5), .O(gate27inter4));
  nand2 gate194(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate195(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate196(.a(N142), .O(gate27inter7));
  inv1  gate197(.a(N82), .O(gate27inter8));
  nand2 gate198(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate199(.a(s_5), .b(gate27inter3), .O(gate27inter10));
  nor2  gate200(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate201(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate202(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate315(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate316(.a(gate36inter0), .b(s_22), .O(gate36inter1));
  and2  gate317(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate318(.a(s_22), .O(gate36inter3));
  inv1  gate319(.a(s_23), .O(gate36inter4));
  nand2 gate320(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate321(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate322(.a(N60), .O(gate36inter7));
  inv1  gate323(.a(N135), .O(gate36inter8));
  nand2 gate324(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate325(.a(s_23), .b(gate36inter3), .O(gate36inter10));
  nor2  gate326(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate327(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate328(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate231(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate232(.a(gate40inter0), .b(s_10), .O(gate40inter1));
  and2  gate233(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate234(.a(s_10), .O(gate40inter3));
  inv1  gate235(.a(s_11), .O(gate40inter4));
  nand2 gate236(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate237(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate238(.a(N86), .O(gate40inter7));
  inv1  gate239(.a(N143), .O(gate40inter8));
  nand2 gate240(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate241(.a(s_11), .b(gate40inter3), .O(gate40inter10));
  nor2  gate242(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate243(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate244(.a(gate40inter12), .b(gate40inter1), .O(N193));
nor2 gate41( .a(N92), .b(N143), .O(N194) );

  xor2  gate413(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate414(.a(gate42inter0), .b(s_36), .O(gate42inter1));
  and2  gate415(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate416(.a(s_36), .O(gate42inter3));
  inv1  gate417(.a(s_37), .O(gate42inter4));
  nand2 gate418(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate419(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate420(.a(N99), .O(gate42inter7));
  inv1  gate421(.a(N147), .O(gate42inter8));
  nand2 gate422(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate423(.a(s_37), .b(gate42inter3), .O(gate42inter10));
  nor2  gate424(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate425(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate426(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );

  xor2  gate259(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate260(.a(gate44inter0), .b(s_14), .O(gate44inter1));
  and2  gate261(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate262(.a(s_14), .O(gate44inter3));
  inv1  gate263(.a(s_15), .O(gate44inter4));
  nand2 gate264(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate265(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate266(.a(N112), .O(gate44inter7));
  inv1  gate267(.a(N151), .O(gate44inter8));
  nand2 gate268(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate269(.a(s_15), .b(gate44inter3), .O(gate44inter10));
  nor2  gate270(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate271(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate272(.a(gate44inter12), .b(gate44inter1), .O(N197));
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );

  xor2  gate399(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate400(.a(gate57inter0), .b(s_34), .O(gate57inter1));
  and2  gate401(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate402(.a(s_34), .O(gate57inter3));
  inv1  gate403(.a(s_35), .O(gate57inter4));
  nand2 gate404(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate405(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate406(.a(N203), .O(gate57inter7));
  inv1  gate407(.a(N174), .O(gate57inter8));
  nand2 gate408(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate409(.a(s_35), .b(gate57inter3), .O(gate57inter10));
  nor2  gate410(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate411(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate412(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );

  xor2  gate371(.a(N180), .b(N203), .O(gate61inter0));
  nand2 gate372(.a(gate61inter0), .b(s_30), .O(gate61inter1));
  and2  gate373(.a(N180), .b(N203), .O(gate61inter2));
  inv1  gate374(.a(s_30), .O(gate61inter3));
  inv1  gate375(.a(s_31), .O(gate61inter4));
  nand2 gate376(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate377(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate378(.a(N203), .O(gate61inter7));
  inv1  gate379(.a(N180), .O(gate61inter8));
  nand2 gate380(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate381(.a(s_31), .b(gate61inter3), .O(gate61inter10));
  nor2  gate382(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate383(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate384(.a(gate61inter12), .b(gate61inter1), .O(N251));
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );

  xor2  gate343(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate344(.a(gate67inter0), .b(s_26), .O(gate67inter1));
  and2  gate345(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate346(.a(s_26), .O(gate67inter3));
  inv1  gate347(.a(s_27), .O(gate67inter4));
  nand2 gate348(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate349(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate350(.a(N213), .O(gate67inter7));
  inv1  gate351(.a(N102), .O(gate67inter8));
  nand2 gate352(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate353(.a(s_27), .b(gate67inter3), .O(gate67inter10));
  nor2  gate354(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate355(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate356(.a(gate67inter12), .b(gate67inter1), .O(N259));
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate273(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate274(.a(gate71inter0), .b(s_16), .O(gate71inter1));
  and2  gate275(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate276(.a(s_16), .O(gate71inter3));
  inv1  gate277(.a(s_17), .O(gate71inter4));
  nand2 gate278(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate279(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate280(.a(N230), .O(gate71inter7));
  inv1  gate281(.a(N185), .O(gate71inter8));
  nand2 gate282(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate283(.a(s_17), .b(gate71inter3), .O(gate71inter10));
  nor2  gate284(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate285(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate286(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate357(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate358(.a(gate83inter0), .b(s_28), .O(gate83inter1));
  and2  gate359(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate360(.a(s_28), .O(gate83inter3));
  inv1  gate361(.a(s_29), .O(gate83inter4));
  nand2 gate362(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate363(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate364(.a(N243), .O(gate83inter7));
  inv1  gate365(.a(N194), .O(gate83inter8));
  nand2 gate366(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate367(.a(s_29), .b(gate83inter3), .O(gate83inter10));
  nor2  gate368(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate369(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate370(.a(gate83inter12), .b(gate83inter1), .O(N293));
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate385(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate386(.a(gate99inter0), .b(s_32), .O(gate99inter1));
  and2  gate387(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate388(.a(s_32), .O(gate99inter3));
  inv1  gate389(.a(s_33), .O(gate99inter4));
  nand2 gate390(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate391(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate392(.a(N309), .O(gate99inter7));
  inv1  gate393(.a(N260), .O(gate99inter8));
  nand2 gate394(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate395(.a(s_33), .b(gate99inter3), .O(gate99inter10));
  nor2  gate396(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate397(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate398(.a(gate99inter12), .b(gate99inter1), .O(N330));
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );

  xor2  gate427(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate428(.a(gate104inter0), .b(s_38), .O(gate104inter1));
  and2  gate429(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate430(.a(s_38), .O(gate104inter3));
  inv1  gate431(.a(s_39), .O(gate104inter4));
  nand2 gate432(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate433(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate434(.a(N309), .O(gate104inter7));
  inv1  gate435(.a(N273), .O(gate104inter8));
  nand2 gate436(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate437(.a(s_39), .b(gate104inter3), .O(gate104inter10));
  nor2  gate438(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate439(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate440(.a(gate104inter12), .b(gate104inter1), .O(N335));
nand2 gate105( .a(N319), .b(N21), .O(N336) );

  xor2  gate301(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate302(.a(gate106inter0), .b(s_20), .O(gate106inter1));
  and2  gate303(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate304(.a(s_20), .O(gate106inter3));
  inv1  gate305(.a(s_21), .O(gate106inter4));
  nand2 gate306(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate307(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate308(.a(N309), .O(gate106inter7));
  inv1  gate309(.a(N276), .O(gate106inter8));
  nand2 gate310(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate311(.a(s_21), .b(gate106inter3), .O(gate106inter10));
  nor2  gate312(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate313(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate314(.a(gate106inter12), .b(gate106inter1), .O(N337));
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );

  xor2  gate217(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate218(.a(gate109inter0), .b(s_8), .O(gate109inter1));
  and2  gate219(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate220(.a(s_8), .O(gate109inter3));
  inv1  gate221(.a(s_9), .O(gate109inter4));
  nand2 gate222(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate223(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate224(.a(N319), .O(gate109inter7));
  inv1  gate225(.a(N47), .O(gate109inter8));
  nand2 gate226(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate227(.a(s_9), .b(gate109inter3), .O(gate109inter10));
  nor2  gate228(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate229(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate230(.a(gate109inter12), .b(gate109inter1), .O(N340));
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );

  xor2  gate287(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate288(.a(gate114inter0), .b(s_18), .O(gate114inter1));
  and2  gate289(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate290(.a(s_18), .O(gate114inter3));
  inv1  gate291(.a(s_19), .O(gate114inter4));
  nand2 gate292(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate293(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate294(.a(N319), .O(gate114inter7));
  inv1  gate295(.a(N86), .O(gate114inter8));
  nand2 gate296(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate297(.a(s_19), .b(gate114inter3), .O(gate114inter10));
  nor2  gate298(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate299(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate300(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );

  xor2  gate441(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate442(.a(gate130inter0), .b(s_40), .O(gate130inter1));
  and2  gate443(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate444(.a(s_40), .O(gate130inter3));
  inv1  gate445(.a(s_41), .O(gate130inter4));
  nand2 gate446(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate447(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate448(.a(N360), .O(gate130inter7));
  inv1  gate449(.a(N27), .O(gate130inter8));
  nand2 gate450(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate451(.a(s_41), .b(gate130inter3), .O(gate130inter10));
  nor2  gate452(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate453(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate454(.a(gate130inter12), .b(gate130inter1), .O(N372));
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate175(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate176(.a(gate132inter0), .b(s_2), .O(gate132inter1));
  and2  gate177(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate178(.a(s_2), .O(gate132inter3));
  inv1  gate179(.a(s_3), .O(gate132inter4));
  nand2 gate180(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate181(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate182(.a(N360), .O(gate132inter7));
  inv1  gate183(.a(N53), .O(gate132inter8));
  nand2 gate184(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate185(.a(s_3), .b(gate132inter3), .O(gate132inter10));
  nor2  gate186(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate187(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate188(.a(gate132inter12), .b(gate132inter1), .O(N374));

  xor2  gate203(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate204(.a(gate133inter0), .b(s_6), .O(gate133inter1));
  and2  gate205(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate206(.a(s_6), .O(gate133inter3));
  inv1  gate207(.a(s_7), .O(gate133inter4));
  nand2 gate208(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate209(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate210(.a(N360), .O(gate133inter7));
  inv1  gate211(.a(N66), .O(gate133inter8));
  nand2 gate212(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate213(.a(s_7), .b(gate133inter3), .O(gate133inter10));
  nor2  gate214(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate215(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate216(.a(gate133inter12), .b(gate133inter1), .O(N375));
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );

  xor2  gate245(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate246(.a(gate154inter0), .b(s_12), .O(gate154inter1));
  and2  gate247(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate248(.a(s_12), .O(gate154inter3));
  inv1  gate249(.a(s_13), .O(gate154inter4));
  nand2 gate250(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate251(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate252(.a(N386), .O(gate154inter7));
  inv1  gate253(.a(N417), .O(gate154inter8));
  nand2 gate254(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate255(.a(s_13), .b(gate154inter3), .O(gate154inter10));
  nor2  gate256(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate257(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate258(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule