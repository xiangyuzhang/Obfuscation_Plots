module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1877(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1878(.a(gate13inter0), .b(s_190), .O(gate13inter1));
  and2  gate1879(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1880(.a(s_190), .O(gate13inter3));
  inv1  gate1881(.a(s_191), .O(gate13inter4));
  nand2 gate1882(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1883(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1884(.a(G9), .O(gate13inter7));
  inv1  gate1885(.a(G10), .O(gate13inter8));
  nand2 gate1886(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1887(.a(s_191), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1888(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1889(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1890(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1387(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1388(.a(gate21inter0), .b(s_120), .O(gate21inter1));
  and2  gate1389(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1390(.a(s_120), .O(gate21inter3));
  inv1  gate1391(.a(s_121), .O(gate21inter4));
  nand2 gate1392(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1393(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1394(.a(G25), .O(gate21inter7));
  inv1  gate1395(.a(G26), .O(gate21inter8));
  nand2 gate1396(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1397(.a(s_121), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1398(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1399(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1400(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1191(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1192(.a(gate22inter0), .b(s_92), .O(gate22inter1));
  and2  gate1193(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1194(.a(s_92), .O(gate22inter3));
  inv1  gate1195(.a(s_93), .O(gate22inter4));
  nand2 gate1196(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1197(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1198(.a(G27), .O(gate22inter7));
  inv1  gate1199(.a(G28), .O(gate22inter8));
  nand2 gate1200(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1201(.a(s_93), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1202(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1203(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1204(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2017(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2018(.a(gate24inter0), .b(s_210), .O(gate24inter1));
  and2  gate2019(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2020(.a(s_210), .O(gate24inter3));
  inv1  gate2021(.a(s_211), .O(gate24inter4));
  nand2 gate2022(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2023(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2024(.a(G31), .O(gate24inter7));
  inv1  gate2025(.a(G32), .O(gate24inter8));
  nand2 gate2026(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2027(.a(s_211), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2028(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2029(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2030(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2283(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2284(.a(gate26inter0), .b(s_248), .O(gate26inter1));
  and2  gate2285(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2286(.a(s_248), .O(gate26inter3));
  inv1  gate2287(.a(s_249), .O(gate26inter4));
  nand2 gate2288(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2289(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2290(.a(G9), .O(gate26inter7));
  inv1  gate2291(.a(G13), .O(gate26inter8));
  nand2 gate2292(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2293(.a(s_249), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2294(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2295(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2296(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1373(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1374(.a(gate29inter0), .b(s_118), .O(gate29inter1));
  and2  gate1375(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1376(.a(s_118), .O(gate29inter3));
  inv1  gate1377(.a(s_119), .O(gate29inter4));
  nand2 gate1378(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1379(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1380(.a(G3), .O(gate29inter7));
  inv1  gate1381(.a(G7), .O(gate29inter8));
  nand2 gate1382(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1383(.a(s_119), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1384(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1385(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1386(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1415(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1416(.a(gate32inter0), .b(s_124), .O(gate32inter1));
  and2  gate1417(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1418(.a(s_124), .O(gate32inter3));
  inv1  gate1419(.a(s_125), .O(gate32inter4));
  nand2 gate1420(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1421(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1422(.a(G12), .O(gate32inter7));
  inv1  gate1423(.a(G16), .O(gate32inter8));
  nand2 gate1424(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1425(.a(s_125), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1426(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1427(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1428(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate617(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate618(.a(gate33inter0), .b(s_10), .O(gate33inter1));
  and2  gate619(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate620(.a(s_10), .O(gate33inter3));
  inv1  gate621(.a(s_11), .O(gate33inter4));
  nand2 gate622(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate623(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate624(.a(G17), .O(gate33inter7));
  inv1  gate625(.a(G21), .O(gate33inter8));
  nand2 gate626(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate627(.a(s_11), .b(gate33inter3), .O(gate33inter10));
  nor2  gate628(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate629(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate630(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1499(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1500(.a(gate34inter0), .b(s_136), .O(gate34inter1));
  and2  gate1501(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1502(.a(s_136), .O(gate34inter3));
  inv1  gate1503(.a(s_137), .O(gate34inter4));
  nand2 gate1504(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1505(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1506(.a(G25), .O(gate34inter7));
  inv1  gate1507(.a(G29), .O(gate34inter8));
  nand2 gate1508(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1509(.a(s_137), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1510(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1511(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1512(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate561(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate562(.a(gate35inter0), .b(s_2), .O(gate35inter1));
  and2  gate563(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate564(.a(s_2), .O(gate35inter3));
  inv1  gate565(.a(s_3), .O(gate35inter4));
  nand2 gate566(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate567(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate568(.a(G18), .O(gate35inter7));
  inv1  gate569(.a(G22), .O(gate35inter8));
  nand2 gate570(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate571(.a(s_3), .b(gate35inter3), .O(gate35inter10));
  nor2  gate572(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate573(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate574(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2255(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2256(.a(gate36inter0), .b(s_244), .O(gate36inter1));
  and2  gate2257(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2258(.a(s_244), .O(gate36inter3));
  inv1  gate2259(.a(s_245), .O(gate36inter4));
  nand2 gate2260(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2261(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2262(.a(G26), .O(gate36inter7));
  inv1  gate2263(.a(G30), .O(gate36inter8));
  nand2 gate2264(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2265(.a(s_245), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2266(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2267(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2268(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1513(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1514(.a(gate37inter0), .b(s_138), .O(gate37inter1));
  and2  gate1515(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1516(.a(s_138), .O(gate37inter3));
  inv1  gate1517(.a(s_139), .O(gate37inter4));
  nand2 gate1518(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1519(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1520(.a(G19), .O(gate37inter7));
  inv1  gate1521(.a(G23), .O(gate37inter8));
  nand2 gate1522(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1523(.a(s_139), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1524(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1525(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1526(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1065(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1066(.a(gate38inter0), .b(s_74), .O(gate38inter1));
  and2  gate1067(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1068(.a(s_74), .O(gate38inter3));
  inv1  gate1069(.a(s_75), .O(gate38inter4));
  nand2 gate1070(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1071(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1072(.a(G27), .O(gate38inter7));
  inv1  gate1073(.a(G31), .O(gate38inter8));
  nand2 gate1074(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1075(.a(s_75), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1076(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1077(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1078(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate981(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate982(.a(gate39inter0), .b(s_62), .O(gate39inter1));
  and2  gate983(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate984(.a(s_62), .O(gate39inter3));
  inv1  gate985(.a(s_63), .O(gate39inter4));
  nand2 gate986(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate987(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate988(.a(G20), .O(gate39inter7));
  inv1  gate989(.a(G24), .O(gate39inter8));
  nand2 gate990(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate991(.a(s_63), .b(gate39inter3), .O(gate39inter10));
  nor2  gate992(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate993(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate994(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1135(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1136(.a(gate42inter0), .b(s_84), .O(gate42inter1));
  and2  gate1137(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1138(.a(s_84), .O(gate42inter3));
  inv1  gate1139(.a(s_85), .O(gate42inter4));
  nand2 gate1140(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1141(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1142(.a(G2), .O(gate42inter7));
  inv1  gate1143(.a(G266), .O(gate42inter8));
  nand2 gate1144(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1145(.a(s_85), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1146(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1147(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1148(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1233(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1234(.a(gate43inter0), .b(s_98), .O(gate43inter1));
  and2  gate1235(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1236(.a(s_98), .O(gate43inter3));
  inv1  gate1237(.a(s_99), .O(gate43inter4));
  nand2 gate1238(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1239(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1240(.a(G3), .O(gate43inter7));
  inv1  gate1241(.a(G269), .O(gate43inter8));
  nand2 gate1242(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1243(.a(s_99), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1244(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1245(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1246(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate715(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate716(.a(gate50inter0), .b(s_24), .O(gate50inter1));
  and2  gate717(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate718(.a(s_24), .O(gate50inter3));
  inv1  gate719(.a(s_25), .O(gate50inter4));
  nand2 gate720(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate721(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate722(.a(G10), .O(gate50inter7));
  inv1  gate723(.a(G278), .O(gate50inter8));
  nand2 gate724(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate725(.a(s_25), .b(gate50inter3), .O(gate50inter10));
  nor2  gate726(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate727(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate728(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate729(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate730(.a(gate51inter0), .b(s_26), .O(gate51inter1));
  and2  gate731(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate732(.a(s_26), .O(gate51inter3));
  inv1  gate733(.a(s_27), .O(gate51inter4));
  nand2 gate734(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate735(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate736(.a(G11), .O(gate51inter7));
  inv1  gate737(.a(G281), .O(gate51inter8));
  nand2 gate738(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate739(.a(s_27), .b(gate51inter3), .O(gate51inter10));
  nor2  gate740(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate741(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate742(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1261(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1262(.a(gate52inter0), .b(s_102), .O(gate52inter1));
  and2  gate1263(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1264(.a(s_102), .O(gate52inter3));
  inv1  gate1265(.a(s_103), .O(gate52inter4));
  nand2 gate1266(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1267(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1268(.a(G12), .O(gate52inter7));
  inv1  gate1269(.a(G281), .O(gate52inter8));
  nand2 gate1270(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1271(.a(s_103), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1272(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1273(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1274(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1695(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1696(.a(gate54inter0), .b(s_164), .O(gate54inter1));
  and2  gate1697(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1698(.a(s_164), .O(gate54inter3));
  inv1  gate1699(.a(s_165), .O(gate54inter4));
  nand2 gate1700(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1701(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1702(.a(G14), .O(gate54inter7));
  inv1  gate1703(.a(G284), .O(gate54inter8));
  nand2 gate1704(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1705(.a(s_165), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1706(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1707(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1708(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate2143(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2144(.a(gate57inter0), .b(s_228), .O(gate57inter1));
  and2  gate2145(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2146(.a(s_228), .O(gate57inter3));
  inv1  gate2147(.a(s_229), .O(gate57inter4));
  nand2 gate2148(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2149(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2150(.a(G17), .O(gate57inter7));
  inv1  gate2151(.a(G290), .O(gate57inter8));
  nand2 gate2152(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2153(.a(s_229), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2154(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2155(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2156(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1709(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1710(.a(gate58inter0), .b(s_166), .O(gate58inter1));
  and2  gate1711(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1712(.a(s_166), .O(gate58inter3));
  inv1  gate1713(.a(s_167), .O(gate58inter4));
  nand2 gate1714(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1715(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1716(.a(G18), .O(gate58inter7));
  inv1  gate1717(.a(G290), .O(gate58inter8));
  nand2 gate1718(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1719(.a(s_167), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1720(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1721(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1722(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate897(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate898(.a(gate65inter0), .b(s_50), .O(gate65inter1));
  and2  gate899(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate900(.a(s_50), .O(gate65inter3));
  inv1  gate901(.a(s_51), .O(gate65inter4));
  nand2 gate902(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate903(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate904(.a(G25), .O(gate65inter7));
  inv1  gate905(.a(G302), .O(gate65inter8));
  nand2 gate906(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate907(.a(s_51), .b(gate65inter3), .O(gate65inter10));
  nor2  gate908(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate909(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate910(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate855(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate856(.a(gate66inter0), .b(s_44), .O(gate66inter1));
  and2  gate857(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate858(.a(s_44), .O(gate66inter3));
  inv1  gate859(.a(s_45), .O(gate66inter4));
  nand2 gate860(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate861(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate862(.a(G26), .O(gate66inter7));
  inv1  gate863(.a(G302), .O(gate66inter8));
  nand2 gate864(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate865(.a(s_45), .b(gate66inter3), .O(gate66inter10));
  nor2  gate866(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate867(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate868(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1555(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1556(.a(gate68inter0), .b(s_144), .O(gate68inter1));
  and2  gate1557(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1558(.a(s_144), .O(gate68inter3));
  inv1  gate1559(.a(s_145), .O(gate68inter4));
  nand2 gate1560(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1561(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1562(.a(G28), .O(gate68inter7));
  inv1  gate1563(.a(G305), .O(gate68inter8));
  nand2 gate1564(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1565(.a(s_145), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1566(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1567(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1568(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1611(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1612(.a(gate71inter0), .b(s_152), .O(gate71inter1));
  and2  gate1613(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1614(.a(s_152), .O(gate71inter3));
  inv1  gate1615(.a(s_153), .O(gate71inter4));
  nand2 gate1616(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1617(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1618(.a(G31), .O(gate71inter7));
  inv1  gate1619(.a(G311), .O(gate71inter8));
  nand2 gate1620(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1621(.a(s_153), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1622(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1623(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1624(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1597(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1598(.a(gate77inter0), .b(s_150), .O(gate77inter1));
  and2  gate1599(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1600(.a(s_150), .O(gate77inter3));
  inv1  gate1601(.a(s_151), .O(gate77inter4));
  nand2 gate1602(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1603(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1604(.a(G2), .O(gate77inter7));
  inv1  gate1605(.a(G320), .O(gate77inter8));
  nand2 gate1606(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1607(.a(s_151), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1608(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1609(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1610(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2073(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2074(.a(gate79inter0), .b(s_218), .O(gate79inter1));
  and2  gate2075(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2076(.a(s_218), .O(gate79inter3));
  inv1  gate2077(.a(s_219), .O(gate79inter4));
  nand2 gate2078(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2079(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2080(.a(G10), .O(gate79inter7));
  inv1  gate2081(.a(G323), .O(gate79inter8));
  nand2 gate2082(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2083(.a(s_219), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2084(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2085(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2086(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1681(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1682(.a(gate80inter0), .b(s_162), .O(gate80inter1));
  and2  gate1683(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1684(.a(s_162), .O(gate80inter3));
  inv1  gate1685(.a(s_163), .O(gate80inter4));
  nand2 gate1686(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1687(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1688(.a(G14), .O(gate80inter7));
  inv1  gate1689(.a(G323), .O(gate80inter8));
  nand2 gate1690(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1691(.a(s_163), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1692(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1693(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1694(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate603(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate604(.a(gate86inter0), .b(s_8), .O(gate86inter1));
  and2  gate605(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate606(.a(s_8), .O(gate86inter3));
  inv1  gate607(.a(s_9), .O(gate86inter4));
  nand2 gate608(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate609(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate610(.a(G8), .O(gate86inter7));
  inv1  gate611(.a(G332), .O(gate86inter8));
  nand2 gate612(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate613(.a(s_9), .b(gate86inter3), .O(gate86inter10));
  nor2  gate614(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate615(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate616(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate785(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate786(.a(gate91inter0), .b(s_34), .O(gate91inter1));
  and2  gate787(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate788(.a(s_34), .O(gate91inter3));
  inv1  gate789(.a(s_35), .O(gate91inter4));
  nand2 gate790(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate791(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate792(.a(G25), .O(gate91inter7));
  inv1  gate793(.a(G341), .O(gate91inter8));
  nand2 gate794(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate795(.a(s_35), .b(gate91inter3), .O(gate91inter10));
  nor2  gate796(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate797(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate798(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate813(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate814(.a(gate92inter0), .b(s_38), .O(gate92inter1));
  and2  gate815(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate816(.a(s_38), .O(gate92inter3));
  inv1  gate817(.a(s_39), .O(gate92inter4));
  nand2 gate818(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate819(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate820(.a(G29), .O(gate92inter7));
  inv1  gate821(.a(G341), .O(gate92inter8));
  nand2 gate822(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate823(.a(s_39), .b(gate92inter3), .O(gate92inter10));
  nor2  gate824(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate825(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate826(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1289(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1290(.a(gate100inter0), .b(s_106), .O(gate100inter1));
  and2  gate1291(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1292(.a(s_106), .O(gate100inter3));
  inv1  gate1293(.a(s_107), .O(gate100inter4));
  nand2 gate1294(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1295(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1296(.a(G31), .O(gate100inter7));
  inv1  gate1297(.a(G353), .O(gate100inter8));
  nand2 gate1298(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1299(.a(s_107), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1300(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1301(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1302(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1205(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1206(.a(gate101inter0), .b(s_94), .O(gate101inter1));
  and2  gate1207(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1208(.a(s_94), .O(gate101inter3));
  inv1  gate1209(.a(s_95), .O(gate101inter4));
  nand2 gate1210(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1211(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1212(.a(G20), .O(gate101inter7));
  inv1  gate1213(.a(G356), .O(gate101inter8));
  nand2 gate1214(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1215(.a(s_95), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1216(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1217(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1218(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1401(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1402(.a(gate108inter0), .b(s_122), .O(gate108inter1));
  and2  gate1403(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1404(.a(s_122), .O(gate108inter3));
  inv1  gate1405(.a(s_123), .O(gate108inter4));
  nand2 gate1406(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1407(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1408(.a(G368), .O(gate108inter7));
  inv1  gate1409(.a(G369), .O(gate108inter8));
  nand2 gate1410(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1411(.a(s_123), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1412(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1413(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1414(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1863(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1864(.a(gate109inter0), .b(s_188), .O(gate109inter1));
  and2  gate1865(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1866(.a(s_188), .O(gate109inter3));
  inv1  gate1867(.a(s_189), .O(gate109inter4));
  nand2 gate1868(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1869(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1870(.a(G370), .O(gate109inter7));
  inv1  gate1871(.a(G371), .O(gate109inter8));
  nand2 gate1872(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1873(.a(s_189), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1874(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1875(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1876(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1485(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1486(.a(gate112inter0), .b(s_134), .O(gate112inter1));
  and2  gate1487(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1488(.a(s_134), .O(gate112inter3));
  inv1  gate1489(.a(s_135), .O(gate112inter4));
  nand2 gate1490(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1491(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1492(.a(G376), .O(gate112inter7));
  inv1  gate1493(.a(G377), .O(gate112inter8));
  nand2 gate1494(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1495(.a(s_135), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1496(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1497(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1498(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1527(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1528(.a(gate119inter0), .b(s_140), .O(gate119inter1));
  and2  gate1529(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1530(.a(s_140), .O(gate119inter3));
  inv1  gate1531(.a(s_141), .O(gate119inter4));
  nand2 gate1532(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1533(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1534(.a(G390), .O(gate119inter7));
  inv1  gate1535(.a(G391), .O(gate119inter8));
  nand2 gate1536(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1537(.a(s_141), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1538(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1539(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1540(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1667(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1668(.a(gate120inter0), .b(s_160), .O(gate120inter1));
  and2  gate1669(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1670(.a(s_160), .O(gate120inter3));
  inv1  gate1671(.a(s_161), .O(gate120inter4));
  nand2 gate1672(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1673(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1674(.a(G392), .O(gate120inter7));
  inv1  gate1675(.a(G393), .O(gate120inter8));
  nand2 gate1676(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1677(.a(s_161), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1678(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1679(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1680(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate673(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate674(.a(gate121inter0), .b(s_18), .O(gate121inter1));
  and2  gate675(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate676(.a(s_18), .O(gate121inter3));
  inv1  gate677(.a(s_19), .O(gate121inter4));
  nand2 gate678(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate679(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate680(.a(G394), .O(gate121inter7));
  inv1  gate681(.a(G395), .O(gate121inter8));
  nand2 gate682(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate683(.a(s_19), .b(gate121inter3), .O(gate121inter10));
  nor2  gate684(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate685(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate686(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1639(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1640(.a(gate122inter0), .b(s_156), .O(gate122inter1));
  and2  gate1641(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1642(.a(s_156), .O(gate122inter3));
  inv1  gate1643(.a(s_157), .O(gate122inter4));
  nand2 gate1644(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1645(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1646(.a(G396), .O(gate122inter7));
  inv1  gate1647(.a(G397), .O(gate122inter8));
  nand2 gate1648(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1649(.a(s_157), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1650(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1651(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1652(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate911(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate912(.a(gate130inter0), .b(s_52), .O(gate130inter1));
  and2  gate913(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate914(.a(s_52), .O(gate130inter3));
  inv1  gate915(.a(s_53), .O(gate130inter4));
  nand2 gate916(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate917(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate918(.a(G412), .O(gate130inter7));
  inv1  gate919(.a(G413), .O(gate130inter8));
  nand2 gate920(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate921(.a(s_53), .b(gate130inter3), .O(gate130inter10));
  nor2  gate922(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate923(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate924(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate799(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate800(.a(gate138inter0), .b(s_36), .O(gate138inter1));
  and2  gate801(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate802(.a(s_36), .O(gate138inter3));
  inv1  gate803(.a(s_37), .O(gate138inter4));
  nand2 gate804(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate805(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate806(.a(G432), .O(gate138inter7));
  inv1  gate807(.a(G435), .O(gate138inter8));
  nand2 gate808(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate809(.a(s_37), .b(gate138inter3), .O(gate138inter10));
  nor2  gate810(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate811(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate812(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2185(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2186(.a(gate140inter0), .b(s_234), .O(gate140inter1));
  and2  gate2187(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2188(.a(s_234), .O(gate140inter3));
  inv1  gate2189(.a(s_235), .O(gate140inter4));
  nand2 gate2190(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2191(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2192(.a(G444), .O(gate140inter7));
  inv1  gate2193(.a(G447), .O(gate140inter8));
  nand2 gate2194(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2195(.a(s_235), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2196(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2197(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2198(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1429(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1430(.a(gate141inter0), .b(s_126), .O(gate141inter1));
  and2  gate1431(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1432(.a(s_126), .O(gate141inter3));
  inv1  gate1433(.a(s_127), .O(gate141inter4));
  nand2 gate1434(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1435(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1436(.a(G450), .O(gate141inter7));
  inv1  gate1437(.a(G453), .O(gate141inter8));
  nand2 gate1438(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1439(.a(s_127), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1440(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1441(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1442(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate939(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate940(.a(gate148inter0), .b(s_56), .O(gate148inter1));
  and2  gate941(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate942(.a(s_56), .O(gate148inter3));
  inv1  gate943(.a(s_57), .O(gate148inter4));
  nand2 gate944(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate945(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate946(.a(G492), .O(gate148inter7));
  inv1  gate947(.a(G495), .O(gate148inter8));
  nand2 gate948(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate949(.a(s_57), .b(gate148inter3), .O(gate148inter10));
  nor2  gate950(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate951(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate952(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate827(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate828(.a(gate149inter0), .b(s_40), .O(gate149inter1));
  and2  gate829(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate830(.a(s_40), .O(gate149inter3));
  inv1  gate831(.a(s_41), .O(gate149inter4));
  nand2 gate832(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate833(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate834(.a(G498), .O(gate149inter7));
  inv1  gate835(.a(G501), .O(gate149inter8));
  nand2 gate836(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate837(.a(s_41), .b(gate149inter3), .O(gate149inter10));
  nor2  gate838(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate839(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate840(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1345(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1346(.a(gate153inter0), .b(s_114), .O(gate153inter1));
  and2  gate1347(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1348(.a(s_114), .O(gate153inter3));
  inv1  gate1349(.a(s_115), .O(gate153inter4));
  nand2 gate1350(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1351(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1352(.a(G426), .O(gate153inter7));
  inv1  gate1353(.a(G522), .O(gate153inter8));
  nand2 gate1354(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1355(.a(s_115), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1356(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1357(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1358(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1023(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1024(.a(gate156inter0), .b(s_68), .O(gate156inter1));
  and2  gate1025(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1026(.a(s_68), .O(gate156inter3));
  inv1  gate1027(.a(s_69), .O(gate156inter4));
  nand2 gate1028(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1029(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1030(.a(G435), .O(gate156inter7));
  inv1  gate1031(.a(G525), .O(gate156inter8));
  nand2 gate1032(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1033(.a(s_69), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1034(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1035(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1036(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1835(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1836(.a(gate159inter0), .b(s_184), .O(gate159inter1));
  and2  gate1837(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1838(.a(s_184), .O(gate159inter3));
  inv1  gate1839(.a(s_185), .O(gate159inter4));
  nand2 gate1840(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1841(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1842(.a(G444), .O(gate159inter7));
  inv1  gate1843(.a(G531), .O(gate159inter8));
  nand2 gate1844(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1845(.a(s_185), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1846(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1847(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1848(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1541(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1542(.a(gate163inter0), .b(s_142), .O(gate163inter1));
  and2  gate1543(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1544(.a(s_142), .O(gate163inter3));
  inv1  gate1545(.a(s_143), .O(gate163inter4));
  nand2 gate1546(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1547(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1548(.a(G456), .O(gate163inter7));
  inv1  gate1549(.a(G537), .O(gate163inter8));
  nand2 gate1550(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1551(.a(s_143), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1552(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1553(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1554(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate925(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate926(.a(gate170inter0), .b(s_54), .O(gate170inter1));
  and2  gate927(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate928(.a(s_54), .O(gate170inter3));
  inv1  gate929(.a(s_55), .O(gate170inter4));
  nand2 gate930(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate931(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate932(.a(G477), .O(gate170inter7));
  inv1  gate933(.a(G546), .O(gate170inter8));
  nand2 gate934(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate935(.a(s_55), .b(gate170inter3), .O(gate170inter10));
  nor2  gate936(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate937(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate938(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2101(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2102(.a(gate187inter0), .b(s_222), .O(gate187inter1));
  and2  gate2103(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2104(.a(s_222), .O(gate187inter3));
  inv1  gate2105(.a(s_223), .O(gate187inter4));
  nand2 gate2106(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2107(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2108(.a(G574), .O(gate187inter7));
  inv1  gate2109(.a(G575), .O(gate187inter8));
  nand2 gate2110(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2111(.a(s_223), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2112(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2113(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2114(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1793(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1794(.a(gate189inter0), .b(s_178), .O(gate189inter1));
  and2  gate1795(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1796(.a(s_178), .O(gate189inter3));
  inv1  gate1797(.a(s_179), .O(gate189inter4));
  nand2 gate1798(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1799(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1800(.a(G578), .O(gate189inter7));
  inv1  gate1801(.a(G579), .O(gate189inter8));
  nand2 gate1802(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1803(.a(s_179), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1804(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1805(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1806(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1359(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1360(.a(gate207inter0), .b(s_116), .O(gate207inter1));
  and2  gate1361(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1362(.a(s_116), .O(gate207inter3));
  inv1  gate1363(.a(s_117), .O(gate207inter4));
  nand2 gate1364(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1365(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1366(.a(G622), .O(gate207inter7));
  inv1  gate1367(.a(G632), .O(gate207inter8));
  nand2 gate1368(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1369(.a(s_117), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1370(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1371(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1372(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2087(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2088(.a(gate208inter0), .b(s_220), .O(gate208inter1));
  and2  gate2089(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2090(.a(s_220), .O(gate208inter3));
  inv1  gate2091(.a(s_221), .O(gate208inter4));
  nand2 gate2092(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2093(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2094(.a(G627), .O(gate208inter7));
  inv1  gate2095(.a(G637), .O(gate208inter8));
  nand2 gate2096(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2097(.a(s_221), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2098(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2099(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2100(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate967(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate968(.a(gate214inter0), .b(s_60), .O(gate214inter1));
  and2  gate969(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate970(.a(s_60), .O(gate214inter3));
  inv1  gate971(.a(s_61), .O(gate214inter4));
  nand2 gate972(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate973(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate974(.a(G612), .O(gate214inter7));
  inv1  gate975(.a(G672), .O(gate214inter8));
  nand2 gate976(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate977(.a(s_61), .b(gate214inter3), .O(gate214inter10));
  nor2  gate978(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate979(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate980(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1723(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1724(.a(gate215inter0), .b(s_168), .O(gate215inter1));
  and2  gate1725(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1726(.a(s_168), .O(gate215inter3));
  inv1  gate1727(.a(s_169), .O(gate215inter4));
  nand2 gate1728(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1729(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1730(.a(G607), .O(gate215inter7));
  inv1  gate1731(.a(G675), .O(gate215inter8));
  nand2 gate1732(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1733(.a(s_169), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1734(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1735(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1736(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1919(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1920(.a(gate216inter0), .b(s_196), .O(gate216inter1));
  and2  gate1921(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1922(.a(s_196), .O(gate216inter3));
  inv1  gate1923(.a(s_197), .O(gate216inter4));
  nand2 gate1924(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1925(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1926(.a(G617), .O(gate216inter7));
  inv1  gate1927(.a(G675), .O(gate216inter8));
  nand2 gate1928(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1929(.a(s_197), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1930(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1931(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1932(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1779(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1780(.a(gate217inter0), .b(s_176), .O(gate217inter1));
  and2  gate1781(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1782(.a(s_176), .O(gate217inter3));
  inv1  gate1783(.a(s_177), .O(gate217inter4));
  nand2 gate1784(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1785(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1786(.a(G622), .O(gate217inter7));
  inv1  gate1787(.a(G678), .O(gate217inter8));
  nand2 gate1788(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1789(.a(s_177), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1790(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1791(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1792(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate2227(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2228(.a(gate218inter0), .b(s_240), .O(gate218inter1));
  and2  gate2229(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2230(.a(s_240), .O(gate218inter3));
  inv1  gate2231(.a(s_241), .O(gate218inter4));
  nand2 gate2232(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2233(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2234(.a(G627), .O(gate218inter7));
  inv1  gate2235(.a(G678), .O(gate218inter8));
  nand2 gate2236(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2237(.a(s_241), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2238(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2239(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2240(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1317(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1318(.a(gate220inter0), .b(s_110), .O(gate220inter1));
  and2  gate1319(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1320(.a(s_110), .O(gate220inter3));
  inv1  gate1321(.a(s_111), .O(gate220inter4));
  nand2 gate1322(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1323(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1324(.a(G637), .O(gate220inter7));
  inv1  gate1325(.a(G681), .O(gate220inter8));
  nand2 gate1326(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1327(.a(s_111), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1328(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1329(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1330(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1009(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1010(.a(gate221inter0), .b(s_66), .O(gate221inter1));
  and2  gate1011(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1012(.a(s_66), .O(gate221inter3));
  inv1  gate1013(.a(s_67), .O(gate221inter4));
  nand2 gate1014(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1015(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1016(.a(G622), .O(gate221inter7));
  inv1  gate1017(.a(G684), .O(gate221inter8));
  nand2 gate1018(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1019(.a(s_67), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1020(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1021(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1022(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate2241(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2242(.a(gate222inter0), .b(s_242), .O(gate222inter1));
  and2  gate2243(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2244(.a(s_242), .O(gate222inter3));
  inv1  gate2245(.a(s_243), .O(gate222inter4));
  nand2 gate2246(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2247(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2248(.a(G632), .O(gate222inter7));
  inv1  gate2249(.a(G684), .O(gate222inter8));
  nand2 gate2250(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2251(.a(s_243), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2252(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2253(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2254(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1891(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1892(.a(gate227inter0), .b(s_192), .O(gate227inter1));
  and2  gate1893(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1894(.a(s_192), .O(gate227inter3));
  inv1  gate1895(.a(s_193), .O(gate227inter4));
  nand2 gate1896(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1897(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1898(.a(G694), .O(gate227inter7));
  inv1  gate1899(.a(G695), .O(gate227inter8));
  nand2 gate1900(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1901(.a(s_193), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1902(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1903(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1904(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1457(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1458(.a(gate228inter0), .b(s_130), .O(gate228inter1));
  and2  gate1459(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1460(.a(s_130), .O(gate228inter3));
  inv1  gate1461(.a(s_131), .O(gate228inter4));
  nand2 gate1462(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1463(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1464(.a(G696), .O(gate228inter7));
  inv1  gate1465(.a(G697), .O(gate228inter8));
  nand2 gate1466(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1467(.a(s_131), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1468(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1469(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1470(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1303(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1304(.a(gate230inter0), .b(s_108), .O(gate230inter1));
  and2  gate1305(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1306(.a(s_108), .O(gate230inter3));
  inv1  gate1307(.a(s_109), .O(gate230inter4));
  nand2 gate1308(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1309(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1310(.a(G700), .O(gate230inter7));
  inv1  gate1311(.a(G701), .O(gate230inter8));
  nand2 gate1312(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1313(.a(s_109), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1314(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1315(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1316(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1807(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1808(.a(gate233inter0), .b(s_180), .O(gate233inter1));
  and2  gate1809(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1810(.a(s_180), .O(gate233inter3));
  inv1  gate1811(.a(s_181), .O(gate233inter4));
  nand2 gate1812(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1813(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1814(.a(G242), .O(gate233inter7));
  inv1  gate1815(.a(G718), .O(gate233inter8));
  nand2 gate1816(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1817(.a(s_181), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1818(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1819(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1820(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2031(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2032(.a(gate241inter0), .b(s_212), .O(gate241inter1));
  and2  gate2033(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2034(.a(s_212), .O(gate241inter3));
  inv1  gate2035(.a(s_213), .O(gate241inter4));
  nand2 gate2036(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2037(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2038(.a(G242), .O(gate241inter7));
  inv1  gate2039(.a(G730), .O(gate241inter8));
  nand2 gate2040(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2041(.a(s_213), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2042(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2043(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2044(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate869(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate870(.a(gate243inter0), .b(s_46), .O(gate243inter1));
  and2  gate871(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate872(.a(s_46), .O(gate243inter3));
  inv1  gate873(.a(s_47), .O(gate243inter4));
  nand2 gate874(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate875(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate876(.a(G245), .O(gate243inter7));
  inv1  gate877(.a(G733), .O(gate243inter8));
  nand2 gate878(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate879(.a(s_47), .b(gate243inter3), .O(gate243inter10));
  nor2  gate880(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate881(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate882(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate589(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate590(.a(gate245inter0), .b(s_6), .O(gate245inter1));
  and2  gate591(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate592(.a(s_6), .O(gate245inter3));
  inv1  gate593(.a(s_7), .O(gate245inter4));
  nand2 gate594(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate595(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate596(.a(G248), .O(gate245inter7));
  inv1  gate597(.a(G736), .O(gate245inter8));
  nand2 gate598(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate599(.a(s_7), .b(gate245inter3), .O(gate245inter10));
  nor2  gate600(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate601(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate602(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1051(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1052(.a(gate251inter0), .b(s_72), .O(gate251inter1));
  and2  gate1053(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1054(.a(s_72), .O(gate251inter3));
  inv1  gate1055(.a(s_73), .O(gate251inter4));
  nand2 gate1056(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1057(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1058(.a(G257), .O(gate251inter7));
  inv1  gate1059(.a(G745), .O(gate251inter8));
  nand2 gate1060(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1061(.a(s_73), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1062(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1063(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1064(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1821(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1822(.a(gate255inter0), .b(s_182), .O(gate255inter1));
  and2  gate1823(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1824(.a(s_182), .O(gate255inter3));
  inv1  gate1825(.a(s_183), .O(gate255inter4));
  nand2 gate1826(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1827(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1828(.a(G263), .O(gate255inter7));
  inv1  gate1829(.a(G751), .O(gate255inter8));
  nand2 gate1830(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1831(.a(s_183), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1832(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1833(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1834(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1737(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1738(.a(gate266inter0), .b(s_170), .O(gate266inter1));
  and2  gate1739(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1740(.a(s_170), .O(gate266inter3));
  inv1  gate1741(.a(s_171), .O(gate266inter4));
  nand2 gate1742(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1743(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1744(.a(G645), .O(gate266inter7));
  inv1  gate1745(.a(G773), .O(gate266inter8));
  nand2 gate1746(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1747(.a(s_171), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1748(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1749(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1750(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate883(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate884(.a(gate268inter0), .b(s_48), .O(gate268inter1));
  and2  gate885(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate886(.a(s_48), .O(gate268inter3));
  inv1  gate887(.a(s_49), .O(gate268inter4));
  nand2 gate888(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate889(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate890(.a(G651), .O(gate268inter7));
  inv1  gate891(.a(G779), .O(gate268inter8));
  nand2 gate892(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate893(.a(s_49), .b(gate268inter3), .O(gate268inter10));
  nor2  gate894(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate895(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate896(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1149(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1150(.a(gate269inter0), .b(s_86), .O(gate269inter1));
  and2  gate1151(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1152(.a(s_86), .O(gate269inter3));
  inv1  gate1153(.a(s_87), .O(gate269inter4));
  nand2 gate1154(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1155(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1156(.a(G654), .O(gate269inter7));
  inv1  gate1157(.a(G782), .O(gate269inter8));
  nand2 gate1158(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1159(.a(s_87), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1160(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1161(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1162(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2115(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2116(.a(gate271inter0), .b(s_224), .O(gate271inter1));
  and2  gate2117(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2118(.a(s_224), .O(gate271inter3));
  inv1  gate2119(.a(s_225), .O(gate271inter4));
  nand2 gate2120(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2121(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2122(.a(G660), .O(gate271inter7));
  inv1  gate2123(.a(G788), .O(gate271inter8));
  nand2 gate2124(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2125(.a(s_225), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2126(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2127(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2128(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1093(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1094(.a(gate273inter0), .b(s_78), .O(gate273inter1));
  and2  gate1095(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1096(.a(s_78), .O(gate273inter3));
  inv1  gate1097(.a(s_79), .O(gate273inter4));
  nand2 gate1098(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1099(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1100(.a(G642), .O(gate273inter7));
  inv1  gate1101(.a(G794), .O(gate273inter8));
  nand2 gate1102(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1103(.a(s_79), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1104(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1105(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1106(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1947(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1948(.a(gate282inter0), .b(s_200), .O(gate282inter1));
  and2  gate1949(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1950(.a(s_200), .O(gate282inter3));
  inv1  gate1951(.a(s_201), .O(gate282inter4));
  nand2 gate1952(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1953(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1954(.a(G782), .O(gate282inter7));
  inv1  gate1955(.a(G806), .O(gate282inter8));
  nand2 gate1956(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1957(.a(s_201), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1958(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1959(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1960(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1079(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1080(.a(gate291inter0), .b(s_76), .O(gate291inter1));
  and2  gate1081(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1082(.a(s_76), .O(gate291inter3));
  inv1  gate1083(.a(s_77), .O(gate291inter4));
  nand2 gate1084(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1085(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1086(.a(G822), .O(gate291inter7));
  inv1  gate1087(.a(G823), .O(gate291inter8));
  nand2 gate1088(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1089(.a(s_77), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1090(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1091(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1092(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1443(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1444(.a(gate295inter0), .b(s_128), .O(gate295inter1));
  and2  gate1445(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1446(.a(s_128), .O(gate295inter3));
  inv1  gate1447(.a(s_129), .O(gate295inter4));
  nand2 gate1448(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1449(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1450(.a(G830), .O(gate295inter7));
  inv1  gate1451(.a(G831), .O(gate295inter8));
  nand2 gate1452(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1453(.a(s_129), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1454(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1455(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1456(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1037(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1038(.a(gate387inter0), .b(s_70), .O(gate387inter1));
  and2  gate1039(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1040(.a(s_70), .O(gate387inter3));
  inv1  gate1041(.a(s_71), .O(gate387inter4));
  nand2 gate1042(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1043(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1044(.a(G1), .O(gate387inter7));
  inv1  gate1045(.a(G1036), .O(gate387inter8));
  nand2 gate1046(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1047(.a(s_71), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1048(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1049(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1050(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1765(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1766(.a(gate390inter0), .b(s_174), .O(gate390inter1));
  and2  gate1767(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1768(.a(s_174), .O(gate390inter3));
  inv1  gate1769(.a(s_175), .O(gate390inter4));
  nand2 gate1770(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1771(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1772(.a(G4), .O(gate390inter7));
  inv1  gate1773(.a(G1045), .O(gate390inter8));
  nand2 gate1774(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1775(.a(s_175), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1776(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1777(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1778(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1107(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1108(.a(gate395inter0), .b(s_80), .O(gate395inter1));
  and2  gate1109(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1110(.a(s_80), .O(gate395inter3));
  inv1  gate1111(.a(s_81), .O(gate395inter4));
  nand2 gate1112(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1113(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1114(.a(G9), .O(gate395inter7));
  inv1  gate1115(.a(G1060), .O(gate395inter8));
  nand2 gate1116(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1117(.a(s_81), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1118(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1119(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1120(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate743(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate744(.a(gate399inter0), .b(s_28), .O(gate399inter1));
  and2  gate745(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate746(.a(s_28), .O(gate399inter3));
  inv1  gate747(.a(s_29), .O(gate399inter4));
  nand2 gate748(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate749(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate750(.a(G13), .O(gate399inter7));
  inv1  gate751(.a(G1072), .O(gate399inter8));
  nand2 gate752(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate753(.a(s_29), .b(gate399inter3), .O(gate399inter10));
  nor2  gate754(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate755(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate756(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1583(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1584(.a(gate405inter0), .b(s_148), .O(gate405inter1));
  and2  gate1585(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1586(.a(s_148), .O(gate405inter3));
  inv1  gate1587(.a(s_149), .O(gate405inter4));
  nand2 gate1588(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1589(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1590(.a(G19), .O(gate405inter7));
  inv1  gate1591(.a(G1090), .O(gate405inter8));
  nand2 gate1592(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1593(.a(s_149), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1594(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1595(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1596(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2129(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2130(.a(gate408inter0), .b(s_226), .O(gate408inter1));
  and2  gate2131(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2132(.a(s_226), .O(gate408inter3));
  inv1  gate2133(.a(s_227), .O(gate408inter4));
  nand2 gate2134(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2135(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2136(.a(G22), .O(gate408inter7));
  inv1  gate2137(.a(G1099), .O(gate408inter8));
  nand2 gate2138(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2139(.a(s_227), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2140(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2141(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2142(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate757(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate758(.a(gate412inter0), .b(s_30), .O(gate412inter1));
  and2  gate759(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate760(.a(s_30), .O(gate412inter3));
  inv1  gate761(.a(s_31), .O(gate412inter4));
  nand2 gate762(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate763(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate764(.a(G26), .O(gate412inter7));
  inv1  gate765(.a(G1111), .O(gate412inter8));
  nand2 gate766(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate767(.a(s_31), .b(gate412inter3), .O(gate412inter10));
  nor2  gate768(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate769(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate770(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate645(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate646(.a(gate420inter0), .b(s_14), .O(gate420inter1));
  and2  gate647(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate648(.a(s_14), .O(gate420inter3));
  inv1  gate649(.a(s_15), .O(gate420inter4));
  nand2 gate650(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate651(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate652(.a(G1036), .O(gate420inter7));
  inv1  gate653(.a(G1132), .O(gate420inter8));
  nand2 gate654(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate655(.a(s_15), .b(gate420inter3), .O(gate420inter10));
  nor2  gate656(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate657(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate658(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2157(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2158(.a(gate421inter0), .b(s_230), .O(gate421inter1));
  and2  gate2159(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2160(.a(s_230), .O(gate421inter3));
  inv1  gate2161(.a(s_231), .O(gate421inter4));
  nand2 gate2162(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2163(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2164(.a(G2), .O(gate421inter7));
  inv1  gate2165(.a(G1135), .O(gate421inter8));
  nand2 gate2166(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2167(.a(s_231), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2168(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2169(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2170(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate631(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate632(.a(gate422inter0), .b(s_12), .O(gate422inter1));
  and2  gate633(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate634(.a(s_12), .O(gate422inter3));
  inv1  gate635(.a(s_13), .O(gate422inter4));
  nand2 gate636(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate637(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate638(.a(G1039), .O(gate422inter7));
  inv1  gate639(.a(G1135), .O(gate422inter8));
  nand2 gate640(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate641(.a(s_13), .b(gate422inter3), .O(gate422inter10));
  nor2  gate642(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate643(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate644(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate2059(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2060(.a(gate423inter0), .b(s_216), .O(gate423inter1));
  and2  gate2061(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2062(.a(s_216), .O(gate423inter3));
  inv1  gate2063(.a(s_217), .O(gate423inter4));
  nand2 gate2064(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2065(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2066(.a(G3), .O(gate423inter7));
  inv1  gate2067(.a(G1138), .O(gate423inter8));
  nand2 gate2068(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2069(.a(s_217), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2070(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2071(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2072(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1751(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1752(.a(gate424inter0), .b(s_172), .O(gate424inter1));
  and2  gate1753(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1754(.a(s_172), .O(gate424inter3));
  inv1  gate1755(.a(s_173), .O(gate424inter4));
  nand2 gate1756(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1757(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1758(.a(G1042), .O(gate424inter7));
  inv1  gate1759(.a(G1138), .O(gate424inter8));
  nand2 gate1760(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1761(.a(s_173), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1762(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1763(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1764(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1331(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1332(.a(gate425inter0), .b(s_112), .O(gate425inter1));
  and2  gate1333(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1334(.a(s_112), .O(gate425inter3));
  inv1  gate1335(.a(s_113), .O(gate425inter4));
  nand2 gate1336(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1337(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1338(.a(G4), .O(gate425inter7));
  inv1  gate1339(.a(G1141), .O(gate425inter8));
  nand2 gate1340(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1341(.a(s_113), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1342(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1343(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1344(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate701(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate702(.a(gate426inter0), .b(s_22), .O(gate426inter1));
  and2  gate703(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate704(.a(s_22), .O(gate426inter3));
  inv1  gate705(.a(s_23), .O(gate426inter4));
  nand2 gate706(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate707(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate708(.a(G1045), .O(gate426inter7));
  inv1  gate709(.a(G1141), .O(gate426inter8));
  nand2 gate710(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate711(.a(s_23), .b(gate426inter3), .O(gate426inter10));
  nor2  gate712(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate713(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate714(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1961(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1962(.a(gate428inter0), .b(s_202), .O(gate428inter1));
  and2  gate1963(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1964(.a(s_202), .O(gate428inter3));
  inv1  gate1965(.a(s_203), .O(gate428inter4));
  nand2 gate1966(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1967(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1968(.a(G1048), .O(gate428inter7));
  inv1  gate1969(.a(G1144), .O(gate428inter8));
  nand2 gate1970(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1971(.a(s_203), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1972(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1973(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1974(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate687(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate688(.a(gate433inter0), .b(s_20), .O(gate433inter1));
  and2  gate689(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate690(.a(s_20), .O(gate433inter3));
  inv1  gate691(.a(s_21), .O(gate433inter4));
  nand2 gate692(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate693(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate694(.a(G8), .O(gate433inter7));
  inv1  gate695(.a(G1153), .O(gate433inter8));
  nand2 gate696(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate697(.a(s_21), .b(gate433inter3), .O(gate433inter10));
  nor2  gate698(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate699(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate700(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1177(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1178(.a(gate435inter0), .b(s_90), .O(gate435inter1));
  and2  gate1179(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1180(.a(s_90), .O(gate435inter3));
  inv1  gate1181(.a(s_91), .O(gate435inter4));
  nand2 gate1182(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1183(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1184(.a(G9), .O(gate435inter7));
  inv1  gate1185(.a(G1156), .O(gate435inter8));
  nand2 gate1186(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1187(.a(s_91), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1188(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1189(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1190(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1905(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1906(.a(gate439inter0), .b(s_194), .O(gate439inter1));
  and2  gate1907(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1908(.a(s_194), .O(gate439inter3));
  inv1  gate1909(.a(s_195), .O(gate439inter4));
  nand2 gate1910(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1911(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1912(.a(G11), .O(gate439inter7));
  inv1  gate1913(.a(G1162), .O(gate439inter8));
  nand2 gate1914(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1915(.a(s_195), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1916(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1917(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1918(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1163(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1164(.a(gate444inter0), .b(s_88), .O(gate444inter1));
  and2  gate1165(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1166(.a(s_88), .O(gate444inter3));
  inv1  gate1167(.a(s_89), .O(gate444inter4));
  nand2 gate1168(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1169(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1170(.a(G1072), .O(gate444inter7));
  inv1  gate1171(.a(G1168), .O(gate444inter8));
  nand2 gate1172(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1173(.a(s_89), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1174(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1175(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1176(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1471(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1472(.a(gate449inter0), .b(s_132), .O(gate449inter1));
  and2  gate1473(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1474(.a(s_132), .O(gate449inter3));
  inv1  gate1475(.a(s_133), .O(gate449inter4));
  nand2 gate1476(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1477(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1478(.a(G16), .O(gate449inter7));
  inv1  gate1479(.a(G1177), .O(gate449inter8));
  nand2 gate1480(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1481(.a(s_133), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1482(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1483(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1484(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate841(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate842(.a(gate450inter0), .b(s_42), .O(gate450inter1));
  and2  gate843(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate844(.a(s_42), .O(gate450inter3));
  inv1  gate845(.a(s_43), .O(gate450inter4));
  nand2 gate846(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate847(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate848(.a(G1081), .O(gate450inter7));
  inv1  gate849(.a(G1177), .O(gate450inter8));
  nand2 gate850(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate851(.a(s_43), .b(gate450inter3), .O(gate450inter10));
  nor2  gate852(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate853(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate854(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1121(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1122(.a(gate453inter0), .b(s_82), .O(gate453inter1));
  and2  gate1123(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1124(.a(s_82), .O(gate453inter3));
  inv1  gate1125(.a(s_83), .O(gate453inter4));
  nand2 gate1126(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1127(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1128(.a(G18), .O(gate453inter7));
  inv1  gate1129(.a(G1183), .O(gate453inter8));
  nand2 gate1130(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1131(.a(s_83), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1132(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1133(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1134(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate953(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate954(.a(gate454inter0), .b(s_58), .O(gate454inter1));
  and2  gate955(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate956(.a(s_58), .O(gate454inter3));
  inv1  gate957(.a(s_59), .O(gate454inter4));
  nand2 gate958(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate959(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate960(.a(G1087), .O(gate454inter7));
  inv1  gate961(.a(G1183), .O(gate454inter8));
  nand2 gate962(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate963(.a(s_59), .b(gate454inter3), .O(gate454inter10));
  nor2  gate964(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate965(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate966(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate2297(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2298(.a(gate456inter0), .b(s_250), .O(gate456inter1));
  and2  gate2299(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2300(.a(s_250), .O(gate456inter3));
  inv1  gate2301(.a(s_251), .O(gate456inter4));
  nand2 gate2302(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2303(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2304(.a(G1090), .O(gate456inter7));
  inv1  gate2305(.a(G1186), .O(gate456inter8));
  nand2 gate2306(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2307(.a(s_251), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2308(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2309(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2310(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1275(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1276(.a(gate459inter0), .b(s_104), .O(gate459inter1));
  and2  gate1277(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1278(.a(s_104), .O(gate459inter3));
  inv1  gate1279(.a(s_105), .O(gate459inter4));
  nand2 gate1280(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1281(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1282(.a(G21), .O(gate459inter7));
  inv1  gate1283(.a(G1192), .O(gate459inter8));
  nand2 gate1284(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1285(.a(s_105), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1286(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1287(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1288(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1219(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1220(.a(gate463inter0), .b(s_96), .O(gate463inter1));
  and2  gate1221(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1222(.a(s_96), .O(gate463inter3));
  inv1  gate1223(.a(s_97), .O(gate463inter4));
  nand2 gate1224(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1225(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1226(.a(G23), .O(gate463inter7));
  inv1  gate1227(.a(G1198), .O(gate463inter8));
  nand2 gate1228(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1229(.a(s_97), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1230(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1231(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1232(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1975(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1976(.a(gate467inter0), .b(s_204), .O(gate467inter1));
  and2  gate1977(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1978(.a(s_204), .O(gate467inter3));
  inv1  gate1979(.a(s_205), .O(gate467inter4));
  nand2 gate1980(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1981(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1982(.a(G25), .O(gate467inter7));
  inv1  gate1983(.a(G1204), .O(gate467inter8));
  nand2 gate1984(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1985(.a(s_205), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1986(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1987(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1988(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate995(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate996(.a(gate468inter0), .b(s_64), .O(gate468inter1));
  and2  gate997(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate998(.a(s_64), .O(gate468inter3));
  inv1  gate999(.a(s_65), .O(gate468inter4));
  nand2 gate1000(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1001(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1002(.a(G1108), .O(gate468inter7));
  inv1  gate1003(.a(G1204), .O(gate468inter8));
  nand2 gate1004(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1005(.a(s_65), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1006(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1007(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1008(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1989(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1990(.a(gate475inter0), .b(s_206), .O(gate475inter1));
  and2  gate1991(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1992(.a(s_206), .O(gate475inter3));
  inv1  gate1993(.a(s_207), .O(gate475inter4));
  nand2 gate1994(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1995(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1996(.a(G29), .O(gate475inter7));
  inv1  gate1997(.a(G1216), .O(gate475inter8));
  nand2 gate1998(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1999(.a(s_207), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2000(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2001(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2002(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate659(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate660(.a(gate476inter0), .b(s_16), .O(gate476inter1));
  and2  gate661(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate662(.a(s_16), .O(gate476inter3));
  inv1  gate663(.a(s_17), .O(gate476inter4));
  nand2 gate664(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate665(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate666(.a(G1120), .O(gate476inter7));
  inv1  gate667(.a(G1216), .O(gate476inter8));
  nand2 gate668(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate669(.a(s_17), .b(gate476inter3), .O(gate476inter10));
  nor2  gate670(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate671(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate672(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1625(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1626(.a(gate477inter0), .b(s_154), .O(gate477inter1));
  and2  gate1627(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1628(.a(s_154), .O(gate477inter3));
  inv1  gate1629(.a(s_155), .O(gate477inter4));
  nand2 gate1630(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1631(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1632(.a(G30), .O(gate477inter7));
  inv1  gate1633(.a(G1219), .O(gate477inter8));
  nand2 gate1634(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1635(.a(s_155), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1636(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1637(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1638(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2213(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2214(.a(gate479inter0), .b(s_238), .O(gate479inter1));
  and2  gate2215(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2216(.a(s_238), .O(gate479inter3));
  inv1  gate2217(.a(s_239), .O(gate479inter4));
  nand2 gate2218(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2219(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2220(.a(G31), .O(gate479inter7));
  inv1  gate2221(.a(G1222), .O(gate479inter8));
  nand2 gate2222(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2223(.a(s_239), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2224(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2225(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2226(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate547(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate548(.a(gate481inter0), .b(s_0), .O(gate481inter1));
  and2  gate549(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate550(.a(s_0), .O(gate481inter3));
  inv1  gate551(.a(s_1), .O(gate481inter4));
  nand2 gate552(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate553(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate554(.a(G32), .O(gate481inter7));
  inv1  gate555(.a(G1225), .O(gate481inter8));
  nand2 gate556(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate557(.a(s_1), .b(gate481inter3), .O(gate481inter10));
  nor2  gate558(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate559(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate560(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate2003(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2004(.a(gate482inter0), .b(s_208), .O(gate482inter1));
  and2  gate2005(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2006(.a(s_208), .O(gate482inter3));
  inv1  gate2007(.a(s_209), .O(gate482inter4));
  nand2 gate2008(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2009(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2010(.a(G1129), .O(gate482inter7));
  inv1  gate2011(.a(G1225), .O(gate482inter8));
  nand2 gate2012(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2013(.a(s_209), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2014(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2015(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2016(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate771(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate772(.a(gate488inter0), .b(s_32), .O(gate488inter1));
  and2  gate773(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate774(.a(s_32), .O(gate488inter3));
  inv1  gate775(.a(s_33), .O(gate488inter4));
  nand2 gate776(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate777(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate778(.a(G1238), .O(gate488inter7));
  inv1  gate779(.a(G1239), .O(gate488inter8));
  nand2 gate780(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate781(.a(s_33), .b(gate488inter3), .O(gate488inter10));
  nor2  gate782(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate783(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate784(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1653(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1654(.a(gate489inter0), .b(s_158), .O(gate489inter1));
  and2  gate1655(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1656(.a(s_158), .O(gate489inter3));
  inv1  gate1657(.a(s_159), .O(gate489inter4));
  nand2 gate1658(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1659(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1660(.a(G1240), .O(gate489inter7));
  inv1  gate1661(.a(G1241), .O(gate489inter8));
  nand2 gate1662(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1663(.a(s_159), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1664(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1665(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1666(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate575(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate576(.a(gate492inter0), .b(s_4), .O(gate492inter1));
  and2  gate577(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate578(.a(s_4), .O(gate492inter3));
  inv1  gate579(.a(s_5), .O(gate492inter4));
  nand2 gate580(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate581(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate582(.a(G1246), .O(gate492inter7));
  inv1  gate583(.a(G1247), .O(gate492inter8));
  nand2 gate584(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate585(.a(s_5), .b(gate492inter3), .O(gate492inter10));
  nor2  gate586(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate587(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate588(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1849(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1850(.a(gate495inter0), .b(s_186), .O(gate495inter1));
  and2  gate1851(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1852(.a(s_186), .O(gate495inter3));
  inv1  gate1853(.a(s_187), .O(gate495inter4));
  nand2 gate1854(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1855(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1856(.a(G1252), .O(gate495inter7));
  inv1  gate1857(.a(G1253), .O(gate495inter8));
  nand2 gate1858(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1859(.a(s_187), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1860(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1861(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1862(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1933(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1934(.a(gate498inter0), .b(s_198), .O(gate498inter1));
  and2  gate1935(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1936(.a(s_198), .O(gate498inter3));
  inv1  gate1937(.a(s_199), .O(gate498inter4));
  nand2 gate1938(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1939(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1940(.a(G1258), .O(gate498inter7));
  inv1  gate1941(.a(G1259), .O(gate498inter8));
  nand2 gate1942(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1943(.a(s_199), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1944(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1945(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1946(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2269(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2270(.a(gate501inter0), .b(s_246), .O(gate501inter1));
  and2  gate2271(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2272(.a(s_246), .O(gate501inter3));
  inv1  gate2273(.a(s_247), .O(gate501inter4));
  nand2 gate2274(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2275(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2276(.a(G1264), .O(gate501inter7));
  inv1  gate2277(.a(G1265), .O(gate501inter8));
  nand2 gate2278(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2279(.a(s_247), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2280(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2281(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2282(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2045(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2046(.a(gate508inter0), .b(s_214), .O(gate508inter1));
  and2  gate2047(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2048(.a(s_214), .O(gate508inter3));
  inv1  gate2049(.a(s_215), .O(gate508inter4));
  nand2 gate2050(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2051(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2052(.a(G1278), .O(gate508inter7));
  inv1  gate2053(.a(G1279), .O(gate508inter8));
  nand2 gate2054(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2055(.a(s_215), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2056(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2057(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2058(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2171(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2172(.a(gate510inter0), .b(s_232), .O(gate510inter1));
  and2  gate2173(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2174(.a(s_232), .O(gate510inter3));
  inv1  gate2175(.a(s_233), .O(gate510inter4));
  nand2 gate2176(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2177(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2178(.a(G1282), .O(gate510inter7));
  inv1  gate2179(.a(G1283), .O(gate510inter8));
  nand2 gate2180(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2181(.a(s_233), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2182(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2183(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2184(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1569(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1570(.a(gate511inter0), .b(s_146), .O(gate511inter1));
  and2  gate1571(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1572(.a(s_146), .O(gate511inter3));
  inv1  gate1573(.a(s_147), .O(gate511inter4));
  nand2 gate1574(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1575(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1576(.a(G1284), .O(gate511inter7));
  inv1  gate1577(.a(G1285), .O(gate511inter8));
  nand2 gate1578(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1579(.a(s_147), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1580(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1581(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1582(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1247(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1248(.a(gate513inter0), .b(s_100), .O(gate513inter1));
  and2  gate1249(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1250(.a(s_100), .O(gate513inter3));
  inv1  gate1251(.a(s_101), .O(gate513inter4));
  nand2 gate1252(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1253(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1254(.a(G1288), .O(gate513inter7));
  inv1  gate1255(.a(G1289), .O(gate513inter8));
  nand2 gate1256(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1257(.a(s_101), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1258(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1259(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1260(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate2199(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2200(.a(gate514inter0), .b(s_236), .O(gate514inter1));
  and2  gate2201(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2202(.a(s_236), .O(gate514inter3));
  inv1  gate2203(.a(s_237), .O(gate514inter4));
  nand2 gate2204(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2205(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2206(.a(G1290), .O(gate514inter7));
  inv1  gate2207(.a(G1291), .O(gate514inter8));
  nand2 gate2208(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2209(.a(s_237), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2210(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2211(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2212(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule