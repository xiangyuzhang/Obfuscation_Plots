module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2129(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2130(.a(gate9inter0), .b(s_226), .O(gate9inter1));
  and2  gate2131(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2132(.a(s_226), .O(gate9inter3));
  inv1  gate2133(.a(s_227), .O(gate9inter4));
  nand2 gate2134(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2135(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2136(.a(G1), .O(gate9inter7));
  inv1  gate2137(.a(G2), .O(gate9inter8));
  nand2 gate2138(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2139(.a(s_227), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2140(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2141(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2142(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1233(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1234(.a(gate12inter0), .b(s_98), .O(gate12inter1));
  and2  gate1235(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1236(.a(s_98), .O(gate12inter3));
  inv1  gate1237(.a(s_99), .O(gate12inter4));
  nand2 gate1238(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1239(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1240(.a(G7), .O(gate12inter7));
  inv1  gate1241(.a(G8), .O(gate12inter8));
  nand2 gate1242(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1243(.a(s_99), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1244(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1245(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1246(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1191(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1192(.a(gate13inter0), .b(s_92), .O(gate13inter1));
  and2  gate1193(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1194(.a(s_92), .O(gate13inter3));
  inv1  gate1195(.a(s_93), .O(gate13inter4));
  nand2 gate1196(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1197(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1198(.a(G9), .O(gate13inter7));
  inv1  gate1199(.a(G10), .O(gate13inter8));
  nand2 gate1200(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1201(.a(s_93), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1202(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1203(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1204(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate2675(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2676(.a(gate14inter0), .b(s_304), .O(gate14inter1));
  and2  gate2677(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2678(.a(s_304), .O(gate14inter3));
  inv1  gate2679(.a(s_305), .O(gate14inter4));
  nand2 gate2680(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2681(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2682(.a(G11), .O(gate14inter7));
  inv1  gate2683(.a(G12), .O(gate14inter8));
  nand2 gate2684(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2685(.a(s_305), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2686(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2687(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2688(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2017(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2018(.a(gate19inter0), .b(s_210), .O(gate19inter1));
  and2  gate2019(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2020(.a(s_210), .O(gate19inter3));
  inv1  gate2021(.a(s_211), .O(gate19inter4));
  nand2 gate2022(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2023(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2024(.a(G21), .O(gate19inter7));
  inv1  gate2025(.a(G22), .O(gate19inter8));
  nand2 gate2026(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2027(.a(s_211), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2028(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2029(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2030(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1443(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1444(.a(gate20inter0), .b(s_128), .O(gate20inter1));
  and2  gate1445(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1446(.a(s_128), .O(gate20inter3));
  inv1  gate1447(.a(s_129), .O(gate20inter4));
  nand2 gate1448(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1449(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1450(.a(G23), .O(gate20inter7));
  inv1  gate1451(.a(G24), .O(gate20inter8));
  nand2 gate1452(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1453(.a(s_129), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1454(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1455(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1456(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1807(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1808(.a(gate23inter0), .b(s_180), .O(gate23inter1));
  and2  gate1809(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1810(.a(s_180), .O(gate23inter3));
  inv1  gate1811(.a(s_181), .O(gate23inter4));
  nand2 gate1812(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1813(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1814(.a(G29), .O(gate23inter7));
  inv1  gate1815(.a(G30), .O(gate23inter8));
  nand2 gate1816(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1817(.a(s_181), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1818(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1819(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1820(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2619(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2620(.a(gate25inter0), .b(s_296), .O(gate25inter1));
  and2  gate2621(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2622(.a(s_296), .O(gate25inter3));
  inv1  gate2623(.a(s_297), .O(gate25inter4));
  nand2 gate2624(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2625(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2626(.a(G1), .O(gate25inter7));
  inv1  gate2627(.a(G5), .O(gate25inter8));
  nand2 gate2628(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2629(.a(s_297), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2630(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2631(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2632(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate939(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate940(.a(gate31inter0), .b(s_56), .O(gate31inter1));
  and2  gate941(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate942(.a(s_56), .O(gate31inter3));
  inv1  gate943(.a(s_57), .O(gate31inter4));
  nand2 gate944(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate945(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate946(.a(G4), .O(gate31inter7));
  inv1  gate947(.a(G8), .O(gate31inter8));
  nand2 gate948(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate949(.a(s_57), .b(gate31inter3), .O(gate31inter10));
  nor2  gate950(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate951(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate952(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate925(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate926(.a(gate35inter0), .b(s_54), .O(gate35inter1));
  and2  gate927(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate928(.a(s_54), .O(gate35inter3));
  inv1  gate929(.a(s_55), .O(gate35inter4));
  nand2 gate930(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate931(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate932(.a(G18), .O(gate35inter7));
  inv1  gate933(.a(G22), .O(gate35inter8));
  nand2 gate934(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate935(.a(s_55), .b(gate35inter3), .O(gate35inter10));
  nor2  gate936(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate937(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate938(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1485(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1486(.a(gate37inter0), .b(s_134), .O(gate37inter1));
  and2  gate1487(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1488(.a(s_134), .O(gate37inter3));
  inv1  gate1489(.a(s_135), .O(gate37inter4));
  nand2 gate1490(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1491(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1492(.a(G19), .O(gate37inter7));
  inv1  gate1493(.a(G23), .O(gate37inter8));
  nand2 gate1494(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1495(.a(s_135), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1496(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1497(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1498(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate813(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate814(.a(gate40inter0), .b(s_38), .O(gate40inter1));
  and2  gate815(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate816(.a(s_38), .O(gate40inter3));
  inv1  gate817(.a(s_39), .O(gate40inter4));
  nand2 gate818(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate819(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate820(.a(G28), .O(gate40inter7));
  inv1  gate821(.a(G32), .O(gate40inter8));
  nand2 gate822(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate823(.a(s_39), .b(gate40inter3), .O(gate40inter10));
  nor2  gate824(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate825(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate826(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1415(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1416(.a(gate41inter0), .b(s_124), .O(gate41inter1));
  and2  gate1417(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1418(.a(s_124), .O(gate41inter3));
  inv1  gate1419(.a(s_125), .O(gate41inter4));
  nand2 gate1420(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1421(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1422(.a(G1), .O(gate41inter7));
  inv1  gate1423(.a(G266), .O(gate41inter8));
  nand2 gate1424(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1425(.a(s_125), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1426(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1427(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1428(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1513(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1514(.a(gate43inter0), .b(s_138), .O(gate43inter1));
  and2  gate1515(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1516(.a(s_138), .O(gate43inter3));
  inv1  gate1517(.a(s_139), .O(gate43inter4));
  nand2 gate1518(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1519(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1520(.a(G3), .O(gate43inter7));
  inv1  gate1521(.a(G269), .O(gate43inter8));
  nand2 gate1522(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1523(.a(s_139), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1524(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1525(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1526(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate631(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate632(.a(gate44inter0), .b(s_12), .O(gate44inter1));
  and2  gate633(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate634(.a(s_12), .O(gate44inter3));
  inv1  gate635(.a(s_13), .O(gate44inter4));
  nand2 gate636(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate637(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate638(.a(G4), .O(gate44inter7));
  inv1  gate639(.a(G269), .O(gate44inter8));
  nand2 gate640(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate641(.a(s_13), .b(gate44inter3), .O(gate44inter10));
  nor2  gate642(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate643(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate644(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1933(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1934(.a(gate46inter0), .b(s_198), .O(gate46inter1));
  and2  gate1935(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1936(.a(s_198), .O(gate46inter3));
  inv1  gate1937(.a(s_199), .O(gate46inter4));
  nand2 gate1938(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1939(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1940(.a(G6), .O(gate46inter7));
  inv1  gate1941(.a(G272), .O(gate46inter8));
  nand2 gate1942(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1943(.a(s_199), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1944(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1945(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1946(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1989(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1990(.a(gate55inter0), .b(s_206), .O(gate55inter1));
  and2  gate1991(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1992(.a(s_206), .O(gate55inter3));
  inv1  gate1993(.a(s_207), .O(gate55inter4));
  nand2 gate1994(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1995(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1996(.a(G15), .O(gate55inter7));
  inv1  gate1997(.a(G287), .O(gate55inter8));
  nand2 gate1998(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1999(.a(s_207), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2000(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2001(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2002(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1135(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1136(.a(gate57inter0), .b(s_84), .O(gate57inter1));
  and2  gate1137(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1138(.a(s_84), .O(gate57inter3));
  inv1  gate1139(.a(s_85), .O(gate57inter4));
  nand2 gate1140(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1141(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1142(.a(G17), .O(gate57inter7));
  inv1  gate1143(.a(G290), .O(gate57inter8));
  nand2 gate1144(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1145(.a(s_85), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1146(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1147(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1148(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate2059(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2060(.a(gate58inter0), .b(s_216), .O(gate58inter1));
  and2  gate2061(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2062(.a(s_216), .O(gate58inter3));
  inv1  gate2063(.a(s_217), .O(gate58inter4));
  nand2 gate2064(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2065(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2066(.a(G18), .O(gate58inter7));
  inv1  gate2067(.a(G290), .O(gate58inter8));
  nand2 gate2068(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2069(.a(s_217), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2070(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2071(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2072(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate2409(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2410(.a(gate65inter0), .b(s_266), .O(gate65inter1));
  and2  gate2411(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2412(.a(s_266), .O(gate65inter3));
  inv1  gate2413(.a(s_267), .O(gate65inter4));
  nand2 gate2414(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2415(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2416(.a(G25), .O(gate65inter7));
  inv1  gate2417(.a(G302), .O(gate65inter8));
  nand2 gate2418(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2419(.a(s_267), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2420(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2421(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2422(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2661(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2662(.a(gate67inter0), .b(s_302), .O(gate67inter1));
  and2  gate2663(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2664(.a(s_302), .O(gate67inter3));
  inv1  gate2665(.a(s_303), .O(gate67inter4));
  nand2 gate2666(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2667(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2668(.a(G27), .O(gate67inter7));
  inv1  gate2669(.a(G305), .O(gate67inter8));
  nand2 gate2670(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2671(.a(s_303), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2672(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2673(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2674(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate2325(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2326(.a(gate68inter0), .b(s_254), .O(gate68inter1));
  and2  gate2327(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2328(.a(s_254), .O(gate68inter3));
  inv1  gate2329(.a(s_255), .O(gate68inter4));
  nand2 gate2330(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2331(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2332(.a(G28), .O(gate68inter7));
  inv1  gate2333(.a(G305), .O(gate68inter8));
  nand2 gate2334(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2335(.a(s_255), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2336(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2337(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2338(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate687(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate688(.a(gate69inter0), .b(s_20), .O(gate69inter1));
  and2  gate689(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate690(.a(s_20), .O(gate69inter3));
  inv1  gate691(.a(s_21), .O(gate69inter4));
  nand2 gate692(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate693(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate694(.a(G29), .O(gate69inter7));
  inv1  gate695(.a(G308), .O(gate69inter8));
  nand2 gate696(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate697(.a(s_21), .b(gate69inter3), .O(gate69inter10));
  nor2  gate698(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate699(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate700(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2451(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2452(.a(gate70inter0), .b(s_272), .O(gate70inter1));
  and2  gate2453(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2454(.a(s_272), .O(gate70inter3));
  inv1  gate2455(.a(s_273), .O(gate70inter4));
  nand2 gate2456(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2457(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2458(.a(G30), .O(gate70inter7));
  inv1  gate2459(.a(G308), .O(gate70inter8));
  nand2 gate2460(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2461(.a(s_273), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2462(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2463(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2464(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1709(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1710(.a(gate77inter0), .b(s_166), .O(gate77inter1));
  and2  gate1711(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1712(.a(s_166), .O(gate77inter3));
  inv1  gate1713(.a(s_167), .O(gate77inter4));
  nand2 gate1714(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1715(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1716(.a(G2), .O(gate77inter7));
  inv1  gate1717(.a(G320), .O(gate77inter8));
  nand2 gate1718(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1719(.a(s_167), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1720(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1721(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1722(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate967(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate968(.a(gate80inter0), .b(s_60), .O(gate80inter1));
  and2  gate969(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate970(.a(s_60), .O(gate80inter3));
  inv1  gate971(.a(s_61), .O(gate80inter4));
  nand2 gate972(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate973(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate974(.a(G14), .O(gate80inter7));
  inv1  gate975(.a(G323), .O(gate80inter8));
  nand2 gate976(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate977(.a(s_61), .b(gate80inter3), .O(gate80inter10));
  nor2  gate978(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate979(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate980(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1289(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1290(.a(gate85inter0), .b(s_106), .O(gate85inter1));
  and2  gate1291(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1292(.a(s_106), .O(gate85inter3));
  inv1  gate1293(.a(s_107), .O(gate85inter4));
  nand2 gate1294(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1295(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1296(.a(G4), .O(gate85inter7));
  inv1  gate1297(.a(G332), .O(gate85inter8));
  nand2 gate1298(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1299(.a(s_107), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1300(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1301(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1302(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1555(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1556(.a(gate87inter0), .b(s_144), .O(gate87inter1));
  and2  gate1557(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1558(.a(s_144), .O(gate87inter3));
  inv1  gate1559(.a(s_145), .O(gate87inter4));
  nand2 gate1560(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1561(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1562(.a(G12), .O(gate87inter7));
  inv1  gate1563(.a(G335), .O(gate87inter8));
  nand2 gate1564(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1565(.a(s_145), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1566(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1567(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1568(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate2297(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2298(.a(gate88inter0), .b(s_250), .O(gate88inter1));
  and2  gate2299(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2300(.a(s_250), .O(gate88inter3));
  inv1  gate2301(.a(s_251), .O(gate88inter4));
  nand2 gate2302(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2303(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2304(.a(G16), .O(gate88inter7));
  inv1  gate2305(.a(G335), .O(gate88inter8));
  nand2 gate2306(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2307(.a(s_251), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2308(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2309(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2310(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate645(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate646(.a(gate89inter0), .b(s_14), .O(gate89inter1));
  and2  gate647(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate648(.a(s_14), .O(gate89inter3));
  inv1  gate649(.a(s_15), .O(gate89inter4));
  nand2 gate650(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate651(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate652(.a(G17), .O(gate89inter7));
  inv1  gate653(.a(G338), .O(gate89inter8));
  nand2 gate654(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate655(.a(s_15), .b(gate89inter3), .O(gate89inter10));
  nor2  gate656(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate657(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate658(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1527(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1528(.a(gate90inter0), .b(s_140), .O(gate90inter1));
  and2  gate1529(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1530(.a(s_140), .O(gate90inter3));
  inv1  gate1531(.a(s_141), .O(gate90inter4));
  nand2 gate1532(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1533(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1534(.a(G21), .O(gate90inter7));
  inv1  gate1535(.a(G338), .O(gate90inter8));
  nand2 gate1536(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1537(.a(s_141), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1538(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1539(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1540(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1317(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1318(.a(gate94inter0), .b(s_110), .O(gate94inter1));
  and2  gate1319(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1320(.a(s_110), .O(gate94inter3));
  inv1  gate1321(.a(s_111), .O(gate94inter4));
  nand2 gate1322(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1323(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1324(.a(G22), .O(gate94inter7));
  inv1  gate1325(.a(G344), .O(gate94inter8));
  nand2 gate1326(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1327(.a(s_111), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1328(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1329(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1330(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2003(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2004(.a(gate96inter0), .b(s_208), .O(gate96inter1));
  and2  gate2005(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2006(.a(s_208), .O(gate96inter3));
  inv1  gate2007(.a(s_209), .O(gate96inter4));
  nand2 gate2008(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2009(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2010(.a(G30), .O(gate96inter7));
  inv1  gate2011(.a(G347), .O(gate96inter8));
  nand2 gate2012(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2013(.a(s_209), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2014(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2015(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2016(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1863(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1864(.a(gate97inter0), .b(s_188), .O(gate97inter1));
  and2  gate1865(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1866(.a(s_188), .O(gate97inter3));
  inv1  gate1867(.a(s_189), .O(gate97inter4));
  nand2 gate1868(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1869(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1870(.a(G19), .O(gate97inter7));
  inv1  gate1871(.a(G350), .O(gate97inter8));
  nand2 gate1872(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1873(.a(s_189), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1874(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1875(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1876(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2073(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2074(.a(gate99inter0), .b(s_218), .O(gate99inter1));
  and2  gate2075(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2076(.a(s_218), .O(gate99inter3));
  inv1  gate2077(.a(s_219), .O(gate99inter4));
  nand2 gate2078(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2079(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2080(.a(G27), .O(gate99inter7));
  inv1  gate2081(.a(G353), .O(gate99inter8));
  nand2 gate2082(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2083(.a(s_219), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2084(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2085(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2086(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate981(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate982(.a(gate101inter0), .b(s_62), .O(gate101inter1));
  and2  gate983(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate984(.a(s_62), .O(gate101inter3));
  inv1  gate985(.a(s_63), .O(gate101inter4));
  nand2 gate986(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate987(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate988(.a(G20), .O(gate101inter7));
  inv1  gate989(.a(G356), .O(gate101inter8));
  nand2 gate990(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate991(.a(s_63), .b(gate101inter3), .O(gate101inter10));
  nor2  gate992(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate993(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate994(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate547(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate548(.a(gate102inter0), .b(s_0), .O(gate102inter1));
  and2  gate549(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate550(.a(s_0), .O(gate102inter3));
  inv1  gate551(.a(s_1), .O(gate102inter4));
  nand2 gate552(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate553(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate554(.a(G24), .O(gate102inter7));
  inv1  gate555(.a(G356), .O(gate102inter8));
  nand2 gate556(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate557(.a(s_1), .b(gate102inter3), .O(gate102inter10));
  nor2  gate558(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate559(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate560(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate2731(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2732(.a(gate103inter0), .b(s_312), .O(gate103inter1));
  and2  gate2733(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2734(.a(s_312), .O(gate103inter3));
  inv1  gate2735(.a(s_313), .O(gate103inter4));
  nand2 gate2736(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2737(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2738(.a(G28), .O(gate103inter7));
  inv1  gate2739(.a(G359), .O(gate103inter8));
  nand2 gate2740(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2741(.a(s_313), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2742(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2743(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2744(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2367(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2368(.a(gate104inter0), .b(s_260), .O(gate104inter1));
  and2  gate2369(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2370(.a(s_260), .O(gate104inter3));
  inv1  gate2371(.a(s_261), .O(gate104inter4));
  nand2 gate2372(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2373(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2374(.a(G32), .O(gate104inter7));
  inv1  gate2375(.a(G359), .O(gate104inter8));
  nand2 gate2376(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2377(.a(s_261), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2378(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2379(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2380(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1821(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1822(.a(gate105inter0), .b(s_182), .O(gate105inter1));
  and2  gate1823(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1824(.a(s_182), .O(gate105inter3));
  inv1  gate1825(.a(s_183), .O(gate105inter4));
  nand2 gate1826(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1827(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1828(.a(G362), .O(gate105inter7));
  inv1  gate1829(.a(G363), .O(gate105inter8));
  nand2 gate1830(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1831(.a(s_183), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1832(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1833(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1834(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1275(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1276(.a(gate107inter0), .b(s_104), .O(gate107inter1));
  and2  gate1277(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1278(.a(s_104), .O(gate107inter3));
  inv1  gate1279(.a(s_105), .O(gate107inter4));
  nand2 gate1280(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1281(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1282(.a(G366), .O(gate107inter7));
  inv1  gate1283(.a(G367), .O(gate107inter8));
  nand2 gate1284(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1285(.a(s_105), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1286(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1287(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1288(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate2269(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2270(.a(gate108inter0), .b(s_246), .O(gate108inter1));
  and2  gate2271(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2272(.a(s_246), .O(gate108inter3));
  inv1  gate2273(.a(s_247), .O(gate108inter4));
  nand2 gate2274(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2275(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2276(.a(G368), .O(gate108inter7));
  inv1  gate2277(.a(G369), .O(gate108inter8));
  nand2 gate2278(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2279(.a(s_247), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2280(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2281(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2282(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate953(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate954(.a(gate110inter0), .b(s_58), .O(gate110inter1));
  and2  gate955(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate956(.a(s_58), .O(gate110inter3));
  inv1  gate957(.a(s_59), .O(gate110inter4));
  nand2 gate958(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate959(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate960(.a(G372), .O(gate110inter7));
  inv1  gate961(.a(G373), .O(gate110inter8));
  nand2 gate962(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate963(.a(s_59), .b(gate110inter3), .O(gate110inter10));
  nor2  gate964(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate965(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate966(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate799(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate800(.a(gate117inter0), .b(s_36), .O(gate117inter1));
  and2  gate801(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate802(.a(s_36), .O(gate117inter3));
  inv1  gate803(.a(s_37), .O(gate117inter4));
  nand2 gate804(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate805(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate806(.a(G386), .O(gate117inter7));
  inv1  gate807(.a(G387), .O(gate117inter8));
  nand2 gate808(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate809(.a(s_37), .b(gate117inter3), .O(gate117inter10));
  nor2  gate810(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate811(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate812(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate897(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate898(.a(gate119inter0), .b(s_50), .O(gate119inter1));
  and2  gate899(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate900(.a(s_50), .O(gate119inter3));
  inv1  gate901(.a(s_51), .O(gate119inter4));
  nand2 gate902(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate903(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate904(.a(G390), .O(gate119inter7));
  inv1  gate905(.a(G391), .O(gate119inter8));
  nand2 gate906(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate907(.a(s_51), .b(gate119inter3), .O(gate119inter10));
  nor2  gate908(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate909(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate910(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate841(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate842(.a(gate120inter0), .b(s_42), .O(gate120inter1));
  and2  gate843(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate844(.a(s_42), .O(gate120inter3));
  inv1  gate845(.a(s_43), .O(gate120inter4));
  nand2 gate846(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate847(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate848(.a(G392), .O(gate120inter7));
  inv1  gate849(.a(G393), .O(gate120inter8));
  nand2 gate850(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate851(.a(s_43), .b(gate120inter3), .O(gate120inter10));
  nor2  gate852(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate853(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate854(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1093(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1094(.a(gate126inter0), .b(s_78), .O(gate126inter1));
  and2  gate1095(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1096(.a(s_78), .O(gate126inter3));
  inv1  gate1097(.a(s_79), .O(gate126inter4));
  nand2 gate1098(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1099(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1100(.a(G404), .O(gate126inter7));
  inv1  gate1101(.a(G405), .O(gate126inter8));
  nand2 gate1102(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1103(.a(s_79), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1104(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1105(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1106(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2087(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2088(.a(gate129inter0), .b(s_220), .O(gate129inter1));
  and2  gate2089(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2090(.a(s_220), .O(gate129inter3));
  inv1  gate2091(.a(s_221), .O(gate129inter4));
  nand2 gate2092(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2093(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2094(.a(G410), .O(gate129inter7));
  inv1  gate2095(.a(G411), .O(gate129inter8));
  nand2 gate2096(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2097(.a(s_221), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2098(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2099(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2100(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1107(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1108(.a(gate133inter0), .b(s_80), .O(gate133inter1));
  and2  gate1109(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1110(.a(s_80), .O(gate133inter3));
  inv1  gate1111(.a(s_81), .O(gate133inter4));
  nand2 gate1112(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1113(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1114(.a(G418), .O(gate133inter7));
  inv1  gate1115(.a(G419), .O(gate133inter8));
  nand2 gate1116(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1117(.a(s_81), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1118(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1119(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1120(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1765(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1766(.a(gate134inter0), .b(s_174), .O(gate134inter1));
  and2  gate1767(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1768(.a(s_174), .O(gate134inter3));
  inv1  gate1769(.a(s_175), .O(gate134inter4));
  nand2 gate1770(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1771(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1772(.a(G420), .O(gate134inter7));
  inv1  gate1773(.a(G421), .O(gate134inter8));
  nand2 gate1774(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1775(.a(s_175), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1776(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1777(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1778(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate673(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate674(.a(gate139inter0), .b(s_18), .O(gate139inter1));
  and2  gate675(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate676(.a(s_18), .O(gate139inter3));
  inv1  gate677(.a(s_19), .O(gate139inter4));
  nand2 gate678(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate679(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate680(.a(G438), .O(gate139inter7));
  inv1  gate681(.a(G441), .O(gate139inter8));
  nand2 gate682(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate683(.a(s_19), .b(gate139inter3), .O(gate139inter10));
  nor2  gate684(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate685(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate686(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1163(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1164(.a(gate140inter0), .b(s_88), .O(gate140inter1));
  and2  gate1165(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1166(.a(s_88), .O(gate140inter3));
  inv1  gate1167(.a(s_89), .O(gate140inter4));
  nand2 gate1168(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1169(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1170(.a(G444), .O(gate140inter7));
  inv1  gate1171(.a(G447), .O(gate140inter8));
  nand2 gate1172(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1173(.a(s_89), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1174(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1175(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1176(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1121(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1122(.a(gate143inter0), .b(s_82), .O(gate143inter1));
  and2  gate1123(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1124(.a(s_82), .O(gate143inter3));
  inv1  gate1125(.a(s_83), .O(gate143inter4));
  nand2 gate1126(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1127(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1128(.a(G462), .O(gate143inter7));
  inv1  gate1129(.a(G465), .O(gate143inter8));
  nand2 gate1130(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1131(.a(s_83), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1132(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1133(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1134(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate855(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate856(.a(gate146inter0), .b(s_44), .O(gate146inter1));
  and2  gate857(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate858(.a(s_44), .O(gate146inter3));
  inv1  gate859(.a(s_45), .O(gate146inter4));
  nand2 gate860(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate861(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate862(.a(G480), .O(gate146inter7));
  inv1  gate863(.a(G483), .O(gate146inter8));
  nand2 gate864(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate865(.a(s_45), .b(gate146inter3), .O(gate146inter10));
  nor2  gate866(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate867(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate868(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2759(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2760(.a(gate148inter0), .b(s_316), .O(gate148inter1));
  and2  gate2761(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2762(.a(s_316), .O(gate148inter3));
  inv1  gate2763(.a(s_317), .O(gate148inter4));
  nand2 gate2764(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2765(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2766(.a(G492), .O(gate148inter7));
  inv1  gate2767(.a(G495), .O(gate148inter8));
  nand2 gate2768(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2769(.a(s_317), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2770(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2771(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2772(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2437(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2438(.a(gate151inter0), .b(s_270), .O(gate151inter1));
  and2  gate2439(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2440(.a(s_270), .O(gate151inter3));
  inv1  gate2441(.a(s_271), .O(gate151inter4));
  nand2 gate2442(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2443(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2444(.a(G510), .O(gate151inter7));
  inv1  gate2445(.a(G513), .O(gate151inter8));
  nand2 gate2446(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2447(.a(s_271), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2448(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2449(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2450(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate729(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate730(.a(gate152inter0), .b(s_26), .O(gate152inter1));
  and2  gate731(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate732(.a(s_26), .O(gate152inter3));
  inv1  gate733(.a(s_27), .O(gate152inter4));
  nand2 gate734(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate735(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate736(.a(G516), .O(gate152inter7));
  inv1  gate737(.a(G519), .O(gate152inter8));
  nand2 gate738(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate739(.a(s_27), .b(gate152inter3), .O(gate152inter10));
  nor2  gate740(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate741(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate742(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate1583(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1584(.a(gate153inter0), .b(s_148), .O(gate153inter1));
  and2  gate1585(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1586(.a(s_148), .O(gate153inter3));
  inv1  gate1587(.a(s_149), .O(gate153inter4));
  nand2 gate1588(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1589(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1590(.a(G426), .O(gate153inter7));
  inv1  gate1591(.a(G522), .O(gate153inter8));
  nand2 gate1592(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1593(.a(s_149), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1594(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1595(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1596(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1639(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1640(.a(gate156inter0), .b(s_156), .O(gate156inter1));
  and2  gate1641(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1642(.a(s_156), .O(gate156inter3));
  inv1  gate1643(.a(s_157), .O(gate156inter4));
  nand2 gate1644(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1645(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1646(.a(G435), .O(gate156inter7));
  inv1  gate1647(.a(G525), .O(gate156inter8));
  nand2 gate1648(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1649(.a(s_157), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1650(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1651(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1652(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate561(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate562(.a(gate157inter0), .b(s_2), .O(gate157inter1));
  and2  gate563(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate564(.a(s_2), .O(gate157inter3));
  inv1  gate565(.a(s_3), .O(gate157inter4));
  nand2 gate566(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate567(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate568(.a(G438), .O(gate157inter7));
  inv1  gate569(.a(G528), .O(gate157inter8));
  nand2 gate570(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate571(.a(s_3), .b(gate157inter3), .O(gate157inter10));
  nor2  gate572(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate573(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate574(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1597(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1598(.a(gate163inter0), .b(s_150), .O(gate163inter1));
  and2  gate1599(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1600(.a(s_150), .O(gate163inter3));
  inv1  gate1601(.a(s_151), .O(gate163inter4));
  nand2 gate1602(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1603(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1604(.a(G456), .O(gate163inter7));
  inv1  gate1605(.a(G537), .O(gate163inter8));
  nand2 gate1606(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1607(.a(s_151), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1608(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1609(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1610(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate1779(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1780(.a(gate164inter0), .b(s_176), .O(gate164inter1));
  and2  gate1781(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1782(.a(s_176), .O(gate164inter3));
  inv1  gate1783(.a(s_177), .O(gate164inter4));
  nand2 gate1784(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1785(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1786(.a(G459), .O(gate164inter7));
  inv1  gate1787(.a(G537), .O(gate164inter8));
  nand2 gate1788(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1789(.a(s_177), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1790(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1791(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1792(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2745(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2746(.a(gate166inter0), .b(s_314), .O(gate166inter1));
  and2  gate2747(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2748(.a(s_314), .O(gate166inter3));
  inv1  gate2749(.a(s_315), .O(gate166inter4));
  nand2 gate2750(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2751(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2752(.a(G465), .O(gate166inter7));
  inv1  gate2753(.a(G540), .O(gate166inter8));
  nand2 gate2754(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2755(.a(s_315), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2756(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2757(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2758(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1247(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1248(.a(gate167inter0), .b(s_100), .O(gate167inter1));
  and2  gate1249(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1250(.a(s_100), .O(gate167inter3));
  inv1  gate1251(.a(s_101), .O(gate167inter4));
  nand2 gate1252(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1253(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1254(.a(G468), .O(gate167inter7));
  inv1  gate1255(.a(G543), .O(gate167inter8));
  nand2 gate1256(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1257(.a(s_101), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1258(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1259(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1260(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2563(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2564(.a(gate170inter0), .b(s_288), .O(gate170inter1));
  and2  gate2565(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2566(.a(s_288), .O(gate170inter3));
  inv1  gate2567(.a(s_289), .O(gate170inter4));
  nand2 gate2568(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2569(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2570(.a(G477), .O(gate170inter7));
  inv1  gate2571(.a(G546), .O(gate170inter8));
  nand2 gate2572(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2573(.a(s_289), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2574(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2575(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2576(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1373(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1374(.a(gate172inter0), .b(s_118), .O(gate172inter1));
  and2  gate1375(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1376(.a(s_118), .O(gate172inter3));
  inv1  gate1377(.a(s_119), .O(gate172inter4));
  nand2 gate1378(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1379(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1380(.a(G483), .O(gate172inter7));
  inv1  gate1381(.a(G549), .O(gate172inter8));
  nand2 gate1382(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1383(.a(s_119), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1384(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1385(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1386(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2787(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2788(.a(gate173inter0), .b(s_320), .O(gate173inter1));
  and2  gate2789(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2790(.a(s_320), .O(gate173inter3));
  inv1  gate2791(.a(s_321), .O(gate173inter4));
  nand2 gate2792(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2793(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2794(.a(G486), .O(gate173inter7));
  inv1  gate2795(.a(G552), .O(gate173inter8));
  nand2 gate2796(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2797(.a(s_321), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2798(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2799(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2800(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate715(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate716(.a(gate174inter0), .b(s_24), .O(gate174inter1));
  and2  gate717(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate718(.a(s_24), .O(gate174inter3));
  inv1  gate719(.a(s_25), .O(gate174inter4));
  nand2 gate720(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate721(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate722(.a(G489), .O(gate174inter7));
  inv1  gate723(.a(G552), .O(gate174inter8));
  nand2 gate724(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate725(.a(s_25), .b(gate174inter3), .O(gate174inter10));
  nor2  gate726(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate727(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate728(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate743(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate744(.a(gate178inter0), .b(s_28), .O(gate178inter1));
  and2  gate745(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate746(.a(s_28), .O(gate178inter3));
  inv1  gate747(.a(s_29), .O(gate178inter4));
  nand2 gate748(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate749(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate750(.a(G501), .O(gate178inter7));
  inv1  gate751(.a(G558), .O(gate178inter8));
  nand2 gate752(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate753(.a(s_29), .b(gate178inter3), .O(gate178inter10));
  nor2  gate754(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate755(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate756(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1681(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1682(.a(gate180inter0), .b(s_162), .O(gate180inter1));
  and2  gate1683(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1684(.a(s_162), .O(gate180inter3));
  inv1  gate1685(.a(s_163), .O(gate180inter4));
  nand2 gate1686(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1687(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1688(.a(G507), .O(gate180inter7));
  inv1  gate1689(.a(G561), .O(gate180inter8));
  nand2 gate1690(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1691(.a(s_163), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1692(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1693(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1694(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2031(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2032(.a(gate182inter0), .b(s_212), .O(gate182inter1));
  and2  gate2033(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2034(.a(s_212), .O(gate182inter3));
  inv1  gate2035(.a(s_213), .O(gate182inter4));
  nand2 gate2036(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2037(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2038(.a(G513), .O(gate182inter7));
  inv1  gate2039(.a(G564), .O(gate182inter8));
  nand2 gate2040(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2041(.a(s_213), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2042(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2043(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2044(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2227(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2228(.a(gate185inter0), .b(s_240), .O(gate185inter1));
  and2  gate2229(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2230(.a(s_240), .O(gate185inter3));
  inv1  gate2231(.a(s_241), .O(gate185inter4));
  nand2 gate2232(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2233(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2234(.a(G570), .O(gate185inter7));
  inv1  gate2235(.a(G571), .O(gate185inter8));
  nand2 gate2236(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2237(.a(s_241), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2238(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2239(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2240(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2199(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2200(.a(gate186inter0), .b(s_236), .O(gate186inter1));
  and2  gate2201(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2202(.a(s_236), .O(gate186inter3));
  inv1  gate2203(.a(s_237), .O(gate186inter4));
  nand2 gate2204(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2205(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2206(.a(G572), .O(gate186inter7));
  inv1  gate2207(.a(G573), .O(gate186inter8));
  nand2 gate2208(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2209(.a(s_237), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2210(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2211(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2212(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate617(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate618(.a(gate196inter0), .b(s_10), .O(gate196inter1));
  and2  gate619(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate620(.a(s_10), .O(gate196inter3));
  inv1  gate621(.a(s_11), .O(gate196inter4));
  nand2 gate622(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate623(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate624(.a(G592), .O(gate196inter7));
  inv1  gate625(.a(G593), .O(gate196inter8));
  nand2 gate626(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate627(.a(s_11), .b(gate196inter3), .O(gate196inter10));
  nor2  gate628(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate629(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate630(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate2465(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2466(.a(gate202inter0), .b(s_274), .O(gate202inter1));
  and2  gate2467(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2468(.a(s_274), .O(gate202inter3));
  inv1  gate2469(.a(s_275), .O(gate202inter4));
  nand2 gate2470(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2471(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2472(.a(G612), .O(gate202inter7));
  inv1  gate2473(.a(G617), .O(gate202inter8));
  nand2 gate2474(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2475(.a(s_275), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2476(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2477(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2478(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1303(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1304(.a(gate206inter0), .b(s_108), .O(gate206inter1));
  and2  gate1305(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1306(.a(s_108), .O(gate206inter3));
  inv1  gate1307(.a(s_109), .O(gate206inter4));
  nand2 gate1308(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1309(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1310(.a(G632), .O(gate206inter7));
  inv1  gate1311(.a(G637), .O(gate206inter8));
  nand2 gate1312(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1313(.a(s_109), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1314(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1315(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1316(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate757(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate758(.a(gate210inter0), .b(s_30), .O(gate210inter1));
  and2  gate759(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate760(.a(s_30), .O(gate210inter3));
  inv1  gate761(.a(s_31), .O(gate210inter4));
  nand2 gate762(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate763(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate764(.a(G607), .O(gate210inter7));
  inv1  gate765(.a(G666), .O(gate210inter8));
  nand2 gate766(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate767(.a(s_31), .b(gate210inter3), .O(gate210inter10));
  nor2  gate768(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate769(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate770(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1737(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1738(.a(gate211inter0), .b(s_170), .O(gate211inter1));
  and2  gate1739(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1740(.a(s_170), .O(gate211inter3));
  inv1  gate1741(.a(s_171), .O(gate211inter4));
  nand2 gate1742(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1743(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1744(.a(G612), .O(gate211inter7));
  inv1  gate1745(.a(G669), .O(gate211inter8));
  nand2 gate1746(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1747(.a(s_171), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1748(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1749(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1750(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1009(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1010(.a(gate212inter0), .b(s_66), .O(gate212inter1));
  and2  gate1011(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1012(.a(s_66), .O(gate212inter3));
  inv1  gate1013(.a(s_67), .O(gate212inter4));
  nand2 gate1014(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1015(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1016(.a(G617), .O(gate212inter7));
  inv1  gate1017(.a(G669), .O(gate212inter8));
  nand2 gate1018(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1019(.a(s_67), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1020(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1021(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1022(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2703(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2704(.a(gate214inter0), .b(s_308), .O(gate214inter1));
  and2  gate2705(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2706(.a(s_308), .O(gate214inter3));
  inv1  gate2707(.a(s_309), .O(gate214inter4));
  nand2 gate2708(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2709(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2710(.a(G612), .O(gate214inter7));
  inv1  gate2711(.a(G672), .O(gate214inter8));
  nand2 gate2712(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2713(.a(s_309), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2714(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2715(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2716(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2633(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2634(.a(gate215inter0), .b(s_298), .O(gate215inter1));
  and2  gate2635(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2636(.a(s_298), .O(gate215inter3));
  inv1  gate2637(.a(s_299), .O(gate215inter4));
  nand2 gate2638(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2639(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2640(.a(G607), .O(gate215inter7));
  inv1  gate2641(.a(G675), .O(gate215inter8));
  nand2 gate2642(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2643(.a(s_299), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2644(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2645(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2646(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate2045(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2046(.a(gate216inter0), .b(s_214), .O(gate216inter1));
  and2  gate2047(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2048(.a(s_214), .O(gate216inter3));
  inv1  gate2049(.a(s_215), .O(gate216inter4));
  nand2 gate2050(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2051(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2052(.a(G617), .O(gate216inter7));
  inv1  gate2053(.a(G675), .O(gate216inter8));
  nand2 gate2054(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2055(.a(s_215), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2056(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2057(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2058(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate575(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate576(.a(gate218inter0), .b(s_4), .O(gate218inter1));
  and2  gate577(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate578(.a(s_4), .O(gate218inter3));
  inv1  gate579(.a(s_5), .O(gate218inter4));
  nand2 gate580(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate581(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate582(.a(G627), .O(gate218inter7));
  inv1  gate583(.a(G678), .O(gate218inter8));
  nand2 gate584(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate585(.a(s_5), .b(gate218inter3), .O(gate218inter10));
  nor2  gate586(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate587(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate588(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1877(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1878(.a(gate221inter0), .b(s_190), .O(gate221inter1));
  and2  gate1879(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1880(.a(s_190), .O(gate221inter3));
  inv1  gate1881(.a(s_191), .O(gate221inter4));
  nand2 gate1882(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1883(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1884(.a(G622), .O(gate221inter7));
  inv1  gate1885(.a(G684), .O(gate221inter8));
  nand2 gate1886(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1887(.a(s_191), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1888(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1889(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1890(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate771(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate772(.a(gate225inter0), .b(s_32), .O(gate225inter1));
  and2  gate773(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate774(.a(s_32), .O(gate225inter3));
  inv1  gate775(.a(s_33), .O(gate225inter4));
  nand2 gate776(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate777(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate778(.a(G690), .O(gate225inter7));
  inv1  gate779(.a(G691), .O(gate225inter8));
  nand2 gate780(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate781(.a(s_33), .b(gate225inter3), .O(gate225inter10));
  nor2  gate782(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate783(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate784(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate589(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate590(.a(gate226inter0), .b(s_6), .O(gate226inter1));
  and2  gate591(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate592(.a(s_6), .O(gate226inter3));
  inv1  gate593(.a(s_7), .O(gate226inter4));
  nand2 gate594(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate595(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate596(.a(G692), .O(gate226inter7));
  inv1  gate597(.a(G693), .O(gate226inter8));
  nand2 gate598(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate599(.a(s_7), .b(gate226inter3), .O(gate226inter10));
  nor2  gate600(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate601(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate602(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1079(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1080(.a(gate234inter0), .b(s_76), .O(gate234inter1));
  and2  gate1081(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1082(.a(s_76), .O(gate234inter3));
  inv1  gate1083(.a(s_77), .O(gate234inter4));
  nand2 gate1084(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1085(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1086(.a(G245), .O(gate234inter7));
  inv1  gate1087(.a(G721), .O(gate234inter8));
  nand2 gate1088(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1089(.a(s_77), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1090(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1091(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1092(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1919(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1920(.a(gate235inter0), .b(s_196), .O(gate235inter1));
  and2  gate1921(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1922(.a(s_196), .O(gate235inter3));
  inv1  gate1923(.a(s_197), .O(gate235inter4));
  nand2 gate1924(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1925(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1926(.a(G248), .O(gate235inter7));
  inv1  gate1927(.a(G724), .O(gate235inter8));
  nand2 gate1928(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1929(.a(s_197), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1930(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1931(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1932(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2353(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2354(.a(gate236inter0), .b(s_258), .O(gate236inter1));
  and2  gate2355(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2356(.a(s_258), .O(gate236inter3));
  inv1  gate2357(.a(s_259), .O(gate236inter4));
  nand2 gate2358(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2359(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2360(.a(G251), .O(gate236inter7));
  inv1  gate2361(.a(G727), .O(gate236inter8));
  nand2 gate2362(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2363(.a(s_259), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2364(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2365(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2366(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1387(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1388(.a(gate237inter0), .b(s_120), .O(gate237inter1));
  and2  gate1389(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1390(.a(s_120), .O(gate237inter3));
  inv1  gate1391(.a(s_121), .O(gate237inter4));
  nand2 gate1392(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1393(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1394(.a(G254), .O(gate237inter7));
  inv1  gate1395(.a(G706), .O(gate237inter8));
  nand2 gate1396(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1397(.a(s_121), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1398(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1399(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1400(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1653(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1654(.a(gate243inter0), .b(s_158), .O(gate243inter1));
  and2  gate1655(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1656(.a(s_158), .O(gate243inter3));
  inv1  gate1657(.a(s_159), .O(gate243inter4));
  nand2 gate1658(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1659(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1660(.a(G245), .O(gate243inter7));
  inv1  gate1661(.a(G733), .O(gate243inter8));
  nand2 gate1662(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1663(.a(s_159), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1664(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1665(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1666(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2381(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2382(.a(gate245inter0), .b(s_262), .O(gate245inter1));
  and2  gate2383(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2384(.a(s_262), .O(gate245inter3));
  inv1  gate2385(.a(s_263), .O(gate245inter4));
  nand2 gate2386(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2387(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2388(.a(G248), .O(gate245inter7));
  inv1  gate2389(.a(G736), .O(gate245inter8));
  nand2 gate2390(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2391(.a(s_263), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2392(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2393(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2394(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1569(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1570(.a(gate247inter0), .b(s_146), .O(gate247inter1));
  and2  gate1571(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1572(.a(s_146), .O(gate247inter3));
  inv1  gate1573(.a(s_147), .O(gate247inter4));
  nand2 gate1574(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1575(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1576(.a(G251), .O(gate247inter7));
  inv1  gate1577(.a(G739), .O(gate247inter8));
  nand2 gate1578(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1579(.a(s_147), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1580(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1581(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1582(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2605(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2606(.a(gate250inter0), .b(s_294), .O(gate250inter1));
  and2  gate2607(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2608(.a(s_294), .O(gate250inter3));
  inv1  gate2609(.a(s_295), .O(gate250inter4));
  nand2 gate2610(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2611(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2612(.a(G706), .O(gate250inter7));
  inv1  gate2613(.a(G742), .O(gate250inter8));
  nand2 gate2614(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2615(.a(s_295), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2616(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2617(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2618(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2283(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2284(.a(gate254inter0), .b(s_248), .O(gate254inter1));
  and2  gate2285(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2286(.a(s_248), .O(gate254inter3));
  inv1  gate2287(.a(s_249), .O(gate254inter4));
  nand2 gate2288(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2289(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2290(.a(G712), .O(gate254inter7));
  inv1  gate2291(.a(G748), .O(gate254inter8));
  nand2 gate2292(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2293(.a(s_249), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2294(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2295(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2296(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1611(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1612(.a(gate256inter0), .b(s_152), .O(gate256inter1));
  and2  gate1613(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1614(.a(s_152), .O(gate256inter3));
  inv1  gate1615(.a(s_153), .O(gate256inter4));
  nand2 gate1616(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1617(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1618(.a(G715), .O(gate256inter7));
  inv1  gate1619(.a(G751), .O(gate256inter8));
  nand2 gate1620(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1621(.a(s_153), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1622(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1623(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1624(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1345(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1346(.a(gate258inter0), .b(s_114), .O(gate258inter1));
  and2  gate1347(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1348(.a(s_114), .O(gate258inter3));
  inv1  gate1349(.a(s_115), .O(gate258inter4));
  nand2 gate1350(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1351(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1352(.a(G756), .O(gate258inter7));
  inv1  gate1353(.a(G757), .O(gate258inter8));
  nand2 gate1354(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1355(.a(s_115), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1356(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1357(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1358(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1429(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1430(.a(gate262inter0), .b(s_126), .O(gate262inter1));
  and2  gate1431(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1432(.a(s_126), .O(gate262inter3));
  inv1  gate1433(.a(s_127), .O(gate262inter4));
  nand2 gate1434(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1435(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1436(.a(G764), .O(gate262inter7));
  inv1  gate1437(.a(G765), .O(gate262inter8));
  nand2 gate1438(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1439(.a(s_127), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1440(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1441(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1442(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1975(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1976(.a(gate265inter0), .b(s_204), .O(gate265inter1));
  and2  gate1977(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1978(.a(s_204), .O(gate265inter3));
  inv1  gate1979(.a(s_205), .O(gate265inter4));
  nand2 gate1980(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1981(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1982(.a(G642), .O(gate265inter7));
  inv1  gate1983(.a(G770), .O(gate265inter8));
  nand2 gate1984(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1985(.a(s_205), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1986(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1987(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1988(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1667(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1668(.a(gate267inter0), .b(s_160), .O(gate267inter1));
  and2  gate1669(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1670(.a(s_160), .O(gate267inter3));
  inv1  gate1671(.a(s_161), .O(gate267inter4));
  nand2 gate1672(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1673(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1674(.a(G648), .O(gate267inter7));
  inv1  gate1675(.a(G776), .O(gate267inter8));
  nand2 gate1676(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1677(.a(s_161), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1678(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1679(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1680(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2171(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2172(.a(gate268inter0), .b(s_232), .O(gate268inter1));
  and2  gate2173(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2174(.a(s_232), .O(gate268inter3));
  inv1  gate2175(.a(s_233), .O(gate268inter4));
  nand2 gate2176(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2177(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2178(.a(G651), .O(gate268inter7));
  inv1  gate2179(.a(G779), .O(gate268inter8));
  nand2 gate2180(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2181(.a(s_233), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2182(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2183(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2184(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2507(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2508(.a(gate272inter0), .b(s_280), .O(gate272inter1));
  and2  gate2509(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2510(.a(s_280), .O(gate272inter3));
  inv1  gate2511(.a(s_281), .O(gate272inter4));
  nand2 gate2512(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2513(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2514(.a(G663), .O(gate272inter7));
  inv1  gate2515(.a(G791), .O(gate272inter8));
  nand2 gate2516(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2517(.a(s_281), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2518(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2519(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2520(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1065(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1066(.a(gate278inter0), .b(s_74), .O(gate278inter1));
  and2  gate1067(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1068(.a(s_74), .O(gate278inter3));
  inv1  gate1069(.a(s_75), .O(gate278inter4));
  nand2 gate1070(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1071(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1072(.a(G776), .O(gate278inter7));
  inv1  gate1073(.a(G800), .O(gate278inter8));
  nand2 gate1074(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1075(.a(s_75), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1076(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1077(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1078(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2255(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2256(.a(gate282inter0), .b(s_244), .O(gate282inter1));
  and2  gate2257(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2258(.a(s_244), .O(gate282inter3));
  inv1  gate2259(.a(s_245), .O(gate282inter4));
  nand2 gate2260(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2261(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2262(.a(G782), .O(gate282inter7));
  inv1  gate2263(.a(G806), .O(gate282inter8));
  nand2 gate2264(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2265(.a(s_245), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2266(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2267(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2268(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2101(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2102(.a(gate285inter0), .b(s_222), .O(gate285inter1));
  and2  gate2103(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2104(.a(s_222), .O(gate285inter3));
  inv1  gate2105(.a(s_223), .O(gate285inter4));
  nand2 gate2106(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2107(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2108(.a(G660), .O(gate285inter7));
  inv1  gate2109(.a(G812), .O(gate285inter8));
  nand2 gate2110(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2111(.a(s_223), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2112(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2113(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2114(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2647(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2648(.a(gate287inter0), .b(s_300), .O(gate287inter1));
  and2  gate2649(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2650(.a(s_300), .O(gate287inter3));
  inv1  gate2651(.a(s_301), .O(gate287inter4));
  nand2 gate2652(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2653(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2654(.a(G663), .O(gate287inter7));
  inv1  gate2655(.a(G815), .O(gate287inter8));
  nand2 gate2656(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2657(.a(s_301), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2658(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2659(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2660(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2143(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2144(.a(gate293inter0), .b(s_228), .O(gate293inter1));
  and2  gate2145(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2146(.a(s_228), .O(gate293inter3));
  inv1  gate2147(.a(s_229), .O(gate293inter4));
  nand2 gate2148(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2149(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2150(.a(G828), .O(gate293inter7));
  inv1  gate2151(.a(G829), .O(gate293inter8));
  nand2 gate2152(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2153(.a(s_229), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2154(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2155(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2156(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1261(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1262(.a(gate295inter0), .b(s_102), .O(gate295inter1));
  and2  gate1263(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1264(.a(s_102), .O(gate295inter3));
  inv1  gate1265(.a(s_103), .O(gate295inter4));
  nand2 gate1266(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1267(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1268(.a(G830), .O(gate295inter7));
  inv1  gate1269(.a(G831), .O(gate295inter8));
  nand2 gate1270(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1271(.a(s_103), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1272(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1273(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1274(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate2549(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2550(.a(gate296inter0), .b(s_286), .O(gate296inter1));
  and2  gate2551(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2552(.a(s_286), .O(gate296inter3));
  inv1  gate2553(.a(s_287), .O(gate296inter4));
  nand2 gate2554(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2555(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2556(.a(G826), .O(gate296inter7));
  inv1  gate2557(.a(G827), .O(gate296inter8));
  nand2 gate2558(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2559(.a(s_287), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2560(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2561(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2562(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2591(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2592(.a(gate388inter0), .b(s_292), .O(gate388inter1));
  and2  gate2593(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2594(.a(s_292), .O(gate388inter3));
  inv1  gate2595(.a(s_293), .O(gate388inter4));
  nand2 gate2596(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2597(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2598(.a(G2), .O(gate388inter7));
  inv1  gate2599(.a(G1039), .O(gate388inter8));
  nand2 gate2600(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2601(.a(s_293), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2602(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2603(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2604(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2241(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2242(.a(gate389inter0), .b(s_242), .O(gate389inter1));
  and2  gate2243(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2244(.a(s_242), .O(gate389inter3));
  inv1  gate2245(.a(s_243), .O(gate389inter4));
  nand2 gate2246(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2247(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2248(.a(G3), .O(gate389inter7));
  inv1  gate2249(.a(G1042), .O(gate389inter8));
  nand2 gate2250(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2251(.a(s_243), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2252(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2253(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2254(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1359(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1360(.a(gate390inter0), .b(s_116), .O(gate390inter1));
  and2  gate1361(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1362(.a(s_116), .O(gate390inter3));
  inv1  gate1363(.a(s_117), .O(gate390inter4));
  nand2 gate1364(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1365(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1366(.a(G4), .O(gate390inter7));
  inv1  gate1367(.a(G1045), .O(gate390inter8));
  nand2 gate1368(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1369(.a(s_117), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1370(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1371(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1372(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1051(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1052(.a(gate391inter0), .b(s_72), .O(gate391inter1));
  and2  gate1053(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1054(.a(s_72), .O(gate391inter3));
  inv1  gate1055(.a(s_73), .O(gate391inter4));
  nand2 gate1056(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1057(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1058(.a(G5), .O(gate391inter7));
  inv1  gate1059(.a(G1048), .O(gate391inter8));
  nand2 gate1060(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1061(.a(s_73), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1062(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1063(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1064(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate2157(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2158(.a(gate393inter0), .b(s_230), .O(gate393inter1));
  and2  gate2159(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2160(.a(s_230), .O(gate393inter3));
  inv1  gate2161(.a(s_231), .O(gate393inter4));
  nand2 gate2162(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2163(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2164(.a(G7), .O(gate393inter7));
  inv1  gate2165(.a(G1054), .O(gate393inter8));
  nand2 gate2166(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2167(.a(s_231), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2168(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2169(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2170(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1149(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1150(.a(gate394inter0), .b(s_86), .O(gate394inter1));
  and2  gate1151(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1152(.a(s_86), .O(gate394inter3));
  inv1  gate1153(.a(s_87), .O(gate394inter4));
  nand2 gate1154(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1155(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1156(.a(G8), .O(gate394inter7));
  inv1  gate1157(.a(G1057), .O(gate394inter8));
  nand2 gate1158(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1159(.a(s_87), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1160(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1161(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1162(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1891(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1892(.a(gate395inter0), .b(s_192), .O(gate395inter1));
  and2  gate1893(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1894(.a(s_192), .O(gate395inter3));
  inv1  gate1895(.a(s_193), .O(gate395inter4));
  nand2 gate1896(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1897(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1898(.a(G9), .O(gate395inter7));
  inv1  gate1899(.a(G1060), .O(gate395inter8));
  nand2 gate1900(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1901(.a(s_193), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1902(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1903(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1904(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2213(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2214(.a(gate396inter0), .b(s_238), .O(gate396inter1));
  and2  gate2215(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2216(.a(s_238), .O(gate396inter3));
  inv1  gate2217(.a(s_239), .O(gate396inter4));
  nand2 gate2218(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2219(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2220(.a(G10), .O(gate396inter7));
  inv1  gate2221(.a(G1063), .O(gate396inter8));
  nand2 gate2222(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2223(.a(s_239), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2224(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2225(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2226(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2689(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2690(.a(gate398inter0), .b(s_306), .O(gate398inter1));
  and2  gate2691(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2692(.a(s_306), .O(gate398inter3));
  inv1  gate2693(.a(s_307), .O(gate398inter4));
  nand2 gate2694(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2695(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2696(.a(G12), .O(gate398inter7));
  inv1  gate2697(.a(G1069), .O(gate398inter8));
  nand2 gate2698(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2699(.a(s_307), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2700(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2701(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2702(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1457(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1458(.a(gate399inter0), .b(s_130), .O(gate399inter1));
  and2  gate1459(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1460(.a(s_130), .O(gate399inter3));
  inv1  gate1461(.a(s_131), .O(gate399inter4));
  nand2 gate1462(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1463(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1464(.a(G13), .O(gate399inter7));
  inv1  gate1465(.a(G1072), .O(gate399inter8));
  nand2 gate1466(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1467(.a(s_131), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1468(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1469(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1470(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1331(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1332(.a(gate400inter0), .b(s_112), .O(gate400inter1));
  and2  gate1333(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1334(.a(s_112), .O(gate400inter3));
  inv1  gate1335(.a(s_113), .O(gate400inter4));
  nand2 gate1336(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1337(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1338(.a(G14), .O(gate400inter7));
  inv1  gate1339(.a(G1075), .O(gate400inter8));
  nand2 gate1340(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1341(.a(s_113), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1342(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1343(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1344(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1947(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1948(.a(gate406inter0), .b(s_200), .O(gate406inter1));
  and2  gate1949(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1950(.a(s_200), .O(gate406inter3));
  inv1  gate1951(.a(s_201), .O(gate406inter4));
  nand2 gate1952(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1953(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1954(.a(G20), .O(gate406inter7));
  inv1  gate1955(.a(G1093), .O(gate406inter8));
  nand2 gate1956(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1957(.a(s_201), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1958(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1959(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1960(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2535(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2536(.a(gate410inter0), .b(s_284), .O(gate410inter1));
  and2  gate2537(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2538(.a(s_284), .O(gate410inter3));
  inv1  gate2539(.a(s_285), .O(gate410inter4));
  nand2 gate2540(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2541(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2542(.a(G24), .O(gate410inter7));
  inv1  gate2543(.a(G1105), .O(gate410inter8));
  nand2 gate2544(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2545(.a(s_285), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2546(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2547(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2548(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate883(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate884(.a(gate412inter0), .b(s_48), .O(gate412inter1));
  and2  gate885(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate886(.a(s_48), .O(gate412inter3));
  inv1  gate887(.a(s_49), .O(gate412inter4));
  nand2 gate888(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate889(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate890(.a(G26), .O(gate412inter7));
  inv1  gate891(.a(G1111), .O(gate412inter8));
  nand2 gate892(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate893(.a(s_49), .b(gate412inter3), .O(gate412inter10));
  nor2  gate894(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate895(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate896(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate995(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate996(.a(gate414inter0), .b(s_64), .O(gate414inter1));
  and2  gate997(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate998(.a(s_64), .O(gate414inter3));
  inv1  gate999(.a(s_65), .O(gate414inter4));
  nand2 gate1000(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1001(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1002(.a(G28), .O(gate414inter7));
  inv1  gate1003(.a(G1117), .O(gate414inter8));
  nand2 gate1004(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1005(.a(s_65), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1006(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1007(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1008(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1023(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1024(.a(gate418inter0), .b(s_68), .O(gate418inter1));
  and2  gate1025(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1026(.a(s_68), .O(gate418inter3));
  inv1  gate1027(.a(s_69), .O(gate418inter4));
  nand2 gate1028(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1029(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1030(.a(G32), .O(gate418inter7));
  inv1  gate1031(.a(G1129), .O(gate418inter8));
  nand2 gate1032(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1033(.a(s_69), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1034(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1035(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1036(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2115(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2116(.a(gate419inter0), .b(s_224), .O(gate419inter1));
  and2  gate2117(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2118(.a(s_224), .O(gate419inter3));
  inv1  gate2119(.a(s_225), .O(gate419inter4));
  nand2 gate2120(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2121(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2122(.a(G1), .O(gate419inter7));
  inv1  gate2123(.a(G1132), .O(gate419inter8));
  nand2 gate2124(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2125(.a(s_225), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2126(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2127(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2128(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1037(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1038(.a(gate428inter0), .b(s_70), .O(gate428inter1));
  and2  gate1039(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1040(.a(s_70), .O(gate428inter3));
  inv1  gate1041(.a(s_71), .O(gate428inter4));
  nand2 gate1042(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1043(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1044(.a(G1048), .O(gate428inter7));
  inv1  gate1045(.a(G1144), .O(gate428inter8));
  nand2 gate1046(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1047(.a(s_71), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1048(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1049(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1050(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2311(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2312(.a(gate431inter0), .b(s_252), .O(gate431inter1));
  and2  gate2313(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2314(.a(s_252), .O(gate431inter3));
  inv1  gate2315(.a(s_253), .O(gate431inter4));
  nand2 gate2316(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2317(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2318(.a(G7), .O(gate431inter7));
  inv1  gate2319(.a(G1150), .O(gate431inter8));
  nand2 gate2320(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2321(.a(s_253), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2322(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2323(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2324(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1849(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1850(.a(gate432inter0), .b(s_186), .O(gate432inter1));
  and2  gate1851(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1852(.a(s_186), .O(gate432inter3));
  inv1  gate1853(.a(s_187), .O(gate432inter4));
  nand2 gate1854(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1855(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1856(.a(G1054), .O(gate432inter7));
  inv1  gate1857(.a(G1150), .O(gate432inter8));
  nand2 gate1858(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1859(.a(s_187), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1860(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1861(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1862(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2185(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2186(.a(gate433inter0), .b(s_234), .O(gate433inter1));
  and2  gate2187(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2188(.a(s_234), .O(gate433inter3));
  inv1  gate2189(.a(s_235), .O(gate433inter4));
  nand2 gate2190(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2191(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2192(.a(G8), .O(gate433inter7));
  inv1  gate2193(.a(G1153), .O(gate433inter8));
  nand2 gate2194(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2195(.a(s_235), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2196(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2197(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2198(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate2479(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2480(.a(gate434inter0), .b(s_276), .O(gate434inter1));
  and2  gate2481(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2482(.a(s_276), .O(gate434inter3));
  inv1  gate2483(.a(s_277), .O(gate434inter4));
  nand2 gate2484(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2485(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2486(.a(G1057), .O(gate434inter7));
  inv1  gate2487(.a(G1153), .O(gate434inter8));
  nand2 gate2488(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2489(.a(s_277), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2490(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2491(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2492(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1695(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1696(.a(gate436inter0), .b(s_164), .O(gate436inter1));
  and2  gate1697(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1698(.a(s_164), .O(gate436inter3));
  inv1  gate1699(.a(s_165), .O(gate436inter4));
  nand2 gate1700(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1701(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1702(.a(G1060), .O(gate436inter7));
  inv1  gate1703(.a(G1156), .O(gate436inter8));
  nand2 gate1704(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1705(.a(s_165), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1706(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1707(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1708(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2773(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2774(.a(gate442inter0), .b(s_318), .O(gate442inter1));
  and2  gate2775(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2776(.a(s_318), .O(gate442inter3));
  inv1  gate2777(.a(s_319), .O(gate442inter4));
  nand2 gate2778(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2779(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2780(.a(G1069), .O(gate442inter7));
  inv1  gate2781(.a(G1165), .O(gate442inter8));
  nand2 gate2782(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2783(.a(s_319), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2784(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2785(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2786(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1751(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1752(.a(gate443inter0), .b(s_172), .O(gate443inter1));
  and2  gate1753(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1754(.a(s_172), .O(gate443inter3));
  inv1  gate1755(.a(s_173), .O(gate443inter4));
  nand2 gate1756(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1757(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1758(.a(G13), .O(gate443inter7));
  inv1  gate1759(.a(G1168), .O(gate443inter8));
  nand2 gate1760(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1761(.a(s_173), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1762(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1763(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1764(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1219(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1220(.a(gate445inter0), .b(s_96), .O(gate445inter1));
  and2  gate1221(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1222(.a(s_96), .O(gate445inter3));
  inv1  gate1223(.a(s_97), .O(gate445inter4));
  nand2 gate1224(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1225(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1226(.a(G14), .O(gate445inter7));
  inv1  gate1227(.a(G1171), .O(gate445inter8));
  nand2 gate1228(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1229(.a(s_97), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1230(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1231(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1232(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1541(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1542(.a(gate447inter0), .b(s_142), .O(gate447inter1));
  and2  gate1543(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1544(.a(s_142), .O(gate447inter3));
  inv1  gate1545(.a(s_143), .O(gate447inter4));
  nand2 gate1546(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1547(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1548(.a(G15), .O(gate447inter7));
  inv1  gate1549(.a(G1174), .O(gate447inter8));
  nand2 gate1550(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1551(.a(s_143), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1552(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1553(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1554(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2521(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2522(.a(gate448inter0), .b(s_282), .O(gate448inter1));
  and2  gate2523(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2524(.a(s_282), .O(gate448inter3));
  inv1  gate2525(.a(s_283), .O(gate448inter4));
  nand2 gate2526(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2527(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2528(.a(G1078), .O(gate448inter7));
  inv1  gate2529(.a(G1174), .O(gate448inter8));
  nand2 gate2530(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2531(.a(s_283), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2532(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2533(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2534(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate603(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate604(.a(gate451inter0), .b(s_8), .O(gate451inter1));
  and2  gate605(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate606(.a(s_8), .O(gate451inter3));
  inv1  gate607(.a(s_9), .O(gate451inter4));
  nand2 gate608(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate609(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate610(.a(G17), .O(gate451inter7));
  inv1  gate611(.a(G1180), .O(gate451inter8));
  nand2 gate612(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate613(.a(s_9), .b(gate451inter3), .O(gate451inter10));
  nor2  gate614(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate615(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate616(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1177(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1178(.a(gate455inter0), .b(s_90), .O(gate455inter1));
  and2  gate1179(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1180(.a(s_90), .O(gate455inter3));
  inv1  gate1181(.a(s_91), .O(gate455inter4));
  nand2 gate1182(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1183(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1184(.a(G19), .O(gate455inter7));
  inv1  gate1185(.a(G1186), .O(gate455inter8));
  nand2 gate1186(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1187(.a(s_91), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1188(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1189(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1190(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1723(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1724(.a(gate457inter0), .b(s_168), .O(gate457inter1));
  and2  gate1725(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1726(.a(s_168), .O(gate457inter3));
  inv1  gate1727(.a(s_169), .O(gate457inter4));
  nand2 gate1728(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1729(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1730(.a(G20), .O(gate457inter7));
  inv1  gate1731(.a(G1189), .O(gate457inter8));
  nand2 gate1732(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1733(.a(s_169), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1734(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1735(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1736(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate701(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate702(.a(gate458inter0), .b(s_22), .O(gate458inter1));
  and2  gate703(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate704(.a(s_22), .O(gate458inter3));
  inv1  gate705(.a(s_23), .O(gate458inter4));
  nand2 gate706(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate707(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate708(.a(G1093), .O(gate458inter7));
  inv1  gate709(.a(G1189), .O(gate458inter8));
  nand2 gate710(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate711(.a(s_23), .b(gate458inter3), .O(gate458inter10));
  nor2  gate712(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate713(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate714(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1471(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1472(.a(gate463inter0), .b(s_132), .O(gate463inter1));
  and2  gate1473(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1474(.a(s_132), .O(gate463inter3));
  inv1  gate1475(.a(s_133), .O(gate463inter4));
  nand2 gate1476(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1477(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1478(.a(G23), .O(gate463inter7));
  inv1  gate1479(.a(G1198), .O(gate463inter8));
  nand2 gate1480(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1481(.a(s_133), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1482(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1483(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1484(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1625(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1626(.a(gate466inter0), .b(s_154), .O(gate466inter1));
  and2  gate1627(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1628(.a(s_154), .O(gate466inter3));
  inv1  gate1629(.a(s_155), .O(gate466inter4));
  nand2 gate1630(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1631(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1632(.a(G1105), .O(gate466inter7));
  inv1  gate1633(.a(G1201), .O(gate466inter8));
  nand2 gate1634(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1635(.a(s_155), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1636(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1637(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1638(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2577(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2578(.a(gate467inter0), .b(s_290), .O(gate467inter1));
  and2  gate2579(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2580(.a(s_290), .O(gate467inter3));
  inv1  gate2581(.a(s_291), .O(gate467inter4));
  nand2 gate2582(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2583(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2584(.a(G25), .O(gate467inter7));
  inv1  gate2585(.a(G1204), .O(gate467inter8));
  nand2 gate2586(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2587(.a(s_291), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2588(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2589(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2590(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate911(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate912(.a(gate470inter0), .b(s_52), .O(gate470inter1));
  and2  gate913(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate914(.a(s_52), .O(gate470inter3));
  inv1  gate915(.a(s_53), .O(gate470inter4));
  nand2 gate916(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate917(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate918(.a(G1111), .O(gate470inter7));
  inv1  gate919(.a(G1207), .O(gate470inter8));
  nand2 gate920(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate921(.a(s_53), .b(gate470inter3), .O(gate470inter10));
  nor2  gate922(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate923(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate924(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2395(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2396(.a(gate479inter0), .b(s_264), .O(gate479inter1));
  and2  gate2397(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2398(.a(s_264), .O(gate479inter3));
  inv1  gate2399(.a(s_265), .O(gate479inter4));
  nand2 gate2400(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2401(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2402(.a(G31), .O(gate479inter7));
  inv1  gate2403(.a(G1222), .O(gate479inter8));
  nand2 gate2404(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2405(.a(s_265), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2406(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2407(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2408(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate869(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate870(.a(gate482inter0), .b(s_46), .O(gate482inter1));
  and2  gate871(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate872(.a(s_46), .O(gate482inter3));
  inv1  gate873(.a(s_47), .O(gate482inter4));
  nand2 gate874(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate875(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate876(.a(G1129), .O(gate482inter7));
  inv1  gate877(.a(G1225), .O(gate482inter8));
  nand2 gate878(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate879(.a(s_47), .b(gate482inter3), .O(gate482inter10));
  nor2  gate880(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate881(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate882(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate659(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate660(.a(gate486inter0), .b(s_16), .O(gate486inter1));
  and2  gate661(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate662(.a(s_16), .O(gate486inter3));
  inv1  gate663(.a(s_17), .O(gate486inter4));
  nand2 gate664(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate665(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate666(.a(G1234), .O(gate486inter7));
  inv1  gate667(.a(G1235), .O(gate486inter8));
  nand2 gate668(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate669(.a(s_17), .b(gate486inter3), .O(gate486inter10));
  nor2  gate670(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate671(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate672(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1205(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1206(.a(gate489inter0), .b(s_94), .O(gate489inter1));
  and2  gate1207(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1208(.a(s_94), .O(gate489inter3));
  inv1  gate1209(.a(s_95), .O(gate489inter4));
  nand2 gate1210(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1211(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1212(.a(G1240), .O(gate489inter7));
  inv1  gate1213(.a(G1241), .O(gate489inter8));
  nand2 gate1214(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1215(.a(s_95), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1216(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1217(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1218(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate827(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate828(.a(gate491inter0), .b(s_40), .O(gate491inter1));
  and2  gate829(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate830(.a(s_40), .O(gate491inter3));
  inv1  gate831(.a(s_41), .O(gate491inter4));
  nand2 gate832(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate833(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate834(.a(G1244), .O(gate491inter7));
  inv1  gate835(.a(G1245), .O(gate491inter8));
  nand2 gate836(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate837(.a(s_41), .b(gate491inter3), .O(gate491inter10));
  nor2  gate838(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate839(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate840(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1835(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1836(.a(gate492inter0), .b(s_184), .O(gate492inter1));
  and2  gate1837(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1838(.a(s_184), .O(gate492inter3));
  inv1  gate1839(.a(s_185), .O(gate492inter4));
  nand2 gate1840(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1841(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1842(.a(G1246), .O(gate492inter7));
  inv1  gate1843(.a(G1247), .O(gate492inter8));
  nand2 gate1844(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1845(.a(s_185), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1846(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1847(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1848(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate2717(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2718(.a(gate495inter0), .b(s_310), .O(gate495inter1));
  and2  gate2719(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2720(.a(s_310), .O(gate495inter3));
  inv1  gate2721(.a(s_311), .O(gate495inter4));
  nand2 gate2722(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2723(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2724(.a(G1252), .O(gate495inter7));
  inv1  gate2725(.a(G1253), .O(gate495inter8));
  nand2 gate2726(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2727(.a(s_311), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2728(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2729(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2730(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate1905(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1906(.a(gate496inter0), .b(s_194), .O(gate496inter1));
  and2  gate1907(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1908(.a(s_194), .O(gate496inter3));
  inv1  gate1909(.a(s_195), .O(gate496inter4));
  nand2 gate1910(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1911(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1912(.a(G1254), .O(gate496inter7));
  inv1  gate1913(.a(G1255), .O(gate496inter8));
  nand2 gate1914(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1915(.a(s_195), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1916(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1917(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1918(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate2423(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2424(.a(gate497inter0), .b(s_268), .O(gate497inter1));
  and2  gate2425(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2426(.a(s_268), .O(gate497inter3));
  inv1  gate2427(.a(s_269), .O(gate497inter4));
  nand2 gate2428(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2429(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2430(.a(G1256), .O(gate497inter7));
  inv1  gate2431(.a(G1257), .O(gate497inter8));
  nand2 gate2432(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2433(.a(s_269), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2434(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2435(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2436(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1401(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1402(.a(gate498inter0), .b(s_122), .O(gate498inter1));
  and2  gate1403(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1404(.a(s_122), .O(gate498inter3));
  inv1  gate1405(.a(s_123), .O(gate498inter4));
  nand2 gate1406(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1407(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1408(.a(G1258), .O(gate498inter7));
  inv1  gate1409(.a(G1259), .O(gate498inter8));
  nand2 gate1410(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1411(.a(s_123), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1412(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1413(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1414(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2339(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2340(.a(gate500inter0), .b(s_256), .O(gate500inter1));
  and2  gate2341(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2342(.a(s_256), .O(gate500inter3));
  inv1  gate2343(.a(s_257), .O(gate500inter4));
  nand2 gate2344(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2345(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2346(.a(G1262), .O(gate500inter7));
  inv1  gate2347(.a(G1263), .O(gate500inter8));
  nand2 gate2348(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2349(.a(s_257), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2350(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2351(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2352(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1793(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1794(.a(gate503inter0), .b(s_178), .O(gate503inter1));
  and2  gate1795(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1796(.a(s_178), .O(gate503inter3));
  inv1  gate1797(.a(s_179), .O(gate503inter4));
  nand2 gate1798(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1799(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1800(.a(G1268), .O(gate503inter7));
  inv1  gate1801(.a(G1269), .O(gate503inter8));
  nand2 gate1802(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1803(.a(s_179), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1804(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1805(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1806(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2493(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2494(.a(gate508inter0), .b(s_278), .O(gate508inter1));
  and2  gate2495(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2496(.a(s_278), .O(gate508inter3));
  inv1  gate2497(.a(s_279), .O(gate508inter4));
  nand2 gate2498(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2499(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2500(.a(G1278), .O(gate508inter7));
  inv1  gate2501(.a(G1279), .O(gate508inter8));
  nand2 gate2502(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2503(.a(s_279), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2504(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2505(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2506(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1961(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1962(.a(gate509inter0), .b(s_202), .O(gate509inter1));
  and2  gate1963(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1964(.a(s_202), .O(gate509inter3));
  inv1  gate1965(.a(s_203), .O(gate509inter4));
  nand2 gate1966(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1967(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1968(.a(G1280), .O(gate509inter7));
  inv1  gate1969(.a(G1281), .O(gate509inter8));
  nand2 gate1970(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1971(.a(s_203), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1972(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1973(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1974(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate785(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate786(.a(gate510inter0), .b(s_34), .O(gate510inter1));
  and2  gate787(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate788(.a(s_34), .O(gate510inter3));
  inv1  gate789(.a(s_35), .O(gate510inter4));
  nand2 gate790(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate791(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate792(.a(G1282), .O(gate510inter7));
  inv1  gate793(.a(G1283), .O(gate510inter8));
  nand2 gate794(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate795(.a(s_35), .b(gate510inter3), .O(gate510inter10));
  nor2  gate796(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate797(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate798(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1499(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1500(.a(gate513inter0), .b(s_136), .O(gate513inter1));
  and2  gate1501(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1502(.a(s_136), .O(gate513inter3));
  inv1  gate1503(.a(s_137), .O(gate513inter4));
  nand2 gate1504(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1505(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1506(.a(G1288), .O(gate513inter7));
  inv1  gate1507(.a(G1289), .O(gate513inter8));
  nand2 gate1508(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1509(.a(s_137), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1510(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1511(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1512(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule