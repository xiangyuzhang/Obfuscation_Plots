module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate981(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate982(.a(gate13inter0), .b(s_62), .O(gate13inter1));
  and2  gate983(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate984(.a(s_62), .O(gate13inter3));
  inv1  gate985(.a(s_63), .O(gate13inter4));
  nand2 gate986(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate987(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate988(.a(G9), .O(gate13inter7));
  inv1  gate989(.a(G10), .O(gate13inter8));
  nand2 gate990(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate991(.a(s_63), .b(gate13inter3), .O(gate13inter10));
  nor2  gate992(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate993(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate994(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate603(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate604(.a(gate16inter0), .b(s_8), .O(gate16inter1));
  and2  gate605(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate606(.a(s_8), .O(gate16inter3));
  inv1  gate607(.a(s_9), .O(gate16inter4));
  nand2 gate608(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate609(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate610(.a(G15), .O(gate16inter7));
  inv1  gate611(.a(G16), .O(gate16inter8));
  nand2 gate612(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate613(.a(s_9), .b(gate16inter3), .O(gate16inter10));
  nor2  gate614(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate615(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate616(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate729(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate730(.a(gate29inter0), .b(s_26), .O(gate29inter1));
  and2  gate731(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate732(.a(s_26), .O(gate29inter3));
  inv1  gate733(.a(s_27), .O(gate29inter4));
  nand2 gate734(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate735(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate736(.a(G3), .O(gate29inter7));
  inv1  gate737(.a(G7), .O(gate29inter8));
  nand2 gate738(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate739(.a(s_27), .b(gate29inter3), .O(gate29inter10));
  nor2  gate740(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate741(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate742(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1051(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1052(.a(gate37inter0), .b(s_72), .O(gate37inter1));
  and2  gate1053(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1054(.a(s_72), .O(gate37inter3));
  inv1  gate1055(.a(s_73), .O(gate37inter4));
  nand2 gate1056(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1057(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1058(.a(G19), .O(gate37inter7));
  inv1  gate1059(.a(G23), .O(gate37inter8));
  nand2 gate1060(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1061(.a(s_73), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1062(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1063(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1064(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1107(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1108(.a(gate55inter0), .b(s_80), .O(gate55inter1));
  and2  gate1109(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1110(.a(s_80), .O(gate55inter3));
  inv1  gate1111(.a(s_81), .O(gate55inter4));
  nand2 gate1112(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1113(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1114(.a(G15), .O(gate55inter7));
  inv1  gate1115(.a(G287), .O(gate55inter8));
  nand2 gate1116(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1117(.a(s_81), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1118(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1119(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1120(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1023(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1024(.a(gate65inter0), .b(s_68), .O(gate65inter1));
  and2  gate1025(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1026(.a(s_68), .O(gate65inter3));
  inv1  gate1027(.a(s_69), .O(gate65inter4));
  nand2 gate1028(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1029(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1030(.a(G25), .O(gate65inter7));
  inv1  gate1031(.a(G302), .O(gate65inter8));
  nand2 gate1032(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1033(.a(s_69), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1034(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1035(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1036(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate771(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate772(.a(gate94inter0), .b(s_32), .O(gate94inter1));
  and2  gate773(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate774(.a(s_32), .O(gate94inter3));
  inv1  gate775(.a(s_33), .O(gate94inter4));
  nand2 gate776(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate777(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate778(.a(G22), .O(gate94inter7));
  inv1  gate779(.a(G344), .O(gate94inter8));
  nand2 gate780(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate781(.a(s_33), .b(gate94inter3), .O(gate94inter10));
  nor2  gate782(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate783(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate784(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate701(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate702(.a(gate109inter0), .b(s_22), .O(gate109inter1));
  and2  gate703(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate704(.a(s_22), .O(gate109inter3));
  inv1  gate705(.a(s_23), .O(gate109inter4));
  nand2 gate706(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate707(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate708(.a(G370), .O(gate109inter7));
  inv1  gate709(.a(G371), .O(gate109inter8));
  nand2 gate710(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate711(.a(s_23), .b(gate109inter3), .O(gate109inter10));
  nor2  gate712(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate713(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate714(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate617(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate618(.a(gate113inter0), .b(s_10), .O(gate113inter1));
  and2  gate619(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate620(.a(s_10), .O(gate113inter3));
  inv1  gate621(.a(s_11), .O(gate113inter4));
  nand2 gate622(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate623(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate624(.a(G378), .O(gate113inter7));
  inv1  gate625(.a(G379), .O(gate113inter8));
  nand2 gate626(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate627(.a(s_11), .b(gate113inter3), .O(gate113inter10));
  nor2  gate628(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate629(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate630(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1093(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1094(.a(gate120inter0), .b(s_78), .O(gate120inter1));
  and2  gate1095(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1096(.a(s_78), .O(gate120inter3));
  inv1  gate1097(.a(s_79), .O(gate120inter4));
  nand2 gate1098(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1099(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1100(.a(G392), .O(gate120inter7));
  inv1  gate1101(.a(G393), .O(gate120inter8));
  nand2 gate1102(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1103(.a(s_79), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1104(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1105(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1106(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate855(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate856(.a(gate122inter0), .b(s_44), .O(gate122inter1));
  and2  gate857(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate858(.a(s_44), .O(gate122inter3));
  inv1  gate859(.a(s_45), .O(gate122inter4));
  nand2 gate860(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate861(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate862(.a(G396), .O(gate122inter7));
  inv1  gate863(.a(G397), .O(gate122inter8));
  nand2 gate864(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate865(.a(s_45), .b(gate122inter3), .O(gate122inter10));
  nor2  gate866(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate867(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate868(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate911(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate912(.a(gate150inter0), .b(s_52), .O(gate150inter1));
  and2  gate913(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate914(.a(s_52), .O(gate150inter3));
  inv1  gate915(.a(s_53), .O(gate150inter4));
  nand2 gate916(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate917(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate918(.a(G504), .O(gate150inter7));
  inv1  gate919(.a(G507), .O(gate150inter8));
  nand2 gate920(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate921(.a(s_53), .b(gate150inter3), .O(gate150inter10));
  nor2  gate922(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate923(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate924(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate897(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate898(.a(gate154inter0), .b(s_50), .O(gate154inter1));
  and2  gate899(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate900(.a(s_50), .O(gate154inter3));
  inv1  gate901(.a(s_51), .O(gate154inter4));
  nand2 gate902(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate903(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate904(.a(G429), .O(gate154inter7));
  inv1  gate905(.a(G522), .O(gate154inter8));
  nand2 gate906(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate907(.a(s_51), .b(gate154inter3), .O(gate154inter10));
  nor2  gate908(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate909(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate910(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate673(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate674(.a(gate158inter0), .b(s_18), .O(gate158inter1));
  and2  gate675(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate676(.a(s_18), .O(gate158inter3));
  inv1  gate677(.a(s_19), .O(gate158inter4));
  nand2 gate678(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate679(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate680(.a(G441), .O(gate158inter7));
  inv1  gate681(.a(G528), .O(gate158inter8));
  nand2 gate682(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate683(.a(s_19), .b(gate158inter3), .O(gate158inter10));
  nor2  gate684(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate685(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate686(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate645(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate646(.a(gate166inter0), .b(s_14), .O(gate166inter1));
  and2  gate647(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate648(.a(s_14), .O(gate166inter3));
  inv1  gate649(.a(s_15), .O(gate166inter4));
  nand2 gate650(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate651(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate652(.a(G465), .O(gate166inter7));
  inv1  gate653(.a(G540), .O(gate166inter8));
  nand2 gate654(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate655(.a(s_15), .b(gate166inter3), .O(gate166inter10));
  nor2  gate656(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate657(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate658(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate575(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate576(.a(gate175inter0), .b(s_4), .O(gate175inter1));
  and2  gate577(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate578(.a(s_4), .O(gate175inter3));
  inv1  gate579(.a(s_5), .O(gate175inter4));
  nand2 gate580(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate581(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate582(.a(G492), .O(gate175inter7));
  inv1  gate583(.a(G555), .O(gate175inter8));
  nand2 gate584(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate585(.a(s_5), .b(gate175inter3), .O(gate175inter10));
  nor2  gate586(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate587(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate588(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1037(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1038(.a(gate196inter0), .b(s_70), .O(gate196inter1));
  and2  gate1039(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1040(.a(s_70), .O(gate196inter3));
  inv1  gate1041(.a(s_71), .O(gate196inter4));
  nand2 gate1042(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1043(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1044(.a(G592), .O(gate196inter7));
  inv1  gate1045(.a(G593), .O(gate196inter8));
  nand2 gate1046(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1047(.a(s_71), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1048(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1049(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1050(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate687(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate688(.a(gate202inter0), .b(s_20), .O(gate202inter1));
  and2  gate689(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate690(.a(s_20), .O(gate202inter3));
  inv1  gate691(.a(s_21), .O(gate202inter4));
  nand2 gate692(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate693(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate694(.a(G612), .O(gate202inter7));
  inv1  gate695(.a(G617), .O(gate202inter8));
  nand2 gate696(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate697(.a(s_21), .b(gate202inter3), .O(gate202inter10));
  nor2  gate698(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate699(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate700(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate869(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate870(.a(gate213inter0), .b(s_46), .O(gate213inter1));
  and2  gate871(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate872(.a(s_46), .O(gate213inter3));
  inv1  gate873(.a(s_47), .O(gate213inter4));
  nand2 gate874(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate875(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate876(.a(G602), .O(gate213inter7));
  inv1  gate877(.a(G672), .O(gate213inter8));
  nand2 gate878(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate879(.a(s_47), .b(gate213inter3), .O(gate213inter10));
  nor2  gate880(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate881(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate882(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate883(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate884(.a(gate220inter0), .b(s_48), .O(gate220inter1));
  and2  gate885(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate886(.a(s_48), .O(gate220inter3));
  inv1  gate887(.a(s_49), .O(gate220inter4));
  nand2 gate888(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate889(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate890(.a(G637), .O(gate220inter7));
  inv1  gate891(.a(G681), .O(gate220inter8));
  nand2 gate892(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate893(.a(s_49), .b(gate220inter3), .O(gate220inter10));
  nor2  gate894(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate895(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate896(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate841(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate842(.a(gate224inter0), .b(s_42), .O(gate224inter1));
  and2  gate843(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate844(.a(s_42), .O(gate224inter3));
  inv1  gate845(.a(s_43), .O(gate224inter4));
  nand2 gate846(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate847(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate848(.a(G637), .O(gate224inter7));
  inv1  gate849(.a(G687), .O(gate224inter8));
  nand2 gate850(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate851(.a(s_43), .b(gate224inter3), .O(gate224inter10));
  nor2  gate852(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate853(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate854(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate939(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate940(.a(gate232inter0), .b(s_56), .O(gate232inter1));
  and2  gate941(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate942(.a(s_56), .O(gate232inter3));
  inv1  gate943(.a(s_57), .O(gate232inter4));
  nand2 gate944(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate945(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate946(.a(G704), .O(gate232inter7));
  inv1  gate947(.a(G705), .O(gate232inter8));
  nand2 gate948(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate949(.a(s_57), .b(gate232inter3), .O(gate232inter10));
  nor2  gate950(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate951(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate952(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1065(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1066(.a(gate237inter0), .b(s_74), .O(gate237inter1));
  and2  gate1067(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1068(.a(s_74), .O(gate237inter3));
  inv1  gate1069(.a(s_75), .O(gate237inter4));
  nand2 gate1070(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1071(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1072(.a(G254), .O(gate237inter7));
  inv1  gate1073(.a(G706), .O(gate237inter8));
  nand2 gate1074(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1075(.a(s_75), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1076(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1077(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1078(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate757(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate758(.a(gate246inter0), .b(s_30), .O(gate246inter1));
  and2  gate759(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate760(.a(s_30), .O(gate246inter3));
  inv1  gate761(.a(s_31), .O(gate246inter4));
  nand2 gate762(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate763(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate764(.a(G724), .O(gate246inter7));
  inv1  gate765(.a(G736), .O(gate246inter8));
  nand2 gate766(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate767(.a(s_31), .b(gate246inter3), .O(gate246inter10));
  nor2  gate768(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate769(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate770(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate967(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate968(.a(gate250inter0), .b(s_60), .O(gate250inter1));
  and2  gate969(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate970(.a(s_60), .O(gate250inter3));
  inv1  gate971(.a(s_61), .O(gate250inter4));
  nand2 gate972(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate973(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate974(.a(G706), .O(gate250inter7));
  inv1  gate975(.a(G742), .O(gate250inter8));
  nand2 gate976(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate977(.a(s_61), .b(gate250inter3), .O(gate250inter10));
  nor2  gate978(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate979(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate980(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate953(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate954(.a(gate256inter0), .b(s_58), .O(gate256inter1));
  and2  gate955(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate956(.a(s_58), .O(gate256inter3));
  inv1  gate957(.a(s_59), .O(gate256inter4));
  nand2 gate958(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate959(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate960(.a(G715), .O(gate256inter7));
  inv1  gate961(.a(G751), .O(gate256inter8));
  nand2 gate962(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate963(.a(s_59), .b(gate256inter3), .O(gate256inter10));
  nor2  gate964(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate965(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate966(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate659(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate660(.a(gate287inter0), .b(s_16), .O(gate287inter1));
  and2  gate661(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate662(.a(s_16), .O(gate287inter3));
  inv1  gate663(.a(s_17), .O(gate287inter4));
  nand2 gate664(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate665(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate666(.a(G663), .O(gate287inter7));
  inv1  gate667(.a(G815), .O(gate287inter8));
  nand2 gate668(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate669(.a(s_17), .b(gate287inter3), .O(gate287inter10));
  nor2  gate670(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate671(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate672(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate631(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate632(.a(gate290inter0), .b(s_12), .O(gate290inter1));
  and2  gate633(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate634(.a(s_12), .O(gate290inter3));
  inv1  gate635(.a(s_13), .O(gate290inter4));
  nand2 gate636(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate637(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate638(.a(G820), .O(gate290inter7));
  inv1  gate639(.a(G821), .O(gate290inter8));
  nand2 gate640(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate641(.a(s_13), .b(gate290inter3), .O(gate290inter10));
  nor2  gate642(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate643(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate644(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate547(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate548(.a(gate291inter0), .b(s_0), .O(gate291inter1));
  and2  gate549(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate550(.a(s_0), .O(gate291inter3));
  inv1  gate551(.a(s_1), .O(gate291inter4));
  nand2 gate552(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate553(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate554(.a(G822), .O(gate291inter7));
  inv1  gate555(.a(G823), .O(gate291inter8));
  nand2 gate556(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate557(.a(s_1), .b(gate291inter3), .O(gate291inter10));
  nor2  gate558(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate559(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate560(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1079(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1080(.a(gate292inter0), .b(s_76), .O(gate292inter1));
  and2  gate1081(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1082(.a(s_76), .O(gate292inter3));
  inv1  gate1083(.a(s_77), .O(gate292inter4));
  nand2 gate1084(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1085(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1086(.a(G824), .O(gate292inter7));
  inv1  gate1087(.a(G825), .O(gate292inter8));
  nand2 gate1088(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1089(.a(s_77), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1090(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1091(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1092(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate995(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate996(.a(gate402inter0), .b(s_64), .O(gate402inter1));
  and2  gate997(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate998(.a(s_64), .O(gate402inter3));
  inv1  gate999(.a(s_65), .O(gate402inter4));
  nand2 gate1000(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1001(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1002(.a(G16), .O(gate402inter7));
  inv1  gate1003(.a(G1081), .O(gate402inter8));
  nand2 gate1004(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1005(.a(s_65), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1006(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1007(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1008(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate827(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate828(.a(gate417inter0), .b(s_40), .O(gate417inter1));
  and2  gate829(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate830(.a(s_40), .O(gate417inter3));
  inv1  gate831(.a(s_41), .O(gate417inter4));
  nand2 gate832(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate833(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate834(.a(G31), .O(gate417inter7));
  inv1  gate835(.a(G1126), .O(gate417inter8));
  nand2 gate836(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate837(.a(s_41), .b(gate417inter3), .O(gate417inter10));
  nor2  gate838(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate839(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate840(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1009(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1010(.a(gate419inter0), .b(s_66), .O(gate419inter1));
  and2  gate1011(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1012(.a(s_66), .O(gate419inter3));
  inv1  gate1013(.a(s_67), .O(gate419inter4));
  nand2 gate1014(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1015(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1016(.a(G1), .O(gate419inter7));
  inv1  gate1017(.a(G1132), .O(gate419inter8));
  nand2 gate1018(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1019(.a(s_67), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1020(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1021(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1022(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate785(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate786(.a(gate428inter0), .b(s_34), .O(gate428inter1));
  and2  gate787(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate788(.a(s_34), .O(gate428inter3));
  inv1  gate789(.a(s_35), .O(gate428inter4));
  nand2 gate790(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate791(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate792(.a(G1048), .O(gate428inter7));
  inv1  gate793(.a(G1144), .O(gate428inter8));
  nand2 gate794(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate795(.a(s_35), .b(gate428inter3), .O(gate428inter10));
  nor2  gate796(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate797(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate798(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate813(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate814(.a(gate434inter0), .b(s_38), .O(gate434inter1));
  and2  gate815(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate816(.a(s_38), .O(gate434inter3));
  inv1  gate817(.a(s_39), .O(gate434inter4));
  nand2 gate818(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate819(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate820(.a(G1057), .O(gate434inter7));
  inv1  gate821(.a(G1153), .O(gate434inter8));
  nand2 gate822(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate823(.a(s_39), .b(gate434inter3), .O(gate434inter10));
  nor2  gate824(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate825(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate826(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate561(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate562(.a(gate473inter0), .b(s_2), .O(gate473inter1));
  and2  gate563(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate564(.a(s_2), .O(gate473inter3));
  inv1  gate565(.a(s_3), .O(gate473inter4));
  nand2 gate566(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate567(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate568(.a(G28), .O(gate473inter7));
  inv1  gate569(.a(G1213), .O(gate473inter8));
  nand2 gate570(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate571(.a(s_3), .b(gate473inter3), .O(gate473inter10));
  nor2  gate572(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate573(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate574(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate715(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate716(.a(gate479inter0), .b(s_24), .O(gate479inter1));
  and2  gate717(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate718(.a(s_24), .O(gate479inter3));
  inv1  gate719(.a(s_25), .O(gate479inter4));
  nand2 gate720(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate721(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate722(.a(G31), .O(gate479inter7));
  inv1  gate723(.a(G1222), .O(gate479inter8));
  nand2 gate724(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate725(.a(s_25), .b(gate479inter3), .O(gate479inter10));
  nor2  gate726(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate727(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate728(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate589(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate590(.a(gate495inter0), .b(s_6), .O(gate495inter1));
  and2  gate591(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate592(.a(s_6), .O(gate495inter3));
  inv1  gate593(.a(s_7), .O(gate495inter4));
  nand2 gate594(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate595(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate596(.a(G1252), .O(gate495inter7));
  inv1  gate597(.a(G1253), .O(gate495inter8));
  nand2 gate598(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate599(.a(s_7), .b(gate495inter3), .O(gate495inter10));
  nor2  gate600(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate601(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate602(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate743(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate744(.a(gate499inter0), .b(s_28), .O(gate499inter1));
  and2  gate745(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate746(.a(s_28), .O(gate499inter3));
  inv1  gate747(.a(s_29), .O(gate499inter4));
  nand2 gate748(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate749(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate750(.a(G1260), .O(gate499inter7));
  inv1  gate751(.a(G1261), .O(gate499inter8));
  nand2 gate752(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate753(.a(s_29), .b(gate499inter3), .O(gate499inter10));
  nor2  gate754(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate755(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate756(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate925(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate926(.a(gate510inter0), .b(s_54), .O(gate510inter1));
  and2  gate927(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate928(.a(s_54), .O(gate510inter3));
  inv1  gate929(.a(s_55), .O(gate510inter4));
  nand2 gate930(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate931(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate932(.a(G1282), .O(gate510inter7));
  inv1  gate933(.a(G1283), .O(gate510inter8));
  nand2 gate934(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate935(.a(s_55), .b(gate510inter3), .O(gate510inter10));
  nor2  gate936(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate937(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate938(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate799(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate800(.a(gate512inter0), .b(s_36), .O(gate512inter1));
  and2  gate801(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate802(.a(s_36), .O(gate512inter3));
  inv1  gate803(.a(s_37), .O(gate512inter4));
  nand2 gate804(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate805(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate806(.a(G1286), .O(gate512inter7));
  inv1  gate807(.a(G1287), .O(gate512inter8));
  nand2 gate808(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate809(.a(s_37), .b(gate512inter3), .O(gate512inter10));
  nor2  gate810(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate811(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate812(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule