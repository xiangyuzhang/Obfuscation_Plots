module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1695(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1696(.a(gate9inter0), .b(s_164), .O(gate9inter1));
  and2  gate1697(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1698(.a(s_164), .O(gate9inter3));
  inv1  gate1699(.a(s_165), .O(gate9inter4));
  nand2 gate1700(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1701(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1702(.a(G1), .O(gate9inter7));
  inv1  gate1703(.a(G2), .O(gate9inter8));
  nand2 gate1704(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1705(.a(s_165), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1706(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1707(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1708(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1555(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1556(.a(gate13inter0), .b(s_144), .O(gate13inter1));
  and2  gate1557(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1558(.a(s_144), .O(gate13inter3));
  inv1  gate1559(.a(s_145), .O(gate13inter4));
  nand2 gate1560(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1561(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1562(.a(G9), .O(gate13inter7));
  inv1  gate1563(.a(G10), .O(gate13inter8));
  nand2 gate1564(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1565(.a(s_145), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1566(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1567(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1568(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate687(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate688(.a(gate16inter0), .b(s_20), .O(gate16inter1));
  and2  gate689(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate690(.a(s_20), .O(gate16inter3));
  inv1  gate691(.a(s_21), .O(gate16inter4));
  nand2 gate692(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate693(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate694(.a(G15), .O(gate16inter7));
  inv1  gate695(.a(G16), .O(gate16inter8));
  nand2 gate696(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate697(.a(s_21), .b(gate16inter3), .O(gate16inter10));
  nor2  gate698(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate699(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate700(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1807(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1808(.a(gate18inter0), .b(s_180), .O(gate18inter1));
  and2  gate1809(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1810(.a(s_180), .O(gate18inter3));
  inv1  gate1811(.a(s_181), .O(gate18inter4));
  nand2 gate1812(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1813(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1814(.a(G19), .O(gate18inter7));
  inv1  gate1815(.a(G20), .O(gate18inter8));
  nand2 gate1816(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1817(.a(s_181), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1818(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1819(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1820(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1709(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1710(.a(gate32inter0), .b(s_166), .O(gate32inter1));
  and2  gate1711(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1712(.a(s_166), .O(gate32inter3));
  inv1  gate1713(.a(s_167), .O(gate32inter4));
  nand2 gate1714(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1715(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1716(.a(G12), .O(gate32inter7));
  inv1  gate1717(.a(G16), .O(gate32inter8));
  nand2 gate1718(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1719(.a(s_167), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1720(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1721(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1722(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1667(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1668(.a(gate34inter0), .b(s_160), .O(gate34inter1));
  and2  gate1669(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1670(.a(s_160), .O(gate34inter3));
  inv1  gate1671(.a(s_161), .O(gate34inter4));
  nand2 gate1672(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1673(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1674(.a(G25), .O(gate34inter7));
  inv1  gate1675(.a(G29), .O(gate34inter8));
  nand2 gate1676(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1677(.a(s_161), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1678(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1679(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1680(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1751(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1752(.a(gate36inter0), .b(s_172), .O(gate36inter1));
  and2  gate1753(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1754(.a(s_172), .O(gate36inter3));
  inv1  gate1755(.a(s_173), .O(gate36inter4));
  nand2 gate1756(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1757(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1758(.a(G26), .O(gate36inter7));
  inv1  gate1759(.a(G30), .O(gate36inter8));
  nand2 gate1760(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1761(.a(s_173), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1762(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1763(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1764(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1275(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1276(.a(gate38inter0), .b(s_104), .O(gate38inter1));
  and2  gate1277(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1278(.a(s_104), .O(gate38inter3));
  inv1  gate1279(.a(s_105), .O(gate38inter4));
  nand2 gate1280(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1281(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1282(.a(G27), .O(gate38inter7));
  inv1  gate1283(.a(G31), .O(gate38inter8));
  nand2 gate1284(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1285(.a(s_105), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1286(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1287(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1288(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate799(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate800(.a(gate39inter0), .b(s_36), .O(gate39inter1));
  and2  gate801(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate802(.a(s_36), .O(gate39inter3));
  inv1  gate803(.a(s_37), .O(gate39inter4));
  nand2 gate804(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate805(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate806(.a(G20), .O(gate39inter7));
  inv1  gate807(.a(G24), .O(gate39inter8));
  nand2 gate808(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate809(.a(s_37), .b(gate39inter3), .O(gate39inter10));
  nor2  gate810(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate811(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate812(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1499(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1500(.a(gate45inter0), .b(s_136), .O(gate45inter1));
  and2  gate1501(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1502(.a(s_136), .O(gate45inter3));
  inv1  gate1503(.a(s_137), .O(gate45inter4));
  nand2 gate1504(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1505(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1506(.a(G5), .O(gate45inter7));
  inv1  gate1507(.a(G272), .O(gate45inter8));
  nand2 gate1508(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1509(.a(s_137), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1510(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1511(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1512(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate743(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate744(.a(gate46inter0), .b(s_28), .O(gate46inter1));
  and2  gate745(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate746(.a(s_28), .O(gate46inter3));
  inv1  gate747(.a(s_29), .O(gate46inter4));
  nand2 gate748(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate749(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate750(.a(G6), .O(gate46inter7));
  inv1  gate751(.a(G272), .O(gate46inter8));
  nand2 gate752(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate753(.a(s_29), .b(gate46inter3), .O(gate46inter10));
  nor2  gate754(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate755(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate756(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate855(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate856(.a(gate58inter0), .b(s_44), .O(gate58inter1));
  and2  gate857(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate858(.a(s_44), .O(gate58inter3));
  inv1  gate859(.a(s_45), .O(gate58inter4));
  nand2 gate860(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate861(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate862(.a(G18), .O(gate58inter7));
  inv1  gate863(.a(G290), .O(gate58inter8));
  nand2 gate864(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate865(.a(s_45), .b(gate58inter3), .O(gate58inter10));
  nor2  gate866(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate867(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate868(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1359(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1360(.a(gate62inter0), .b(s_116), .O(gate62inter1));
  and2  gate1361(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1362(.a(s_116), .O(gate62inter3));
  inv1  gate1363(.a(s_117), .O(gate62inter4));
  nand2 gate1364(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1365(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1366(.a(G22), .O(gate62inter7));
  inv1  gate1367(.a(G296), .O(gate62inter8));
  nand2 gate1368(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1369(.a(s_117), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1370(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1371(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1372(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1289(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1290(.a(gate65inter0), .b(s_106), .O(gate65inter1));
  and2  gate1291(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1292(.a(s_106), .O(gate65inter3));
  inv1  gate1293(.a(s_107), .O(gate65inter4));
  nand2 gate1294(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1295(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1296(.a(G25), .O(gate65inter7));
  inv1  gate1297(.a(G302), .O(gate65inter8));
  nand2 gate1298(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1299(.a(s_107), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1300(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1301(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1302(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1625(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1626(.a(gate66inter0), .b(s_154), .O(gate66inter1));
  and2  gate1627(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1628(.a(s_154), .O(gate66inter3));
  inv1  gate1629(.a(s_155), .O(gate66inter4));
  nand2 gate1630(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1631(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1632(.a(G26), .O(gate66inter7));
  inv1  gate1633(.a(G302), .O(gate66inter8));
  nand2 gate1634(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1635(.a(s_155), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1636(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1637(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1638(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1065(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1066(.a(gate67inter0), .b(s_74), .O(gate67inter1));
  and2  gate1067(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1068(.a(s_74), .O(gate67inter3));
  inv1  gate1069(.a(s_75), .O(gate67inter4));
  nand2 gate1070(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1071(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1072(.a(G27), .O(gate67inter7));
  inv1  gate1073(.a(G305), .O(gate67inter8));
  nand2 gate1074(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1075(.a(s_75), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1076(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1077(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1078(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1793(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1794(.a(gate68inter0), .b(s_178), .O(gate68inter1));
  and2  gate1795(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1796(.a(s_178), .O(gate68inter3));
  inv1  gate1797(.a(s_179), .O(gate68inter4));
  nand2 gate1798(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1799(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1800(.a(G28), .O(gate68inter7));
  inv1  gate1801(.a(G305), .O(gate68inter8));
  nand2 gate1802(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1803(.a(s_179), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1804(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1805(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1806(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1457(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1458(.a(gate91inter0), .b(s_130), .O(gate91inter1));
  and2  gate1459(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1460(.a(s_130), .O(gate91inter3));
  inv1  gate1461(.a(s_131), .O(gate91inter4));
  nand2 gate1462(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1463(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1464(.a(G25), .O(gate91inter7));
  inv1  gate1465(.a(G341), .O(gate91inter8));
  nand2 gate1466(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1467(.a(s_131), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1468(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1469(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1470(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate953(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate954(.a(gate96inter0), .b(s_58), .O(gate96inter1));
  and2  gate955(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate956(.a(s_58), .O(gate96inter3));
  inv1  gate957(.a(s_59), .O(gate96inter4));
  nand2 gate958(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate959(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate960(.a(G30), .O(gate96inter7));
  inv1  gate961(.a(G347), .O(gate96inter8));
  nand2 gate962(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate963(.a(s_59), .b(gate96inter3), .O(gate96inter10));
  nor2  gate964(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate965(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate966(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1401(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1402(.a(gate112inter0), .b(s_122), .O(gate112inter1));
  and2  gate1403(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1404(.a(s_122), .O(gate112inter3));
  inv1  gate1405(.a(s_123), .O(gate112inter4));
  nand2 gate1406(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1407(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1408(.a(G376), .O(gate112inter7));
  inv1  gate1409(.a(G377), .O(gate112inter8));
  nand2 gate1410(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1411(.a(s_123), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1412(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1413(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1414(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1527(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1528(.a(gate117inter0), .b(s_140), .O(gate117inter1));
  and2  gate1529(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1530(.a(s_140), .O(gate117inter3));
  inv1  gate1531(.a(s_141), .O(gate117inter4));
  nand2 gate1532(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1533(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1534(.a(G386), .O(gate117inter7));
  inv1  gate1535(.a(G387), .O(gate117inter8));
  nand2 gate1536(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1537(.a(s_141), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1538(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1539(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1540(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate813(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate814(.a(gate124inter0), .b(s_38), .O(gate124inter1));
  and2  gate815(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate816(.a(s_38), .O(gate124inter3));
  inv1  gate817(.a(s_39), .O(gate124inter4));
  nand2 gate818(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate819(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate820(.a(G400), .O(gate124inter7));
  inv1  gate821(.a(G401), .O(gate124inter8));
  nand2 gate822(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate823(.a(s_39), .b(gate124inter3), .O(gate124inter10));
  nor2  gate824(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate825(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate826(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1051(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1052(.a(gate127inter0), .b(s_72), .O(gate127inter1));
  and2  gate1053(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1054(.a(s_72), .O(gate127inter3));
  inv1  gate1055(.a(s_73), .O(gate127inter4));
  nand2 gate1056(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1057(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1058(.a(G406), .O(gate127inter7));
  inv1  gate1059(.a(G407), .O(gate127inter8));
  nand2 gate1060(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1061(.a(s_73), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1062(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1063(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1064(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1177(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1178(.a(gate130inter0), .b(s_90), .O(gate130inter1));
  and2  gate1179(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1180(.a(s_90), .O(gate130inter3));
  inv1  gate1181(.a(s_91), .O(gate130inter4));
  nand2 gate1182(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1183(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1184(.a(G412), .O(gate130inter7));
  inv1  gate1185(.a(G413), .O(gate130inter8));
  nand2 gate1186(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1187(.a(s_91), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1188(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1189(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1190(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate939(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate940(.a(gate133inter0), .b(s_56), .O(gate133inter1));
  and2  gate941(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate942(.a(s_56), .O(gate133inter3));
  inv1  gate943(.a(s_57), .O(gate133inter4));
  nand2 gate944(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate945(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate946(.a(G418), .O(gate133inter7));
  inv1  gate947(.a(G419), .O(gate133inter8));
  nand2 gate948(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate949(.a(s_57), .b(gate133inter3), .O(gate133inter10));
  nor2  gate950(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate951(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate952(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate575(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate576(.a(gate136inter0), .b(s_4), .O(gate136inter1));
  and2  gate577(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate578(.a(s_4), .O(gate136inter3));
  inv1  gate579(.a(s_5), .O(gate136inter4));
  nand2 gate580(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate581(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate582(.a(G424), .O(gate136inter7));
  inv1  gate583(.a(G425), .O(gate136inter8));
  nand2 gate584(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate585(.a(s_5), .b(gate136inter3), .O(gate136inter10));
  nor2  gate586(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate587(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate588(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate715(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate716(.a(gate137inter0), .b(s_24), .O(gate137inter1));
  and2  gate717(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate718(.a(s_24), .O(gate137inter3));
  inv1  gate719(.a(s_25), .O(gate137inter4));
  nand2 gate720(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate721(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate722(.a(G426), .O(gate137inter7));
  inv1  gate723(.a(G429), .O(gate137inter8));
  nand2 gate724(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate725(.a(s_25), .b(gate137inter3), .O(gate137inter10));
  nor2  gate726(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate727(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate728(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate869(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate870(.a(gate138inter0), .b(s_46), .O(gate138inter1));
  and2  gate871(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate872(.a(s_46), .O(gate138inter3));
  inv1  gate873(.a(s_47), .O(gate138inter4));
  nand2 gate874(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate875(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate876(.a(G432), .O(gate138inter7));
  inv1  gate877(.a(G435), .O(gate138inter8));
  nand2 gate878(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate879(.a(s_47), .b(gate138inter3), .O(gate138inter10));
  nor2  gate880(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate881(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate882(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate659(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate660(.a(gate139inter0), .b(s_16), .O(gate139inter1));
  and2  gate661(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate662(.a(s_16), .O(gate139inter3));
  inv1  gate663(.a(s_17), .O(gate139inter4));
  nand2 gate664(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate665(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate666(.a(G438), .O(gate139inter7));
  inv1  gate667(.a(G441), .O(gate139inter8));
  nand2 gate668(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate669(.a(s_17), .b(gate139inter3), .O(gate139inter10));
  nor2  gate670(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate671(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate672(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1485(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1486(.a(gate141inter0), .b(s_134), .O(gate141inter1));
  and2  gate1487(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1488(.a(s_134), .O(gate141inter3));
  inv1  gate1489(.a(s_135), .O(gate141inter4));
  nand2 gate1490(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1491(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1492(.a(G450), .O(gate141inter7));
  inv1  gate1493(.a(G453), .O(gate141inter8));
  nand2 gate1494(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1495(.a(s_135), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1496(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1497(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1498(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1443(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1444(.a(gate143inter0), .b(s_128), .O(gate143inter1));
  and2  gate1445(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1446(.a(s_128), .O(gate143inter3));
  inv1  gate1447(.a(s_129), .O(gate143inter4));
  nand2 gate1448(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1449(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1450(.a(G462), .O(gate143inter7));
  inv1  gate1451(.a(G465), .O(gate143inter8));
  nand2 gate1452(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1453(.a(s_129), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1454(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1455(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1456(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1653(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1654(.a(gate147inter0), .b(s_158), .O(gate147inter1));
  and2  gate1655(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1656(.a(s_158), .O(gate147inter3));
  inv1  gate1657(.a(s_159), .O(gate147inter4));
  nand2 gate1658(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1659(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1660(.a(G486), .O(gate147inter7));
  inv1  gate1661(.a(G489), .O(gate147inter8));
  nand2 gate1662(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1663(.a(s_159), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1664(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1665(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1666(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1037(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1038(.a(gate148inter0), .b(s_70), .O(gate148inter1));
  and2  gate1039(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1040(.a(s_70), .O(gate148inter3));
  inv1  gate1041(.a(s_71), .O(gate148inter4));
  nand2 gate1042(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1043(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1044(.a(G492), .O(gate148inter7));
  inv1  gate1045(.a(G495), .O(gate148inter8));
  nand2 gate1046(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1047(.a(s_71), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1048(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1049(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1050(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1737(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1738(.a(gate157inter0), .b(s_170), .O(gate157inter1));
  and2  gate1739(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1740(.a(s_170), .O(gate157inter3));
  inv1  gate1741(.a(s_171), .O(gate157inter4));
  nand2 gate1742(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1743(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1744(.a(G438), .O(gate157inter7));
  inv1  gate1745(.a(G528), .O(gate157inter8));
  nand2 gate1746(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1747(.a(s_171), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1748(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1749(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1750(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate995(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate996(.a(gate158inter0), .b(s_64), .O(gate158inter1));
  and2  gate997(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate998(.a(s_64), .O(gate158inter3));
  inv1  gate999(.a(s_65), .O(gate158inter4));
  nand2 gate1000(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1001(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1002(.a(G441), .O(gate158inter7));
  inv1  gate1003(.a(G528), .O(gate158inter8));
  nand2 gate1004(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1005(.a(s_65), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1006(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1007(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1008(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate701(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate702(.a(gate170inter0), .b(s_22), .O(gate170inter1));
  and2  gate703(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate704(.a(s_22), .O(gate170inter3));
  inv1  gate705(.a(s_23), .O(gate170inter4));
  nand2 gate706(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate707(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate708(.a(G477), .O(gate170inter7));
  inv1  gate709(.a(G546), .O(gate170inter8));
  nand2 gate710(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate711(.a(s_23), .b(gate170inter3), .O(gate170inter10));
  nor2  gate712(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate713(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate714(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1471(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1472(.a(gate174inter0), .b(s_132), .O(gate174inter1));
  and2  gate1473(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1474(.a(s_132), .O(gate174inter3));
  inv1  gate1475(.a(s_133), .O(gate174inter4));
  nand2 gate1476(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1477(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1478(.a(G489), .O(gate174inter7));
  inv1  gate1479(.a(G552), .O(gate174inter8));
  nand2 gate1480(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1481(.a(s_133), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1482(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1483(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1484(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1779(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1780(.a(gate183inter0), .b(s_176), .O(gate183inter1));
  and2  gate1781(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1782(.a(s_176), .O(gate183inter3));
  inv1  gate1783(.a(s_177), .O(gate183inter4));
  nand2 gate1784(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1785(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1786(.a(G516), .O(gate183inter7));
  inv1  gate1787(.a(G567), .O(gate183inter8));
  nand2 gate1788(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1789(.a(s_177), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1790(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1791(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1792(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1191(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1192(.a(gate188inter0), .b(s_92), .O(gate188inter1));
  and2  gate1193(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1194(.a(s_92), .O(gate188inter3));
  inv1  gate1195(.a(s_93), .O(gate188inter4));
  nand2 gate1196(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1197(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1198(.a(G576), .O(gate188inter7));
  inv1  gate1199(.a(G577), .O(gate188inter8));
  nand2 gate1200(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1201(.a(s_93), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1202(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1203(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1204(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1331(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1332(.a(gate191inter0), .b(s_112), .O(gate191inter1));
  and2  gate1333(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1334(.a(s_112), .O(gate191inter3));
  inv1  gate1335(.a(s_113), .O(gate191inter4));
  nand2 gate1336(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1337(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1338(.a(G582), .O(gate191inter7));
  inv1  gate1339(.a(G583), .O(gate191inter8));
  nand2 gate1340(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1341(.a(s_113), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1342(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1343(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1344(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1023(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1024(.a(gate192inter0), .b(s_68), .O(gate192inter1));
  and2  gate1025(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1026(.a(s_68), .O(gate192inter3));
  inv1  gate1027(.a(s_69), .O(gate192inter4));
  nand2 gate1028(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1029(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1030(.a(G584), .O(gate192inter7));
  inv1  gate1031(.a(G585), .O(gate192inter8));
  nand2 gate1032(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1033(.a(s_69), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1034(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1035(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1036(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1765(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1766(.a(gate198inter0), .b(s_174), .O(gate198inter1));
  and2  gate1767(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1768(.a(s_174), .O(gate198inter3));
  inv1  gate1769(.a(s_175), .O(gate198inter4));
  nand2 gate1770(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1771(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1772(.a(G596), .O(gate198inter7));
  inv1  gate1773(.a(G597), .O(gate198inter8));
  nand2 gate1774(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1775(.a(s_175), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1776(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1777(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1778(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate925(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate926(.a(gate203inter0), .b(s_54), .O(gate203inter1));
  and2  gate927(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate928(.a(s_54), .O(gate203inter3));
  inv1  gate929(.a(s_55), .O(gate203inter4));
  nand2 gate930(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate931(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate932(.a(G602), .O(gate203inter7));
  inv1  gate933(.a(G612), .O(gate203inter8));
  nand2 gate934(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate935(.a(s_55), .b(gate203inter3), .O(gate203inter10));
  nor2  gate936(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate937(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate938(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate883(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate884(.a(gate204inter0), .b(s_48), .O(gate204inter1));
  and2  gate885(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate886(.a(s_48), .O(gate204inter3));
  inv1  gate887(.a(s_49), .O(gate204inter4));
  nand2 gate888(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate889(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate890(.a(G607), .O(gate204inter7));
  inv1  gate891(.a(G617), .O(gate204inter8));
  nand2 gate892(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate893(.a(s_49), .b(gate204inter3), .O(gate204inter10));
  nor2  gate894(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate895(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate896(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1513(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1514(.a(gate205inter0), .b(s_138), .O(gate205inter1));
  and2  gate1515(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1516(.a(s_138), .O(gate205inter3));
  inv1  gate1517(.a(s_139), .O(gate205inter4));
  nand2 gate1518(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1519(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1520(.a(G622), .O(gate205inter7));
  inv1  gate1521(.a(G627), .O(gate205inter8));
  nand2 gate1522(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1523(.a(s_139), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1524(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1525(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1526(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate631(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate632(.a(gate219inter0), .b(s_12), .O(gate219inter1));
  and2  gate633(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate634(.a(s_12), .O(gate219inter3));
  inv1  gate635(.a(s_13), .O(gate219inter4));
  nand2 gate636(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate637(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate638(.a(G632), .O(gate219inter7));
  inv1  gate639(.a(G681), .O(gate219inter8));
  nand2 gate640(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate641(.a(s_13), .b(gate219inter3), .O(gate219inter10));
  nor2  gate642(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate643(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate644(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1597(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1598(.a(gate220inter0), .b(s_150), .O(gate220inter1));
  and2  gate1599(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1600(.a(s_150), .O(gate220inter3));
  inv1  gate1601(.a(s_151), .O(gate220inter4));
  nand2 gate1602(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1603(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1604(.a(G637), .O(gate220inter7));
  inv1  gate1605(.a(G681), .O(gate220inter8));
  nand2 gate1606(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1607(.a(s_151), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1608(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1609(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1610(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1639(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1640(.a(gate232inter0), .b(s_156), .O(gate232inter1));
  and2  gate1641(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1642(.a(s_156), .O(gate232inter3));
  inv1  gate1643(.a(s_157), .O(gate232inter4));
  nand2 gate1644(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1645(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1646(.a(G704), .O(gate232inter7));
  inv1  gate1647(.a(G705), .O(gate232inter8));
  nand2 gate1648(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1649(.a(s_157), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1650(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1651(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1652(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1723(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1724(.a(gate235inter0), .b(s_168), .O(gate235inter1));
  and2  gate1725(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1726(.a(s_168), .O(gate235inter3));
  inv1  gate1727(.a(s_169), .O(gate235inter4));
  nand2 gate1728(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1729(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1730(.a(G248), .O(gate235inter7));
  inv1  gate1731(.a(G724), .O(gate235inter8));
  nand2 gate1732(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1733(.a(s_169), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1734(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1735(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1736(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate729(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate730(.a(gate238inter0), .b(s_26), .O(gate238inter1));
  and2  gate731(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate732(.a(s_26), .O(gate238inter3));
  inv1  gate733(.a(s_27), .O(gate238inter4));
  nand2 gate734(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate735(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate736(.a(G257), .O(gate238inter7));
  inv1  gate737(.a(G709), .O(gate238inter8));
  nand2 gate738(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate739(.a(s_27), .b(gate238inter3), .O(gate238inter10));
  nor2  gate740(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate741(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate742(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1569(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1570(.a(gate239inter0), .b(s_146), .O(gate239inter1));
  and2  gate1571(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1572(.a(s_146), .O(gate239inter3));
  inv1  gate1573(.a(s_147), .O(gate239inter4));
  nand2 gate1574(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1575(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1576(.a(G260), .O(gate239inter7));
  inv1  gate1577(.a(G712), .O(gate239inter8));
  nand2 gate1578(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1579(.a(s_147), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1580(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1581(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1582(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1303(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1304(.a(gate243inter0), .b(s_108), .O(gate243inter1));
  and2  gate1305(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1306(.a(s_108), .O(gate243inter3));
  inv1  gate1307(.a(s_109), .O(gate243inter4));
  nand2 gate1308(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1309(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1310(.a(G245), .O(gate243inter7));
  inv1  gate1311(.a(G733), .O(gate243inter8));
  nand2 gate1312(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1313(.a(s_109), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1314(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1315(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1316(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate841(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate842(.a(gate244inter0), .b(s_42), .O(gate244inter1));
  and2  gate843(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate844(.a(s_42), .O(gate244inter3));
  inv1  gate845(.a(s_43), .O(gate244inter4));
  nand2 gate846(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate847(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate848(.a(G721), .O(gate244inter7));
  inv1  gate849(.a(G733), .O(gate244inter8));
  nand2 gate850(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate851(.a(s_43), .b(gate244inter3), .O(gate244inter10));
  nor2  gate852(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate853(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate854(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1317(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1318(.a(gate247inter0), .b(s_110), .O(gate247inter1));
  and2  gate1319(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1320(.a(s_110), .O(gate247inter3));
  inv1  gate1321(.a(s_111), .O(gate247inter4));
  nand2 gate1322(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1323(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1324(.a(G251), .O(gate247inter7));
  inv1  gate1325(.a(G739), .O(gate247inter8));
  nand2 gate1326(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1327(.a(s_111), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1328(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1329(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1330(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1611(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1612(.a(gate253inter0), .b(s_152), .O(gate253inter1));
  and2  gate1613(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1614(.a(s_152), .O(gate253inter3));
  inv1  gate1615(.a(s_153), .O(gate253inter4));
  nand2 gate1616(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1617(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1618(.a(G260), .O(gate253inter7));
  inv1  gate1619(.a(G748), .O(gate253inter8));
  nand2 gate1620(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1621(.a(s_153), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1622(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1623(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1624(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate771(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate772(.a(gate256inter0), .b(s_32), .O(gate256inter1));
  and2  gate773(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate774(.a(s_32), .O(gate256inter3));
  inv1  gate775(.a(s_33), .O(gate256inter4));
  nand2 gate776(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate777(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate778(.a(G715), .O(gate256inter7));
  inv1  gate779(.a(G751), .O(gate256inter8));
  nand2 gate780(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate781(.a(s_33), .b(gate256inter3), .O(gate256inter10));
  nor2  gate782(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate783(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate784(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate785(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate786(.a(gate261inter0), .b(s_34), .O(gate261inter1));
  and2  gate787(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate788(.a(s_34), .O(gate261inter3));
  inv1  gate789(.a(s_35), .O(gate261inter4));
  nand2 gate790(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate791(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate792(.a(G762), .O(gate261inter7));
  inv1  gate793(.a(G763), .O(gate261inter8));
  nand2 gate794(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate795(.a(s_35), .b(gate261inter3), .O(gate261inter10));
  nor2  gate796(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate797(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate798(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate561(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate562(.a(gate265inter0), .b(s_2), .O(gate265inter1));
  and2  gate563(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate564(.a(s_2), .O(gate265inter3));
  inv1  gate565(.a(s_3), .O(gate265inter4));
  nand2 gate566(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate567(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate568(.a(G642), .O(gate265inter7));
  inv1  gate569(.a(G770), .O(gate265inter8));
  nand2 gate570(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate571(.a(s_3), .b(gate265inter3), .O(gate265inter10));
  nor2  gate572(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate573(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate574(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1429(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1430(.a(gate267inter0), .b(s_126), .O(gate267inter1));
  and2  gate1431(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1432(.a(s_126), .O(gate267inter3));
  inv1  gate1433(.a(s_127), .O(gate267inter4));
  nand2 gate1434(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1435(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1436(.a(G648), .O(gate267inter7));
  inv1  gate1437(.a(G776), .O(gate267inter8));
  nand2 gate1438(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1439(.a(s_127), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1440(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1441(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1442(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1373(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1374(.a(gate269inter0), .b(s_118), .O(gate269inter1));
  and2  gate1375(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1376(.a(s_118), .O(gate269inter3));
  inv1  gate1377(.a(s_119), .O(gate269inter4));
  nand2 gate1378(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1379(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1380(.a(G654), .O(gate269inter7));
  inv1  gate1381(.a(G782), .O(gate269inter8));
  nand2 gate1382(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1383(.a(s_119), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1384(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1385(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1386(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate981(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate982(.a(gate271inter0), .b(s_62), .O(gate271inter1));
  and2  gate983(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate984(.a(s_62), .O(gate271inter3));
  inv1  gate985(.a(s_63), .O(gate271inter4));
  nand2 gate986(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate987(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate988(.a(G660), .O(gate271inter7));
  inv1  gate989(.a(G788), .O(gate271inter8));
  nand2 gate990(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate991(.a(s_63), .b(gate271inter3), .O(gate271inter10));
  nor2  gate992(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate993(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate994(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate617(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate618(.a(gate272inter0), .b(s_10), .O(gate272inter1));
  and2  gate619(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate620(.a(s_10), .O(gate272inter3));
  inv1  gate621(.a(s_11), .O(gate272inter4));
  nand2 gate622(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate623(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate624(.a(G663), .O(gate272inter7));
  inv1  gate625(.a(G791), .O(gate272inter8));
  nand2 gate626(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate627(.a(s_11), .b(gate272inter3), .O(gate272inter10));
  nor2  gate628(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate629(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate630(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1681(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1682(.a(gate277inter0), .b(s_162), .O(gate277inter1));
  and2  gate1683(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1684(.a(s_162), .O(gate277inter3));
  inv1  gate1685(.a(s_163), .O(gate277inter4));
  nand2 gate1686(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1687(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1688(.a(G648), .O(gate277inter7));
  inv1  gate1689(.a(G800), .O(gate277inter8));
  nand2 gate1690(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1691(.a(s_163), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1692(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1693(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1694(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1219(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1220(.a(gate278inter0), .b(s_96), .O(gate278inter1));
  and2  gate1221(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1222(.a(s_96), .O(gate278inter3));
  inv1  gate1223(.a(s_97), .O(gate278inter4));
  nand2 gate1224(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1225(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1226(.a(G776), .O(gate278inter7));
  inv1  gate1227(.a(G800), .O(gate278inter8));
  nand2 gate1228(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1229(.a(s_97), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1230(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1231(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1232(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1247(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1248(.a(gate284inter0), .b(s_100), .O(gate284inter1));
  and2  gate1249(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1250(.a(s_100), .O(gate284inter3));
  inv1  gate1251(.a(s_101), .O(gate284inter4));
  nand2 gate1252(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1253(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1254(.a(G785), .O(gate284inter7));
  inv1  gate1255(.a(G809), .O(gate284inter8));
  nand2 gate1256(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1257(.a(s_101), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1258(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1259(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1260(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1583(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1584(.a(gate287inter0), .b(s_148), .O(gate287inter1));
  and2  gate1585(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1586(.a(s_148), .O(gate287inter3));
  inv1  gate1587(.a(s_149), .O(gate287inter4));
  nand2 gate1588(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1589(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1590(.a(G663), .O(gate287inter7));
  inv1  gate1591(.a(G815), .O(gate287inter8));
  nand2 gate1592(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1593(.a(s_149), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1594(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1595(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1596(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1107(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1108(.a(gate291inter0), .b(s_80), .O(gate291inter1));
  and2  gate1109(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1110(.a(s_80), .O(gate291inter3));
  inv1  gate1111(.a(s_81), .O(gate291inter4));
  nand2 gate1112(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1113(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1114(.a(G822), .O(gate291inter7));
  inv1  gate1115(.a(G823), .O(gate291inter8));
  nand2 gate1116(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1117(.a(s_81), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1118(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1119(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1120(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate589(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate590(.a(gate388inter0), .b(s_6), .O(gate388inter1));
  and2  gate591(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate592(.a(s_6), .O(gate388inter3));
  inv1  gate593(.a(s_7), .O(gate388inter4));
  nand2 gate594(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate595(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate596(.a(G2), .O(gate388inter7));
  inv1  gate597(.a(G1039), .O(gate388inter8));
  nand2 gate598(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate599(.a(s_7), .b(gate388inter3), .O(gate388inter10));
  nor2  gate600(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate601(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate602(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1345(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1346(.a(gate389inter0), .b(s_114), .O(gate389inter1));
  and2  gate1347(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1348(.a(s_114), .O(gate389inter3));
  inv1  gate1349(.a(s_115), .O(gate389inter4));
  nand2 gate1350(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1351(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1352(.a(G3), .O(gate389inter7));
  inv1  gate1353(.a(G1042), .O(gate389inter8));
  nand2 gate1354(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1355(.a(s_115), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1356(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1357(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1358(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1093(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1094(.a(gate391inter0), .b(s_78), .O(gate391inter1));
  and2  gate1095(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1096(.a(s_78), .O(gate391inter3));
  inv1  gate1097(.a(s_79), .O(gate391inter4));
  nand2 gate1098(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1099(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1100(.a(G5), .O(gate391inter7));
  inv1  gate1101(.a(G1048), .O(gate391inter8));
  nand2 gate1102(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1103(.a(s_79), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1104(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1105(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1106(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1387(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1388(.a(gate393inter0), .b(s_120), .O(gate393inter1));
  and2  gate1389(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1390(.a(s_120), .O(gate393inter3));
  inv1  gate1391(.a(s_121), .O(gate393inter4));
  nand2 gate1392(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1393(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1394(.a(G7), .O(gate393inter7));
  inv1  gate1395(.a(G1054), .O(gate393inter8));
  nand2 gate1396(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1397(.a(s_121), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1398(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1399(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1400(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1149(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1150(.a(gate402inter0), .b(s_86), .O(gate402inter1));
  and2  gate1151(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1152(.a(s_86), .O(gate402inter3));
  inv1  gate1153(.a(s_87), .O(gate402inter4));
  nand2 gate1154(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1155(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1156(.a(G16), .O(gate402inter7));
  inv1  gate1157(.a(G1081), .O(gate402inter8));
  nand2 gate1158(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1159(.a(s_87), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1160(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1161(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1162(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate911(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate912(.a(gate411inter0), .b(s_52), .O(gate411inter1));
  and2  gate913(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate914(.a(s_52), .O(gate411inter3));
  inv1  gate915(.a(s_53), .O(gate411inter4));
  nand2 gate916(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate917(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate918(.a(G25), .O(gate411inter7));
  inv1  gate919(.a(G1108), .O(gate411inter8));
  nand2 gate920(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate921(.a(s_53), .b(gate411inter3), .O(gate411inter10));
  nor2  gate922(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate923(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate924(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate967(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate968(.a(gate420inter0), .b(s_60), .O(gate420inter1));
  and2  gate969(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate970(.a(s_60), .O(gate420inter3));
  inv1  gate971(.a(s_61), .O(gate420inter4));
  nand2 gate972(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate973(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate974(.a(G1036), .O(gate420inter7));
  inv1  gate975(.a(G1132), .O(gate420inter8));
  nand2 gate976(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate977(.a(s_61), .b(gate420inter3), .O(gate420inter10));
  nor2  gate978(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate979(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate980(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1541(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1542(.a(gate422inter0), .b(s_142), .O(gate422inter1));
  and2  gate1543(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1544(.a(s_142), .O(gate422inter3));
  inv1  gate1545(.a(s_143), .O(gate422inter4));
  nand2 gate1546(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1547(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1548(.a(G1039), .O(gate422inter7));
  inv1  gate1549(.a(G1135), .O(gate422inter8));
  nand2 gate1550(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1551(.a(s_143), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1552(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1553(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1554(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate603(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate604(.a(gate423inter0), .b(s_8), .O(gate423inter1));
  and2  gate605(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate606(.a(s_8), .O(gate423inter3));
  inv1  gate607(.a(s_9), .O(gate423inter4));
  nand2 gate608(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate609(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate610(.a(G3), .O(gate423inter7));
  inv1  gate611(.a(G1138), .O(gate423inter8));
  nand2 gate612(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate613(.a(s_9), .b(gate423inter3), .O(gate423inter10));
  nor2  gate614(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate615(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate616(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1205(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1206(.a(gate428inter0), .b(s_94), .O(gate428inter1));
  and2  gate1207(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1208(.a(s_94), .O(gate428inter3));
  inv1  gate1209(.a(s_95), .O(gate428inter4));
  nand2 gate1210(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1211(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1212(.a(G1048), .O(gate428inter7));
  inv1  gate1213(.a(G1144), .O(gate428inter8));
  nand2 gate1214(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1215(.a(s_95), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1216(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1217(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1218(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1415(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1416(.a(gate429inter0), .b(s_124), .O(gate429inter1));
  and2  gate1417(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1418(.a(s_124), .O(gate429inter3));
  inv1  gate1419(.a(s_125), .O(gate429inter4));
  nand2 gate1420(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1421(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1422(.a(G6), .O(gate429inter7));
  inv1  gate1423(.a(G1147), .O(gate429inter8));
  nand2 gate1424(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1425(.a(s_125), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1426(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1427(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1428(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate645(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate646(.a(gate432inter0), .b(s_14), .O(gate432inter1));
  and2  gate647(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate648(.a(s_14), .O(gate432inter3));
  inv1  gate649(.a(s_15), .O(gate432inter4));
  nand2 gate650(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate651(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate652(.a(G1054), .O(gate432inter7));
  inv1  gate653(.a(G1150), .O(gate432inter8));
  nand2 gate654(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate655(.a(s_15), .b(gate432inter3), .O(gate432inter10));
  nor2  gate656(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate657(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate658(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1121(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1122(.a(gate447inter0), .b(s_82), .O(gate447inter1));
  and2  gate1123(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1124(.a(s_82), .O(gate447inter3));
  inv1  gate1125(.a(s_83), .O(gate447inter4));
  nand2 gate1126(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1127(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1128(.a(G15), .O(gate447inter7));
  inv1  gate1129(.a(G1174), .O(gate447inter8));
  nand2 gate1130(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1131(.a(s_83), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1132(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1133(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1134(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1135(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1136(.a(gate451inter0), .b(s_84), .O(gate451inter1));
  and2  gate1137(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1138(.a(s_84), .O(gate451inter3));
  inv1  gate1139(.a(s_85), .O(gate451inter4));
  nand2 gate1140(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1141(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1142(.a(G17), .O(gate451inter7));
  inv1  gate1143(.a(G1180), .O(gate451inter8));
  nand2 gate1144(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1145(.a(s_85), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1146(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1147(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1148(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate897(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate898(.a(gate452inter0), .b(s_50), .O(gate452inter1));
  and2  gate899(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate900(.a(s_50), .O(gate452inter3));
  inv1  gate901(.a(s_51), .O(gate452inter4));
  nand2 gate902(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate903(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate904(.a(G1084), .O(gate452inter7));
  inv1  gate905(.a(G1180), .O(gate452inter8));
  nand2 gate906(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate907(.a(s_51), .b(gate452inter3), .O(gate452inter10));
  nor2  gate908(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate909(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate910(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate827(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate828(.a(gate470inter0), .b(s_40), .O(gate470inter1));
  and2  gate829(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate830(.a(s_40), .O(gate470inter3));
  inv1  gate831(.a(s_41), .O(gate470inter4));
  nand2 gate832(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate833(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate834(.a(G1111), .O(gate470inter7));
  inv1  gate835(.a(G1207), .O(gate470inter8));
  nand2 gate836(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate837(.a(s_41), .b(gate470inter3), .O(gate470inter10));
  nor2  gate838(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate839(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate840(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate547(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate548(.a(gate477inter0), .b(s_0), .O(gate477inter1));
  and2  gate549(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate550(.a(s_0), .O(gate477inter3));
  inv1  gate551(.a(s_1), .O(gate477inter4));
  nand2 gate552(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate553(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate554(.a(G30), .O(gate477inter7));
  inv1  gate555(.a(G1219), .O(gate477inter8));
  nand2 gate556(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate557(.a(s_1), .b(gate477inter3), .O(gate477inter10));
  nor2  gate558(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate559(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate560(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1009(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1010(.a(gate485inter0), .b(s_66), .O(gate485inter1));
  and2  gate1011(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1012(.a(s_66), .O(gate485inter3));
  inv1  gate1013(.a(s_67), .O(gate485inter4));
  nand2 gate1014(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1015(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1016(.a(G1232), .O(gate485inter7));
  inv1  gate1017(.a(G1233), .O(gate485inter8));
  nand2 gate1018(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1019(.a(s_67), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1020(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1021(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1022(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1233(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1234(.a(gate493inter0), .b(s_98), .O(gate493inter1));
  and2  gate1235(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1236(.a(s_98), .O(gate493inter3));
  inv1  gate1237(.a(s_99), .O(gate493inter4));
  nand2 gate1238(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1239(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1240(.a(G1248), .O(gate493inter7));
  inv1  gate1241(.a(G1249), .O(gate493inter8));
  nand2 gate1242(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1243(.a(s_99), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1244(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1245(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1246(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1261(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1262(.a(gate496inter0), .b(s_102), .O(gate496inter1));
  and2  gate1263(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1264(.a(s_102), .O(gate496inter3));
  inv1  gate1265(.a(s_103), .O(gate496inter4));
  nand2 gate1266(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1267(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1268(.a(G1254), .O(gate496inter7));
  inv1  gate1269(.a(G1255), .O(gate496inter8));
  nand2 gate1270(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1271(.a(s_103), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1272(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1273(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1274(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate673(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate674(.a(gate499inter0), .b(s_18), .O(gate499inter1));
  and2  gate675(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate676(.a(s_18), .O(gate499inter3));
  inv1  gate677(.a(s_19), .O(gate499inter4));
  nand2 gate678(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate679(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate680(.a(G1260), .O(gate499inter7));
  inv1  gate681(.a(G1261), .O(gate499inter8));
  nand2 gate682(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate683(.a(s_19), .b(gate499inter3), .O(gate499inter10));
  nor2  gate684(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate685(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate686(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1163(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1164(.a(gate502inter0), .b(s_88), .O(gate502inter1));
  and2  gate1165(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1166(.a(s_88), .O(gate502inter3));
  inv1  gate1167(.a(s_89), .O(gate502inter4));
  nand2 gate1168(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1169(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1170(.a(G1266), .O(gate502inter7));
  inv1  gate1171(.a(G1267), .O(gate502inter8));
  nand2 gate1172(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1173(.a(s_89), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1174(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1175(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1176(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate757(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate758(.a(gate508inter0), .b(s_30), .O(gate508inter1));
  and2  gate759(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate760(.a(s_30), .O(gate508inter3));
  inv1  gate761(.a(s_31), .O(gate508inter4));
  nand2 gate762(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate763(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate764(.a(G1278), .O(gate508inter7));
  inv1  gate765(.a(G1279), .O(gate508inter8));
  nand2 gate766(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate767(.a(s_31), .b(gate508inter3), .O(gate508inter10));
  nor2  gate768(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate769(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate770(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1079(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1080(.a(gate510inter0), .b(s_76), .O(gate510inter1));
  and2  gate1081(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1082(.a(s_76), .O(gate510inter3));
  inv1  gate1083(.a(s_77), .O(gate510inter4));
  nand2 gate1084(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1085(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1086(.a(G1282), .O(gate510inter7));
  inv1  gate1087(.a(G1283), .O(gate510inter8));
  nand2 gate1088(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1089(.a(s_77), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1090(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1091(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1092(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule