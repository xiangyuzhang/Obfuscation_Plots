module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate855(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate856(.a(gate13inter0), .b(s_44), .O(gate13inter1));
  and2  gate857(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate858(.a(s_44), .O(gate13inter3));
  inv1  gate859(.a(s_45), .O(gate13inter4));
  nand2 gate860(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate861(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate862(.a(G9), .O(gate13inter7));
  inv1  gate863(.a(G10), .O(gate13inter8));
  nand2 gate864(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate865(.a(s_45), .b(gate13inter3), .O(gate13inter10));
  nor2  gate866(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate867(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate868(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate547(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate548(.a(gate17inter0), .b(s_0), .O(gate17inter1));
  and2  gate549(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate550(.a(s_0), .O(gate17inter3));
  inv1  gate551(.a(s_1), .O(gate17inter4));
  nand2 gate552(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate553(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate554(.a(G17), .O(gate17inter7));
  inv1  gate555(.a(G18), .O(gate17inter8));
  nand2 gate556(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate557(.a(s_1), .b(gate17inter3), .O(gate17inter10));
  nor2  gate558(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate559(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate560(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1709(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1710(.a(gate19inter0), .b(s_166), .O(gate19inter1));
  and2  gate1711(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1712(.a(s_166), .O(gate19inter3));
  inv1  gate1713(.a(s_167), .O(gate19inter4));
  nand2 gate1714(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1715(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1716(.a(G21), .O(gate19inter7));
  inv1  gate1717(.a(G22), .O(gate19inter8));
  nand2 gate1718(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1719(.a(s_167), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1720(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1721(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1722(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2003(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2004(.a(gate22inter0), .b(s_208), .O(gate22inter1));
  and2  gate2005(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2006(.a(s_208), .O(gate22inter3));
  inv1  gate2007(.a(s_209), .O(gate22inter4));
  nand2 gate2008(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2009(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2010(.a(G27), .O(gate22inter7));
  inv1  gate2011(.a(G28), .O(gate22inter8));
  nand2 gate2012(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2013(.a(s_209), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2014(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2015(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2016(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate939(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate940(.a(gate29inter0), .b(s_56), .O(gate29inter1));
  and2  gate941(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate942(.a(s_56), .O(gate29inter3));
  inv1  gate943(.a(s_57), .O(gate29inter4));
  nand2 gate944(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate945(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate946(.a(G3), .O(gate29inter7));
  inv1  gate947(.a(G7), .O(gate29inter8));
  nand2 gate948(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate949(.a(s_57), .b(gate29inter3), .O(gate29inter10));
  nor2  gate950(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate951(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate952(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1989(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1990(.a(gate38inter0), .b(s_206), .O(gate38inter1));
  and2  gate1991(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1992(.a(s_206), .O(gate38inter3));
  inv1  gate1993(.a(s_207), .O(gate38inter4));
  nand2 gate1994(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1995(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1996(.a(G27), .O(gate38inter7));
  inv1  gate1997(.a(G31), .O(gate38inter8));
  nand2 gate1998(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1999(.a(s_207), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2000(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2001(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2002(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1275(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1276(.a(gate42inter0), .b(s_104), .O(gate42inter1));
  and2  gate1277(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1278(.a(s_104), .O(gate42inter3));
  inv1  gate1279(.a(s_105), .O(gate42inter4));
  nand2 gate1280(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1281(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1282(.a(G2), .O(gate42inter7));
  inv1  gate1283(.a(G266), .O(gate42inter8));
  nand2 gate1284(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1285(.a(s_105), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1286(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1287(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1288(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate589(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate590(.a(gate45inter0), .b(s_6), .O(gate45inter1));
  and2  gate591(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate592(.a(s_6), .O(gate45inter3));
  inv1  gate593(.a(s_7), .O(gate45inter4));
  nand2 gate594(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate595(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate596(.a(G5), .O(gate45inter7));
  inv1  gate597(.a(G272), .O(gate45inter8));
  nand2 gate598(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate599(.a(s_7), .b(gate45inter3), .O(gate45inter10));
  nor2  gate600(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate601(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate602(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate645(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate646(.a(gate59inter0), .b(s_14), .O(gate59inter1));
  and2  gate647(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate648(.a(s_14), .O(gate59inter3));
  inv1  gate649(.a(s_15), .O(gate59inter4));
  nand2 gate650(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate651(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate652(.a(G19), .O(gate59inter7));
  inv1  gate653(.a(G293), .O(gate59inter8));
  nand2 gate654(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate655(.a(s_15), .b(gate59inter3), .O(gate59inter10));
  nor2  gate656(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate657(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate658(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate743(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate744(.a(gate62inter0), .b(s_28), .O(gate62inter1));
  and2  gate745(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate746(.a(s_28), .O(gate62inter3));
  inv1  gate747(.a(s_29), .O(gate62inter4));
  nand2 gate748(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate749(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate750(.a(G22), .O(gate62inter7));
  inv1  gate751(.a(G296), .O(gate62inter8));
  nand2 gate752(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate753(.a(s_29), .b(gate62inter3), .O(gate62inter10));
  nor2  gate754(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate755(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate756(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1107(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1108(.a(gate63inter0), .b(s_80), .O(gate63inter1));
  and2  gate1109(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1110(.a(s_80), .O(gate63inter3));
  inv1  gate1111(.a(s_81), .O(gate63inter4));
  nand2 gate1112(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1113(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1114(.a(G23), .O(gate63inter7));
  inv1  gate1115(.a(G299), .O(gate63inter8));
  nand2 gate1116(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1117(.a(s_81), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1118(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1119(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1120(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1023(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1024(.a(gate71inter0), .b(s_68), .O(gate71inter1));
  and2  gate1025(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1026(.a(s_68), .O(gate71inter3));
  inv1  gate1027(.a(s_69), .O(gate71inter4));
  nand2 gate1028(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1029(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1030(.a(G31), .O(gate71inter7));
  inv1  gate1031(.a(G311), .O(gate71inter8));
  nand2 gate1032(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1033(.a(s_69), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1034(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1035(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1036(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1485(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1486(.a(gate72inter0), .b(s_134), .O(gate72inter1));
  and2  gate1487(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1488(.a(s_134), .O(gate72inter3));
  inv1  gate1489(.a(s_135), .O(gate72inter4));
  nand2 gate1490(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1491(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1492(.a(G32), .O(gate72inter7));
  inv1  gate1493(.a(G311), .O(gate72inter8));
  nand2 gate1494(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1495(.a(s_135), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1496(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1497(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1498(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1919(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1920(.a(gate76inter0), .b(s_196), .O(gate76inter1));
  and2  gate1921(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1922(.a(s_196), .O(gate76inter3));
  inv1  gate1923(.a(s_197), .O(gate76inter4));
  nand2 gate1924(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1925(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1926(.a(G13), .O(gate76inter7));
  inv1  gate1927(.a(G317), .O(gate76inter8));
  nand2 gate1928(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1929(.a(s_197), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1930(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1931(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1932(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1401(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1402(.a(gate77inter0), .b(s_122), .O(gate77inter1));
  and2  gate1403(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1404(.a(s_122), .O(gate77inter3));
  inv1  gate1405(.a(s_123), .O(gate77inter4));
  nand2 gate1406(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1407(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1408(.a(G2), .O(gate77inter7));
  inv1  gate1409(.a(G320), .O(gate77inter8));
  nand2 gate1410(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1411(.a(s_123), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1412(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1413(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1414(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1835(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1836(.a(gate78inter0), .b(s_184), .O(gate78inter1));
  and2  gate1837(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1838(.a(s_184), .O(gate78inter3));
  inv1  gate1839(.a(s_185), .O(gate78inter4));
  nand2 gate1840(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1841(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1842(.a(G6), .O(gate78inter7));
  inv1  gate1843(.a(G320), .O(gate78inter8));
  nand2 gate1844(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1845(.a(s_185), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1846(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1847(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1848(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate981(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate982(.a(gate81inter0), .b(s_62), .O(gate81inter1));
  and2  gate983(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate984(.a(s_62), .O(gate81inter3));
  inv1  gate985(.a(s_63), .O(gate81inter4));
  nand2 gate986(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate987(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate988(.a(G3), .O(gate81inter7));
  inv1  gate989(.a(G326), .O(gate81inter8));
  nand2 gate990(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate991(.a(s_63), .b(gate81inter3), .O(gate81inter10));
  nor2  gate992(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate993(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate994(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1723(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1724(.a(gate84inter0), .b(s_168), .O(gate84inter1));
  and2  gate1725(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1726(.a(s_168), .O(gate84inter3));
  inv1  gate1727(.a(s_169), .O(gate84inter4));
  nand2 gate1728(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1729(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1730(.a(G15), .O(gate84inter7));
  inv1  gate1731(.a(G329), .O(gate84inter8));
  nand2 gate1732(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1733(.a(s_169), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1734(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1735(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1736(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1331(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1332(.a(gate86inter0), .b(s_112), .O(gate86inter1));
  and2  gate1333(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1334(.a(s_112), .O(gate86inter3));
  inv1  gate1335(.a(s_113), .O(gate86inter4));
  nand2 gate1336(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1337(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1338(.a(G8), .O(gate86inter7));
  inv1  gate1339(.a(G332), .O(gate86inter8));
  nand2 gate1340(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1341(.a(s_113), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1342(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1343(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1344(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate729(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate730(.a(gate89inter0), .b(s_26), .O(gate89inter1));
  and2  gate731(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate732(.a(s_26), .O(gate89inter3));
  inv1  gate733(.a(s_27), .O(gate89inter4));
  nand2 gate734(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate735(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate736(.a(G17), .O(gate89inter7));
  inv1  gate737(.a(G338), .O(gate89inter8));
  nand2 gate738(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate739(.a(s_27), .b(gate89inter3), .O(gate89inter10));
  nor2  gate740(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate741(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate742(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1821(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1822(.a(gate93inter0), .b(s_182), .O(gate93inter1));
  and2  gate1823(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1824(.a(s_182), .O(gate93inter3));
  inv1  gate1825(.a(s_183), .O(gate93inter4));
  nand2 gate1826(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1827(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1828(.a(G18), .O(gate93inter7));
  inv1  gate1829(.a(G344), .O(gate93inter8));
  nand2 gate1830(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1831(.a(s_183), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1832(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1833(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1834(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate799(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate800(.a(gate94inter0), .b(s_36), .O(gate94inter1));
  and2  gate801(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate802(.a(s_36), .O(gate94inter3));
  inv1  gate803(.a(s_37), .O(gate94inter4));
  nand2 gate804(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate805(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate806(.a(G22), .O(gate94inter7));
  inv1  gate807(.a(G344), .O(gate94inter8));
  nand2 gate808(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate809(.a(s_37), .b(gate94inter3), .O(gate94inter10));
  nor2  gate810(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate811(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate812(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1877(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1878(.a(gate95inter0), .b(s_190), .O(gate95inter1));
  and2  gate1879(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1880(.a(s_190), .O(gate95inter3));
  inv1  gate1881(.a(s_191), .O(gate95inter4));
  nand2 gate1882(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1883(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1884(.a(G26), .O(gate95inter7));
  inv1  gate1885(.a(G347), .O(gate95inter8));
  nand2 gate1886(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1887(.a(s_191), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1888(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1889(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1890(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1695(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1696(.a(gate97inter0), .b(s_164), .O(gate97inter1));
  and2  gate1697(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1698(.a(s_164), .O(gate97inter3));
  inv1  gate1699(.a(s_165), .O(gate97inter4));
  nand2 gate1700(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1701(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1702(.a(G19), .O(gate97inter7));
  inv1  gate1703(.a(G350), .O(gate97inter8));
  nand2 gate1704(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1705(.a(s_165), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1706(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1707(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1708(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1079(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1080(.a(gate98inter0), .b(s_76), .O(gate98inter1));
  and2  gate1081(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1082(.a(s_76), .O(gate98inter3));
  inv1  gate1083(.a(s_77), .O(gate98inter4));
  nand2 gate1084(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1085(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1086(.a(G23), .O(gate98inter7));
  inv1  gate1087(.a(G350), .O(gate98inter8));
  nand2 gate1088(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1089(.a(s_77), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1090(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1091(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1092(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate673(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate674(.a(gate100inter0), .b(s_18), .O(gate100inter1));
  and2  gate675(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate676(.a(s_18), .O(gate100inter3));
  inv1  gate677(.a(s_19), .O(gate100inter4));
  nand2 gate678(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate679(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate680(.a(G31), .O(gate100inter7));
  inv1  gate681(.a(G353), .O(gate100inter8));
  nand2 gate682(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate683(.a(s_19), .b(gate100inter3), .O(gate100inter10));
  nor2  gate684(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate685(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate686(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate687(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate688(.a(gate105inter0), .b(s_20), .O(gate105inter1));
  and2  gate689(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate690(.a(s_20), .O(gate105inter3));
  inv1  gate691(.a(s_21), .O(gate105inter4));
  nand2 gate692(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate693(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate694(.a(G362), .O(gate105inter7));
  inv1  gate695(.a(G363), .O(gate105inter8));
  nand2 gate696(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate697(.a(s_21), .b(gate105inter3), .O(gate105inter10));
  nor2  gate698(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate699(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate700(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate701(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate702(.a(gate111inter0), .b(s_22), .O(gate111inter1));
  and2  gate703(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate704(.a(s_22), .O(gate111inter3));
  inv1  gate705(.a(s_23), .O(gate111inter4));
  nand2 gate706(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate707(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate708(.a(G374), .O(gate111inter7));
  inv1  gate709(.a(G375), .O(gate111inter8));
  nand2 gate710(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate711(.a(s_23), .b(gate111inter3), .O(gate111inter10));
  nor2  gate712(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate713(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate714(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1583(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1584(.a(gate113inter0), .b(s_148), .O(gate113inter1));
  and2  gate1585(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1586(.a(s_148), .O(gate113inter3));
  inv1  gate1587(.a(s_149), .O(gate113inter4));
  nand2 gate1588(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1589(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1590(.a(G378), .O(gate113inter7));
  inv1  gate1591(.a(G379), .O(gate113inter8));
  nand2 gate1592(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1593(.a(s_149), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1594(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1595(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1596(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate1261(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1262(.a(gate114inter0), .b(s_102), .O(gate114inter1));
  and2  gate1263(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1264(.a(s_102), .O(gate114inter3));
  inv1  gate1265(.a(s_103), .O(gate114inter4));
  nand2 gate1266(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1267(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1268(.a(G380), .O(gate114inter7));
  inv1  gate1269(.a(G381), .O(gate114inter8));
  nand2 gate1270(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1271(.a(s_103), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1272(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1273(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1274(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1681(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1682(.a(gate117inter0), .b(s_162), .O(gate117inter1));
  and2  gate1683(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1684(.a(s_162), .O(gate117inter3));
  inv1  gate1685(.a(s_163), .O(gate117inter4));
  nand2 gate1686(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1687(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1688(.a(G386), .O(gate117inter7));
  inv1  gate1689(.a(G387), .O(gate117inter8));
  nand2 gate1690(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1691(.a(s_163), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1692(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1693(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1694(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1317(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1318(.a(gate121inter0), .b(s_110), .O(gate121inter1));
  and2  gate1319(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1320(.a(s_110), .O(gate121inter3));
  inv1  gate1321(.a(s_111), .O(gate121inter4));
  nand2 gate1322(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1323(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1324(.a(G394), .O(gate121inter7));
  inv1  gate1325(.a(G395), .O(gate121inter8));
  nand2 gate1326(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1327(.a(s_111), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1328(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1329(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1330(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1065(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1066(.a(gate123inter0), .b(s_74), .O(gate123inter1));
  and2  gate1067(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1068(.a(s_74), .O(gate123inter3));
  inv1  gate1069(.a(s_75), .O(gate123inter4));
  nand2 gate1070(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1071(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1072(.a(G398), .O(gate123inter7));
  inv1  gate1073(.a(G399), .O(gate123inter8));
  nand2 gate1074(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1075(.a(s_75), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1076(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1077(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1078(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1387(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1388(.a(gate127inter0), .b(s_120), .O(gate127inter1));
  and2  gate1389(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1390(.a(s_120), .O(gate127inter3));
  inv1  gate1391(.a(s_121), .O(gate127inter4));
  nand2 gate1392(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1393(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1394(.a(G406), .O(gate127inter7));
  inv1  gate1395(.a(G407), .O(gate127inter8));
  nand2 gate1396(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1397(.a(s_121), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1398(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1399(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1400(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1051(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1052(.a(gate130inter0), .b(s_72), .O(gate130inter1));
  and2  gate1053(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1054(.a(s_72), .O(gate130inter3));
  inv1  gate1055(.a(s_73), .O(gate130inter4));
  nand2 gate1056(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1057(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1058(.a(G412), .O(gate130inter7));
  inv1  gate1059(.a(G413), .O(gate130inter8));
  nand2 gate1060(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1061(.a(s_73), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1062(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1063(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1064(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1345(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1346(.a(gate131inter0), .b(s_114), .O(gate131inter1));
  and2  gate1347(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1348(.a(s_114), .O(gate131inter3));
  inv1  gate1349(.a(s_115), .O(gate131inter4));
  nand2 gate1350(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1351(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1352(.a(G414), .O(gate131inter7));
  inv1  gate1353(.a(G415), .O(gate131inter8));
  nand2 gate1354(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1355(.a(s_115), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1356(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1357(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1358(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1457(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1458(.a(gate142inter0), .b(s_130), .O(gate142inter1));
  and2  gate1459(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1460(.a(s_130), .O(gate142inter3));
  inv1  gate1461(.a(s_131), .O(gate142inter4));
  nand2 gate1462(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1463(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1464(.a(G456), .O(gate142inter7));
  inv1  gate1465(.a(G459), .O(gate142inter8));
  nand2 gate1466(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1467(.a(s_131), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1468(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1469(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1470(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1121(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1122(.a(gate151inter0), .b(s_82), .O(gate151inter1));
  and2  gate1123(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1124(.a(s_82), .O(gate151inter3));
  inv1  gate1125(.a(s_83), .O(gate151inter4));
  nand2 gate1126(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1127(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1128(.a(G510), .O(gate151inter7));
  inv1  gate1129(.a(G513), .O(gate151inter8));
  nand2 gate1130(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1131(.a(s_83), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1132(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1133(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1134(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1611(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1612(.a(gate156inter0), .b(s_152), .O(gate156inter1));
  and2  gate1613(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1614(.a(s_152), .O(gate156inter3));
  inv1  gate1615(.a(s_153), .O(gate156inter4));
  nand2 gate1616(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1617(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1618(.a(G435), .O(gate156inter7));
  inv1  gate1619(.a(G525), .O(gate156inter8));
  nand2 gate1620(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1621(.a(s_153), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1622(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1623(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1624(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate757(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate758(.a(gate158inter0), .b(s_30), .O(gate158inter1));
  and2  gate759(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate760(.a(s_30), .O(gate158inter3));
  inv1  gate761(.a(s_31), .O(gate158inter4));
  nand2 gate762(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate763(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate764(.a(G441), .O(gate158inter7));
  inv1  gate765(.a(G528), .O(gate158inter8));
  nand2 gate766(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate767(.a(s_31), .b(gate158inter3), .O(gate158inter10));
  nor2  gate768(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate769(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate770(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1541(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1542(.a(gate160inter0), .b(s_142), .O(gate160inter1));
  and2  gate1543(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1544(.a(s_142), .O(gate160inter3));
  inv1  gate1545(.a(s_143), .O(gate160inter4));
  nand2 gate1546(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1547(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1548(.a(G447), .O(gate160inter7));
  inv1  gate1549(.a(G531), .O(gate160inter8));
  nand2 gate1550(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1551(.a(s_143), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1552(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1553(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1554(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate911(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate912(.a(gate166inter0), .b(s_52), .O(gate166inter1));
  and2  gate913(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate914(.a(s_52), .O(gate166inter3));
  inv1  gate915(.a(s_53), .O(gate166inter4));
  nand2 gate916(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate917(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate918(.a(G465), .O(gate166inter7));
  inv1  gate919(.a(G540), .O(gate166inter8));
  nand2 gate920(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate921(.a(s_53), .b(gate166inter3), .O(gate166inter10));
  nor2  gate922(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate923(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate924(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate575(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate576(.a(gate176inter0), .b(s_4), .O(gate176inter1));
  and2  gate577(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate578(.a(s_4), .O(gate176inter3));
  inv1  gate579(.a(s_5), .O(gate176inter4));
  nand2 gate580(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate581(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate582(.a(G495), .O(gate176inter7));
  inv1  gate583(.a(G555), .O(gate176inter8));
  nand2 gate584(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate585(.a(s_5), .b(gate176inter3), .O(gate176inter10));
  nor2  gate586(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate587(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate588(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate813(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate814(.a(gate178inter0), .b(s_38), .O(gate178inter1));
  and2  gate815(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate816(.a(s_38), .O(gate178inter3));
  inv1  gate817(.a(s_39), .O(gate178inter4));
  nand2 gate818(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate819(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate820(.a(G501), .O(gate178inter7));
  inv1  gate821(.a(G558), .O(gate178inter8));
  nand2 gate822(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate823(.a(s_39), .b(gate178inter3), .O(gate178inter10));
  nor2  gate824(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate825(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate826(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1751(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1752(.a(gate189inter0), .b(s_172), .O(gate189inter1));
  and2  gate1753(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1754(.a(s_172), .O(gate189inter3));
  inv1  gate1755(.a(s_173), .O(gate189inter4));
  nand2 gate1756(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1757(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1758(.a(G578), .O(gate189inter7));
  inv1  gate1759(.a(G579), .O(gate189inter8));
  nand2 gate1760(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1761(.a(s_173), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1762(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1763(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1764(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1527(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1528(.a(gate190inter0), .b(s_140), .O(gate190inter1));
  and2  gate1529(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1530(.a(s_140), .O(gate190inter3));
  inv1  gate1531(.a(s_141), .O(gate190inter4));
  nand2 gate1532(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1533(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1534(.a(G580), .O(gate190inter7));
  inv1  gate1535(.a(G581), .O(gate190inter8));
  nand2 gate1536(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1537(.a(s_141), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1538(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1539(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1540(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate771(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate772(.a(gate191inter0), .b(s_32), .O(gate191inter1));
  and2  gate773(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate774(.a(s_32), .O(gate191inter3));
  inv1  gate775(.a(s_33), .O(gate191inter4));
  nand2 gate776(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate777(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate778(.a(G582), .O(gate191inter7));
  inv1  gate779(.a(G583), .O(gate191inter8));
  nand2 gate780(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate781(.a(s_33), .b(gate191inter3), .O(gate191inter10));
  nor2  gate782(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate783(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate784(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate785(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate786(.a(gate192inter0), .b(s_34), .O(gate192inter1));
  and2  gate787(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate788(.a(s_34), .O(gate192inter3));
  inv1  gate789(.a(s_35), .O(gate192inter4));
  nand2 gate790(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate791(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate792(.a(G584), .O(gate192inter7));
  inv1  gate793(.a(G585), .O(gate192inter8));
  nand2 gate794(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate795(.a(s_35), .b(gate192inter3), .O(gate192inter10));
  nor2  gate796(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate797(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate798(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1009(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1010(.a(gate194inter0), .b(s_66), .O(gate194inter1));
  and2  gate1011(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1012(.a(s_66), .O(gate194inter3));
  inv1  gate1013(.a(s_67), .O(gate194inter4));
  nand2 gate1014(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1015(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1016(.a(G588), .O(gate194inter7));
  inv1  gate1017(.a(G589), .O(gate194inter8));
  nand2 gate1018(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1019(.a(s_67), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1020(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1021(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1022(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1359(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1360(.a(gate197inter0), .b(s_116), .O(gate197inter1));
  and2  gate1361(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1362(.a(s_116), .O(gate197inter3));
  inv1  gate1363(.a(s_117), .O(gate197inter4));
  nand2 gate1364(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1365(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1366(.a(G594), .O(gate197inter7));
  inv1  gate1367(.a(G595), .O(gate197inter8));
  nand2 gate1368(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1369(.a(s_117), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1370(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1371(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1372(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate715(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate716(.a(gate204inter0), .b(s_24), .O(gate204inter1));
  and2  gate717(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate718(.a(s_24), .O(gate204inter3));
  inv1  gate719(.a(s_25), .O(gate204inter4));
  nand2 gate720(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate721(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate722(.a(G607), .O(gate204inter7));
  inv1  gate723(.a(G617), .O(gate204inter8));
  nand2 gate724(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate725(.a(s_25), .b(gate204inter3), .O(gate204inter10));
  nor2  gate726(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate727(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate728(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1891(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1892(.a(gate206inter0), .b(s_192), .O(gate206inter1));
  and2  gate1893(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1894(.a(s_192), .O(gate206inter3));
  inv1  gate1895(.a(s_193), .O(gate206inter4));
  nand2 gate1896(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1897(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1898(.a(G632), .O(gate206inter7));
  inv1  gate1899(.a(G637), .O(gate206inter8));
  nand2 gate1900(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1901(.a(s_193), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1902(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1903(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1904(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate603(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate604(.a(gate208inter0), .b(s_8), .O(gate208inter1));
  and2  gate605(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate606(.a(s_8), .O(gate208inter3));
  inv1  gate607(.a(s_9), .O(gate208inter4));
  nand2 gate608(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate609(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate610(.a(G627), .O(gate208inter7));
  inv1  gate611(.a(G637), .O(gate208inter8));
  nand2 gate612(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate613(.a(s_9), .b(gate208inter3), .O(gate208inter10));
  nor2  gate614(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate615(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate616(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1205(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1206(.a(gate209inter0), .b(s_94), .O(gate209inter1));
  and2  gate1207(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1208(.a(s_94), .O(gate209inter3));
  inv1  gate1209(.a(s_95), .O(gate209inter4));
  nand2 gate1210(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1211(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1212(.a(G602), .O(gate209inter7));
  inv1  gate1213(.a(G666), .O(gate209inter8));
  nand2 gate1214(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1215(.a(s_95), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1216(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1217(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1218(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1947(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1948(.a(gate211inter0), .b(s_200), .O(gate211inter1));
  and2  gate1949(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1950(.a(s_200), .O(gate211inter3));
  inv1  gate1951(.a(s_201), .O(gate211inter4));
  nand2 gate1952(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1953(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1954(.a(G612), .O(gate211inter7));
  inv1  gate1955(.a(G669), .O(gate211inter8));
  nand2 gate1956(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1957(.a(s_201), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1958(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1959(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1960(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1905(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1906(.a(gate212inter0), .b(s_194), .O(gate212inter1));
  and2  gate1907(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1908(.a(s_194), .O(gate212inter3));
  inv1  gate1909(.a(s_195), .O(gate212inter4));
  nand2 gate1910(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1911(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1912(.a(G617), .O(gate212inter7));
  inv1  gate1913(.a(G669), .O(gate212inter8));
  nand2 gate1914(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1915(.a(s_195), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1916(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1917(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1918(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1779(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1780(.a(gate213inter0), .b(s_176), .O(gate213inter1));
  and2  gate1781(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1782(.a(s_176), .O(gate213inter3));
  inv1  gate1783(.a(s_177), .O(gate213inter4));
  nand2 gate1784(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1785(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1786(.a(G602), .O(gate213inter7));
  inv1  gate1787(.a(G672), .O(gate213inter8));
  nand2 gate1788(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1789(.a(s_177), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1790(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1791(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1792(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1513(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1514(.a(gate215inter0), .b(s_138), .O(gate215inter1));
  and2  gate1515(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1516(.a(s_138), .O(gate215inter3));
  inv1  gate1517(.a(s_139), .O(gate215inter4));
  nand2 gate1518(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1519(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1520(.a(G607), .O(gate215inter7));
  inv1  gate1521(.a(G675), .O(gate215inter8));
  nand2 gate1522(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1523(.a(s_139), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1524(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1525(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1526(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1667(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1668(.a(gate221inter0), .b(s_160), .O(gate221inter1));
  and2  gate1669(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1670(.a(s_160), .O(gate221inter3));
  inv1  gate1671(.a(s_161), .O(gate221inter4));
  nand2 gate1672(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1673(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1674(.a(G622), .O(gate221inter7));
  inv1  gate1675(.a(G684), .O(gate221inter8));
  nand2 gate1676(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1677(.a(s_161), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1678(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1679(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1680(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1807(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1808(.a(gate223inter0), .b(s_180), .O(gate223inter1));
  and2  gate1809(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1810(.a(s_180), .O(gate223inter3));
  inv1  gate1811(.a(s_181), .O(gate223inter4));
  nand2 gate1812(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1813(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1814(.a(G627), .O(gate223inter7));
  inv1  gate1815(.a(G687), .O(gate223inter8));
  nand2 gate1816(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1817(.a(s_181), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1818(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1819(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1820(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1177(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1178(.a(gate227inter0), .b(s_90), .O(gate227inter1));
  and2  gate1179(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1180(.a(s_90), .O(gate227inter3));
  inv1  gate1181(.a(s_91), .O(gate227inter4));
  nand2 gate1182(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1183(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1184(.a(G694), .O(gate227inter7));
  inv1  gate1185(.a(G695), .O(gate227inter8));
  nand2 gate1186(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1187(.a(s_91), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1188(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1189(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1190(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1499(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1500(.a(gate231inter0), .b(s_136), .O(gate231inter1));
  and2  gate1501(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1502(.a(s_136), .O(gate231inter3));
  inv1  gate1503(.a(s_137), .O(gate231inter4));
  nand2 gate1504(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1505(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1506(.a(G702), .O(gate231inter7));
  inv1  gate1507(.a(G703), .O(gate231inter8));
  nand2 gate1508(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1509(.a(s_137), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1510(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1511(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1512(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1639(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1640(.a(gate237inter0), .b(s_156), .O(gate237inter1));
  and2  gate1641(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1642(.a(s_156), .O(gate237inter3));
  inv1  gate1643(.a(s_157), .O(gate237inter4));
  nand2 gate1644(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1645(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1646(.a(G254), .O(gate237inter7));
  inv1  gate1647(.a(G706), .O(gate237inter8));
  nand2 gate1648(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1649(.a(s_157), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1650(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1651(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1652(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1569(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1570(.a(gate240inter0), .b(s_146), .O(gate240inter1));
  and2  gate1571(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1572(.a(s_146), .O(gate240inter3));
  inv1  gate1573(.a(s_147), .O(gate240inter4));
  nand2 gate1574(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1575(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1576(.a(G263), .O(gate240inter7));
  inv1  gate1577(.a(G715), .O(gate240inter8));
  nand2 gate1578(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1579(.a(s_147), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1580(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1581(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1582(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate953(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate954(.a(gate243inter0), .b(s_58), .O(gate243inter1));
  and2  gate955(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate956(.a(s_58), .O(gate243inter3));
  inv1  gate957(.a(s_59), .O(gate243inter4));
  nand2 gate958(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate959(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate960(.a(G245), .O(gate243inter7));
  inv1  gate961(.a(G733), .O(gate243inter8));
  nand2 gate962(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate963(.a(s_59), .b(gate243inter3), .O(gate243inter10));
  nor2  gate964(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate965(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate966(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate617(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate618(.a(gate247inter0), .b(s_10), .O(gate247inter1));
  and2  gate619(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate620(.a(s_10), .O(gate247inter3));
  inv1  gate621(.a(s_11), .O(gate247inter4));
  nand2 gate622(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate623(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate624(.a(G251), .O(gate247inter7));
  inv1  gate625(.a(G739), .O(gate247inter8));
  nand2 gate626(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate627(.a(s_11), .b(gate247inter3), .O(gate247inter10));
  nor2  gate628(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate629(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate630(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1765(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1766(.a(gate250inter0), .b(s_174), .O(gate250inter1));
  and2  gate1767(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1768(.a(s_174), .O(gate250inter3));
  inv1  gate1769(.a(s_175), .O(gate250inter4));
  nand2 gate1770(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1771(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1772(.a(G706), .O(gate250inter7));
  inv1  gate1773(.a(G742), .O(gate250inter8));
  nand2 gate1774(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1775(.a(s_175), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1776(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1777(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1778(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1471(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1472(.a(gate251inter0), .b(s_132), .O(gate251inter1));
  and2  gate1473(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1474(.a(s_132), .O(gate251inter3));
  inv1  gate1475(.a(s_133), .O(gate251inter4));
  nand2 gate1476(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1477(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1478(.a(G257), .O(gate251inter7));
  inv1  gate1479(.a(G745), .O(gate251inter8));
  nand2 gate1480(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1481(.a(s_133), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1482(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1483(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1484(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1793(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1794(.a(gate253inter0), .b(s_178), .O(gate253inter1));
  and2  gate1795(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1796(.a(s_178), .O(gate253inter3));
  inv1  gate1797(.a(s_179), .O(gate253inter4));
  nand2 gate1798(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1799(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1800(.a(G260), .O(gate253inter7));
  inv1  gate1801(.a(G748), .O(gate253inter8));
  nand2 gate1802(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1803(.a(s_179), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1804(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1805(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1806(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate925(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate926(.a(gate257inter0), .b(s_54), .O(gate257inter1));
  and2  gate927(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate928(.a(s_54), .O(gate257inter3));
  inv1  gate929(.a(s_55), .O(gate257inter4));
  nand2 gate930(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate931(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate932(.a(G754), .O(gate257inter7));
  inv1  gate933(.a(G755), .O(gate257inter8));
  nand2 gate934(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate935(.a(s_55), .b(gate257inter3), .O(gate257inter10));
  nor2  gate936(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate937(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate938(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1415(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1416(.a(gate261inter0), .b(s_124), .O(gate261inter1));
  and2  gate1417(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1418(.a(s_124), .O(gate261inter3));
  inv1  gate1419(.a(s_125), .O(gate261inter4));
  nand2 gate1420(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1421(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1422(.a(G762), .O(gate261inter7));
  inv1  gate1423(.a(G763), .O(gate261inter8));
  nand2 gate1424(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1425(.a(s_125), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1426(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1427(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1428(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate897(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate898(.a(gate265inter0), .b(s_50), .O(gate265inter1));
  and2  gate899(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate900(.a(s_50), .O(gate265inter3));
  inv1  gate901(.a(s_51), .O(gate265inter4));
  nand2 gate902(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate903(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate904(.a(G642), .O(gate265inter7));
  inv1  gate905(.a(G770), .O(gate265inter8));
  nand2 gate906(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate907(.a(s_51), .b(gate265inter3), .O(gate265inter10));
  nor2  gate908(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate909(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate910(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate841(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate842(.a(gate267inter0), .b(s_42), .O(gate267inter1));
  and2  gate843(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate844(.a(s_42), .O(gate267inter3));
  inv1  gate845(.a(s_43), .O(gate267inter4));
  nand2 gate846(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate847(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate848(.a(G648), .O(gate267inter7));
  inv1  gate849(.a(G776), .O(gate267inter8));
  nand2 gate850(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate851(.a(s_43), .b(gate267inter3), .O(gate267inter10));
  nor2  gate852(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate853(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate854(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate883(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate884(.a(gate272inter0), .b(s_48), .O(gate272inter1));
  and2  gate885(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate886(.a(s_48), .O(gate272inter3));
  inv1  gate887(.a(s_49), .O(gate272inter4));
  nand2 gate888(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate889(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate890(.a(G663), .O(gate272inter7));
  inv1  gate891(.a(G791), .O(gate272inter8));
  nand2 gate892(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate893(.a(s_49), .b(gate272inter3), .O(gate272inter10));
  nor2  gate894(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate895(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate896(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1373(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1374(.a(gate276inter0), .b(s_118), .O(gate276inter1));
  and2  gate1375(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1376(.a(s_118), .O(gate276inter3));
  inv1  gate1377(.a(s_119), .O(gate276inter4));
  nand2 gate1378(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1379(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1380(.a(G773), .O(gate276inter7));
  inv1  gate1381(.a(G797), .O(gate276inter8));
  nand2 gate1382(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1383(.a(s_119), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1384(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1385(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1386(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1961(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1962(.a(gate281inter0), .b(s_202), .O(gate281inter1));
  and2  gate1963(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1964(.a(s_202), .O(gate281inter3));
  inv1  gate1965(.a(s_203), .O(gate281inter4));
  nand2 gate1966(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1967(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1968(.a(G654), .O(gate281inter7));
  inv1  gate1969(.a(G806), .O(gate281inter8));
  nand2 gate1970(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1971(.a(s_203), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1972(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1973(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1974(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1863(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1864(.a(gate283inter0), .b(s_188), .O(gate283inter1));
  and2  gate1865(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1866(.a(s_188), .O(gate283inter3));
  inv1  gate1867(.a(s_189), .O(gate283inter4));
  nand2 gate1868(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1869(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1870(.a(G657), .O(gate283inter7));
  inv1  gate1871(.a(G809), .O(gate283inter8));
  nand2 gate1872(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1873(.a(s_189), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1874(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1875(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1876(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate631(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate632(.a(gate286inter0), .b(s_12), .O(gate286inter1));
  and2  gate633(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate634(.a(s_12), .O(gate286inter3));
  inv1  gate635(.a(s_13), .O(gate286inter4));
  nand2 gate636(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate637(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate638(.a(G788), .O(gate286inter7));
  inv1  gate639(.a(G812), .O(gate286inter8));
  nand2 gate640(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate641(.a(s_13), .b(gate286inter3), .O(gate286inter10));
  nor2  gate642(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate643(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate644(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1233(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1234(.a(gate296inter0), .b(s_98), .O(gate296inter1));
  and2  gate1235(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1236(.a(s_98), .O(gate296inter3));
  inv1  gate1237(.a(s_99), .O(gate296inter4));
  nand2 gate1238(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1239(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1240(.a(G826), .O(gate296inter7));
  inv1  gate1241(.a(G827), .O(gate296inter8));
  nand2 gate1242(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1243(.a(s_99), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1244(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1245(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1246(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1737(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1738(.a(gate398inter0), .b(s_170), .O(gate398inter1));
  and2  gate1739(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1740(.a(s_170), .O(gate398inter3));
  inv1  gate1741(.a(s_171), .O(gate398inter4));
  nand2 gate1742(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1743(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1744(.a(G12), .O(gate398inter7));
  inv1  gate1745(.a(G1069), .O(gate398inter8));
  nand2 gate1746(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1747(.a(s_171), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1748(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1749(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1750(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1093(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1094(.a(gate417inter0), .b(s_78), .O(gate417inter1));
  and2  gate1095(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1096(.a(s_78), .O(gate417inter3));
  inv1  gate1097(.a(s_79), .O(gate417inter4));
  nand2 gate1098(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1099(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1100(.a(G31), .O(gate417inter7));
  inv1  gate1101(.a(G1126), .O(gate417inter8));
  nand2 gate1102(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1103(.a(s_79), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1104(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1105(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1106(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1163(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1164(.a(gate418inter0), .b(s_88), .O(gate418inter1));
  and2  gate1165(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1166(.a(s_88), .O(gate418inter3));
  inv1  gate1167(.a(s_89), .O(gate418inter4));
  nand2 gate1168(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1169(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1170(.a(G32), .O(gate418inter7));
  inv1  gate1171(.a(G1129), .O(gate418inter8));
  nand2 gate1172(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1173(.a(s_89), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1174(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1175(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1176(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate995(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate996(.a(gate421inter0), .b(s_64), .O(gate421inter1));
  and2  gate997(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate998(.a(s_64), .O(gate421inter3));
  inv1  gate999(.a(s_65), .O(gate421inter4));
  nand2 gate1000(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1001(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1002(.a(G2), .O(gate421inter7));
  inv1  gate1003(.a(G1135), .O(gate421inter8));
  nand2 gate1004(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1005(.a(s_65), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1006(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1007(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1008(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1597(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1598(.a(gate422inter0), .b(s_150), .O(gate422inter1));
  and2  gate1599(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1600(.a(s_150), .O(gate422inter3));
  inv1  gate1601(.a(s_151), .O(gate422inter4));
  nand2 gate1602(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1603(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1604(.a(G1039), .O(gate422inter7));
  inv1  gate1605(.a(G1135), .O(gate422inter8));
  nand2 gate1606(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1607(.a(s_151), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1608(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1609(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1610(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1653(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1654(.a(gate424inter0), .b(s_158), .O(gate424inter1));
  and2  gate1655(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1656(.a(s_158), .O(gate424inter3));
  inv1  gate1657(.a(s_159), .O(gate424inter4));
  nand2 gate1658(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1659(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1660(.a(G1042), .O(gate424inter7));
  inv1  gate1661(.a(G1138), .O(gate424inter8));
  nand2 gate1662(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1663(.a(s_159), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1664(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1665(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1666(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1429(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1430(.a(gate425inter0), .b(s_126), .O(gate425inter1));
  and2  gate1431(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1432(.a(s_126), .O(gate425inter3));
  inv1  gate1433(.a(s_127), .O(gate425inter4));
  nand2 gate1434(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1435(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1436(.a(G4), .O(gate425inter7));
  inv1  gate1437(.a(G1141), .O(gate425inter8));
  nand2 gate1438(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1439(.a(s_127), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1440(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1441(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1442(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate869(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate870(.a(gate430inter0), .b(s_46), .O(gate430inter1));
  and2  gate871(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate872(.a(s_46), .O(gate430inter3));
  inv1  gate873(.a(s_47), .O(gate430inter4));
  nand2 gate874(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate875(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate876(.a(G1051), .O(gate430inter7));
  inv1  gate877(.a(G1147), .O(gate430inter8));
  nand2 gate878(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate879(.a(s_47), .b(gate430inter3), .O(gate430inter10));
  nor2  gate880(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate881(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate882(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1219(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1220(.a(gate433inter0), .b(s_96), .O(gate433inter1));
  and2  gate1221(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1222(.a(s_96), .O(gate433inter3));
  inv1  gate1223(.a(s_97), .O(gate433inter4));
  nand2 gate1224(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1225(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1226(.a(G8), .O(gate433inter7));
  inv1  gate1227(.a(G1153), .O(gate433inter8));
  nand2 gate1228(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1229(.a(s_97), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1230(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1231(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1232(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1975(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1976(.a(gate436inter0), .b(s_204), .O(gate436inter1));
  and2  gate1977(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1978(.a(s_204), .O(gate436inter3));
  inv1  gate1979(.a(s_205), .O(gate436inter4));
  nand2 gate1980(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1981(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1982(.a(G1060), .O(gate436inter7));
  inv1  gate1983(.a(G1156), .O(gate436inter8));
  nand2 gate1984(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1985(.a(s_205), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1986(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1987(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1988(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1247(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1248(.a(gate441inter0), .b(s_100), .O(gate441inter1));
  and2  gate1249(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1250(.a(s_100), .O(gate441inter3));
  inv1  gate1251(.a(s_101), .O(gate441inter4));
  nand2 gate1252(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1253(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1254(.a(G12), .O(gate441inter7));
  inv1  gate1255(.a(G1165), .O(gate441inter8));
  nand2 gate1256(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1257(.a(s_101), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1258(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1259(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1260(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1191(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1192(.a(gate442inter0), .b(s_92), .O(gate442inter1));
  and2  gate1193(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1194(.a(s_92), .O(gate442inter3));
  inv1  gate1195(.a(s_93), .O(gate442inter4));
  nand2 gate1196(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1197(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1198(.a(G1069), .O(gate442inter7));
  inv1  gate1199(.a(G1165), .O(gate442inter8));
  nand2 gate1200(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1201(.a(s_93), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1202(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1203(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1204(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1303(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1304(.a(gate444inter0), .b(s_108), .O(gate444inter1));
  and2  gate1305(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1306(.a(s_108), .O(gate444inter3));
  inv1  gate1307(.a(s_109), .O(gate444inter4));
  nand2 gate1308(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1309(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1310(.a(G1072), .O(gate444inter7));
  inv1  gate1311(.a(G1168), .O(gate444inter8));
  nand2 gate1312(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1313(.a(s_109), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1314(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1315(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1316(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1037(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1038(.a(gate456inter0), .b(s_70), .O(gate456inter1));
  and2  gate1039(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1040(.a(s_70), .O(gate456inter3));
  inv1  gate1041(.a(s_71), .O(gate456inter4));
  nand2 gate1042(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1043(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1044(.a(G1090), .O(gate456inter7));
  inv1  gate1045(.a(G1186), .O(gate456inter8));
  nand2 gate1046(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1047(.a(s_71), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1048(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1049(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1050(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1625(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1626(.a(gate459inter0), .b(s_154), .O(gate459inter1));
  and2  gate1627(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1628(.a(s_154), .O(gate459inter3));
  inv1  gate1629(.a(s_155), .O(gate459inter4));
  nand2 gate1630(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1631(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1632(.a(G21), .O(gate459inter7));
  inv1  gate1633(.a(G1192), .O(gate459inter8));
  nand2 gate1634(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1635(.a(s_155), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1636(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1637(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1638(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate967(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate968(.a(gate460inter0), .b(s_60), .O(gate460inter1));
  and2  gate969(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate970(.a(s_60), .O(gate460inter3));
  inv1  gate971(.a(s_61), .O(gate460inter4));
  nand2 gate972(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate973(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate974(.a(G1096), .O(gate460inter7));
  inv1  gate975(.a(G1192), .O(gate460inter8));
  nand2 gate976(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate977(.a(s_61), .b(gate460inter3), .O(gate460inter10));
  nor2  gate978(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate979(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate980(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate827(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate828(.a(gate461inter0), .b(s_40), .O(gate461inter1));
  and2  gate829(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate830(.a(s_40), .O(gate461inter3));
  inv1  gate831(.a(s_41), .O(gate461inter4));
  nand2 gate832(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate833(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate834(.a(G22), .O(gate461inter7));
  inv1  gate835(.a(G1195), .O(gate461inter8));
  nand2 gate836(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate837(.a(s_41), .b(gate461inter3), .O(gate461inter10));
  nor2  gate838(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate839(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate840(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1849(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1850(.a(gate463inter0), .b(s_186), .O(gate463inter1));
  and2  gate1851(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1852(.a(s_186), .O(gate463inter3));
  inv1  gate1853(.a(s_187), .O(gate463inter4));
  nand2 gate1854(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1855(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1856(.a(G23), .O(gate463inter7));
  inv1  gate1857(.a(G1198), .O(gate463inter8));
  nand2 gate1858(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1859(.a(s_187), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1860(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1861(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1862(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1933(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1934(.a(gate465inter0), .b(s_198), .O(gate465inter1));
  and2  gate1935(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1936(.a(s_198), .O(gate465inter3));
  inv1  gate1937(.a(s_199), .O(gate465inter4));
  nand2 gate1938(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1939(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1940(.a(G24), .O(gate465inter7));
  inv1  gate1941(.a(G1201), .O(gate465inter8));
  nand2 gate1942(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1943(.a(s_199), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1944(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1945(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1946(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1135(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1136(.a(gate466inter0), .b(s_84), .O(gate466inter1));
  and2  gate1137(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1138(.a(s_84), .O(gate466inter3));
  inv1  gate1139(.a(s_85), .O(gate466inter4));
  nand2 gate1140(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1141(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1142(.a(G1105), .O(gate466inter7));
  inv1  gate1143(.a(G1201), .O(gate466inter8));
  nand2 gate1144(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1145(.a(s_85), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1146(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1147(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1148(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate659(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate660(.a(gate480inter0), .b(s_16), .O(gate480inter1));
  and2  gate661(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate662(.a(s_16), .O(gate480inter3));
  inv1  gate663(.a(s_17), .O(gate480inter4));
  nand2 gate664(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate665(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate666(.a(G1126), .O(gate480inter7));
  inv1  gate667(.a(G1222), .O(gate480inter8));
  nand2 gate668(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate669(.a(s_17), .b(gate480inter3), .O(gate480inter10));
  nor2  gate670(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate671(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate672(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1443(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1444(.a(gate486inter0), .b(s_128), .O(gate486inter1));
  and2  gate1445(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1446(.a(s_128), .O(gate486inter3));
  inv1  gate1447(.a(s_129), .O(gate486inter4));
  nand2 gate1448(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1449(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1450(.a(G1234), .O(gate486inter7));
  inv1  gate1451(.a(G1235), .O(gate486inter8));
  nand2 gate1452(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1453(.a(s_129), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1454(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1455(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1456(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1289(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1290(.a(gate499inter0), .b(s_106), .O(gate499inter1));
  and2  gate1291(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1292(.a(s_106), .O(gate499inter3));
  inv1  gate1293(.a(s_107), .O(gate499inter4));
  nand2 gate1294(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1295(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1296(.a(G1260), .O(gate499inter7));
  inv1  gate1297(.a(G1261), .O(gate499inter8));
  nand2 gate1298(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1299(.a(s_107), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1300(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1301(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1302(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1149(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1150(.a(gate501inter0), .b(s_86), .O(gate501inter1));
  and2  gate1151(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1152(.a(s_86), .O(gate501inter3));
  inv1  gate1153(.a(s_87), .O(gate501inter4));
  nand2 gate1154(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1155(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1156(.a(G1264), .O(gate501inter7));
  inv1  gate1157(.a(G1265), .O(gate501inter8));
  nand2 gate1158(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1159(.a(s_87), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1160(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1161(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1162(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate561(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate562(.a(gate502inter0), .b(s_2), .O(gate502inter1));
  and2  gate563(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate564(.a(s_2), .O(gate502inter3));
  inv1  gate565(.a(s_3), .O(gate502inter4));
  nand2 gate566(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate567(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate568(.a(G1266), .O(gate502inter7));
  inv1  gate569(.a(G1267), .O(gate502inter8));
  nand2 gate570(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate571(.a(s_3), .b(gate502inter3), .O(gate502inter10));
  nor2  gate572(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate573(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate574(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1555(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1556(.a(gate504inter0), .b(s_144), .O(gate504inter1));
  and2  gate1557(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1558(.a(s_144), .O(gate504inter3));
  inv1  gate1559(.a(s_145), .O(gate504inter4));
  nand2 gate1560(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1561(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1562(.a(G1270), .O(gate504inter7));
  inv1  gate1563(.a(G1271), .O(gate504inter8));
  nand2 gate1564(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1565(.a(s_145), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1566(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1567(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1568(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2017(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2018(.a(gate513inter0), .b(s_210), .O(gate513inter1));
  and2  gate2019(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2020(.a(s_210), .O(gate513inter3));
  inv1  gate2021(.a(s_211), .O(gate513inter4));
  nand2 gate2022(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2023(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2024(.a(G1288), .O(gate513inter7));
  inv1  gate2025(.a(G1289), .O(gate513inter8));
  nand2 gate2026(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2027(.a(s_211), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2028(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2029(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2030(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule