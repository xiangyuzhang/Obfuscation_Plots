module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1597(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1598(.a(gate11inter0), .b(s_150), .O(gate11inter1));
  and2  gate1599(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1600(.a(s_150), .O(gate11inter3));
  inv1  gate1601(.a(s_151), .O(gate11inter4));
  nand2 gate1602(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1603(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1604(.a(G5), .O(gate11inter7));
  inv1  gate1605(.a(G6), .O(gate11inter8));
  nand2 gate1606(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1607(.a(s_151), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1608(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1609(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1610(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1513(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1514(.a(gate19inter0), .b(s_138), .O(gate19inter1));
  and2  gate1515(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1516(.a(s_138), .O(gate19inter3));
  inv1  gate1517(.a(s_139), .O(gate19inter4));
  nand2 gate1518(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1519(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1520(.a(G21), .O(gate19inter7));
  inv1  gate1521(.a(G22), .O(gate19inter8));
  nand2 gate1522(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1523(.a(s_139), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1524(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1525(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1526(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1107(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1108(.a(gate22inter0), .b(s_80), .O(gate22inter1));
  and2  gate1109(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1110(.a(s_80), .O(gate22inter3));
  inv1  gate1111(.a(s_81), .O(gate22inter4));
  nand2 gate1112(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1113(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1114(.a(G27), .O(gate22inter7));
  inv1  gate1115(.a(G28), .O(gate22inter8));
  nand2 gate1116(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1117(.a(s_81), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1118(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1119(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1120(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1289(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1290(.a(gate25inter0), .b(s_106), .O(gate25inter1));
  and2  gate1291(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1292(.a(s_106), .O(gate25inter3));
  inv1  gate1293(.a(s_107), .O(gate25inter4));
  nand2 gate1294(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1295(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1296(.a(G1), .O(gate25inter7));
  inv1  gate1297(.a(G5), .O(gate25inter8));
  nand2 gate1298(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1299(.a(s_107), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1300(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1301(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1302(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1541(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1542(.a(gate28inter0), .b(s_142), .O(gate28inter1));
  and2  gate1543(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1544(.a(s_142), .O(gate28inter3));
  inv1  gate1545(.a(s_143), .O(gate28inter4));
  nand2 gate1546(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1547(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1548(.a(G10), .O(gate28inter7));
  inv1  gate1549(.a(G14), .O(gate28inter8));
  nand2 gate1550(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1551(.a(s_143), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1552(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1553(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1554(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1471(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1472(.a(gate33inter0), .b(s_132), .O(gate33inter1));
  and2  gate1473(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1474(.a(s_132), .O(gate33inter3));
  inv1  gate1475(.a(s_133), .O(gate33inter4));
  nand2 gate1476(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1477(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1478(.a(G17), .O(gate33inter7));
  inv1  gate1479(.a(G21), .O(gate33inter8));
  nand2 gate1480(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1481(.a(s_133), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1482(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1483(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1484(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1177(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1178(.a(gate34inter0), .b(s_90), .O(gate34inter1));
  and2  gate1179(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1180(.a(s_90), .O(gate34inter3));
  inv1  gate1181(.a(s_91), .O(gate34inter4));
  nand2 gate1182(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1183(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1184(.a(G25), .O(gate34inter7));
  inv1  gate1185(.a(G29), .O(gate34inter8));
  nand2 gate1186(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1187(.a(s_91), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1188(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1189(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1190(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate631(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate632(.a(gate40inter0), .b(s_12), .O(gate40inter1));
  and2  gate633(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate634(.a(s_12), .O(gate40inter3));
  inv1  gate635(.a(s_13), .O(gate40inter4));
  nand2 gate636(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate637(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate638(.a(G28), .O(gate40inter7));
  inv1  gate639(.a(G32), .O(gate40inter8));
  nand2 gate640(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate641(.a(s_13), .b(gate40inter3), .O(gate40inter10));
  nor2  gate642(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate643(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate644(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1625(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1626(.a(gate49inter0), .b(s_154), .O(gate49inter1));
  and2  gate1627(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1628(.a(s_154), .O(gate49inter3));
  inv1  gate1629(.a(s_155), .O(gate49inter4));
  nand2 gate1630(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1631(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1632(.a(G9), .O(gate49inter7));
  inv1  gate1633(.a(G278), .O(gate49inter8));
  nand2 gate1634(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1635(.a(s_155), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1636(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1637(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1638(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate981(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate982(.a(gate56inter0), .b(s_62), .O(gate56inter1));
  and2  gate983(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate984(.a(s_62), .O(gate56inter3));
  inv1  gate985(.a(s_63), .O(gate56inter4));
  nand2 gate986(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate987(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate988(.a(G16), .O(gate56inter7));
  inv1  gate989(.a(G287), .O(gate56inter8));
  nand2 gate990(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate991(.a(s_63), .b(gate56inter3), .O(gate56inter10));
  nor2  gate992(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate993(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate994(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1247(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1248(.a(gate58inter0), .b(s_100), .O(gate58inter1));
  and2  gate1249(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1250(.a(s_100), .O(gate58inter3));
  inv1  gate1251(.a(s_101), .O(gate58inter4));
  nand2 gate1252(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1253(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1254(.a(G18), .O(gate58inter7));
  inv1  gate1255(.a(G290), .O(gate58inter8));
  nand2 gate1256(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1257(.a(s_101), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1258(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1259(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1260(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1163(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1164(.a(gate64inter0), .b(s_88), .O(gate64inter1));
  and2  gate1165(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1166(.a(s_88), .O(gate64inter3));
  inv1  gate1167(.a(s_89), .O(gate64inter4));
  nand2 gate1168(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1169(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1170(.a(G24), .O(gate64inter7));
  inv1  gate1171(.a(G299), .O(gate64inter8));
  nand2 gate1172(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1173(.a(s_89), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1174(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1175(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1176(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1219(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1220(.a(gate66inter0), .b(s_96), .O(gate66inter1));
  and2  gate1221(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1222(.a(s_96), .O(gate66inter3));
  inv1  gate1223(.a(s_97), .O(gate66inter4));
  nand2 gate1224(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1225(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1226(.a(G26), .O(gate66inter7));
  inv1  gate1227(.a(G302), .O(gate66inter8));
  nand2 gate1228(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1229(.a(s_97), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1230(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1231(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1232(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1429(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1430(.a(gate70inter0), .b(s_126), .O(gate70inter1));
  and2  gate1431(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1432(.a(s_126), .O(gate70inter3));
  inv1  gate1433(.a(s_127), .O(gate70inter4));
  nand2 gate1434(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1435(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1436(.a(G30), .O(gate70inter7));
  inv1  gate1437(.a(G308), .O(gate70inter8));
  nand2 gate1438(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1439(.a(s_127), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1440(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1441(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1442(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1877(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1878(.a(gate74inter0), .b(s_190), .O(gate74inter1));
  and2  gate1879(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1880(.a(s_190), .O(gate74inter3));
  inv1  gate1881(.a(s_191), .O(gate74inter4));
  nand2 gate1882(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1883(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1884(.a(G5), .O(gate74inter7));
  inv1  gate1885(.a(G314), .O(gate74inter8));
  nand2 gate1886(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1887(.a(s_191), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1888(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1889(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1890(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1569(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1570(.a(gate75inter0), .b(s_146), .O(gate75inter1));
  and2  gate1571(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1572(.a(s_146), .O(gate75inter3));
  inv1  gate1573(.a(s_147), .O(gate75inter4));
  nand2 gate1574(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1575(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1576(.a(G9), .O(gate75inter7));
  inv1  gate1577(.a(G317), .O(gate75inter8));
  nand2 gate1578(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1579(.a(s_147), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1580(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1581(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1582(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1653(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1654(.a(gate86inter0), .b(s_158), .O(gate86inter1));
  and2  gate1655(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1656(.a(s_158), .O(gate86inter3));
  inv1  gate1657(.a(s_159), .O(gate86inter4));
  nand2 gate1658(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1659(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1660(.a(G8), .O(gate86inter7));
  inv1  gate1661(.a(G332), .O(gate86inter8));
  nand2 gate1662(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1663(.a(s_159), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1664(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1665(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1666(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1779(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1780(.a(gate87inter0), .b(s_176), .O(gate87inter1));
  and2  gate1781(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1782(.a(s_176), .O(gate87inter3));
  inv1  gate1783(.a(s_177), .O(gate87inter4));
  nand2 gate1784(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1785(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1786(.a(G12), .O(gate87inter7));
  inv1  gate1787(.a(G335), .O(gate87inter8));
  nand2 gate1788(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1789(.a(s_177), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1790(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1791(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1792(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1611(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1612(.a(gate89inter0), .b(s_152), .O(gate89inter1));
  and2  gate1613(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1614(.a(s_152), .O(gate89inter3));
  inv1  gate1615(.a(s_153), .O(gate89inter4));
  nand2 gate1616(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1617(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1618(.a(G17), .O(gate89inter7));
  inv1  gate1619(.a(G338), .O(gate89inter8));
  nand2 gate1620(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1621(.a(s_153), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1622(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1623(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1624(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate771(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate772(.a(gate92inter0), .b(s_32), .O(gate92inter1));
  and2  gate773(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate774(.a(s_32), .O(gate92inter3));
  inv1  gate775(.a(s_33), .O(gate92inter4));
  nand2 gate776(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate777(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate778(.a(G29), .O(gate92inter7));
  inv1  gate779(.a(G341), .O(gate92inter8));
  nand2 gate780(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate781(.a(s_33), .b(gate92inter3), .O(gate92inter10));
  nor2  gate782(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate783(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate784(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1135(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1136(.a(gate96inter0), .b(s_84), .O(gate96inter1));
  and2  gate1137(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1138(.a(s_84), .O(gate96inter3));
  inv1  gate1139(.a(s_85), .O(gate96inter4));
  nand2 gate1140(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1141(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1142(.a(G30), .O(gate96inter7));
  inv1  gate1143(.a(G347), .O(gate96inter8));
  nand2 gate1144(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1145(.a(s_85), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1146(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1147(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1148(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1863(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1864(.a(gate99inter0), .b(s_188), .O(gate99inter1));
  and2  gate1865(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1866(.a(s_188), .O(gate99inter3));
  inv1  gate1867(.a(s_189), .O(gate99inter4));
  nand2 gate1868(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1869(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1870(.a(G27), .O(gate99inter7));
  inv1  gate1871(.a(G353), .O(gate99inter8));
  nand2 gate1872(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1873(.a(s_189), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1874(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1875(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1876(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1023(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1024(.a(gate110inter0), .b(s_68), .O(gate110inter1));
  and2  gate1025(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1026(.a(s_68), .O(gate110inter3));
  inv1  gate1027(.a(s_69), .O(gate110inter4));
  nand2 gate1028(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1029(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1030(.a(G372), .O(gate110inter7));
  inv1  gate1031(.a(G373), .O(gate110inter8));
  nand2 gate1032(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1033(.a(s_69), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1034(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1035(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1036(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1009(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1010(.a(gate113inter0), .b(s_66), .O(gate113inter1));
  and2  gate1011(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1012(.a(s_66), .O(gate113inter3));
  inv1  gate1013(.a(s_67), .O(gate113inter4));
  nand2 gate1014(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1015(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1016(.a(G378), .O(gate113inter7));
  inv1  gate1017(.a(G379), .O(gate113inter8));
  nand2 gate1018(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1019(.a(s_67), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1020(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1021(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1022(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate687(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate688(.a(gate114inter0), .b(s_20), .O(gate114inter1));
  and2  gate689(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate690(.a(s_20), .O(gate114inter3));
  inv1  gate691(.a(s_21), .O(gate114inter4));
  nand2 gate692(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate693(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate694(.a(G380), .O(gate114inter7));
  inv1  gate695(.a(G381), .O(gate114inter8));
  nand2 gate696(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate697(.a(s_21), .b(gate114inter3), .O(gate114inter10));
  nor2  gate698(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate699(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate700(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate939(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate940(.a(gate117inter0), .b(s_56), .O(gate117inter1));
  and2  gate941(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate942(.a(s_56), .O(gate117inter3));
  inv1  gate943(.a(s_57), .O(gate117inter4));
  nand2 gate944(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate945(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate946(.a(G386), .O(gate117inter7));
  inv1  gate947(.a(G387), .O(gate117inter8));
  nand2 gate948(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate949(.a(s_57), .b(gate117inter3), .O(gate117inter10));
  nor2  gate950(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate951(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate952(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1443(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1444(.a(gate121inter0), .b(s_128), .O(gate121inter1));
  and2  gate1445(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1446(.a(s_128), .O(gate121inter3));
  inv1  gate1447(.a(s_129), .O(gate121inter4));
  nand2 gate1448(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1449(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1450(.a(G394), .O(gate121inter7));
  inv1  gate1451(.a(G395), .O(gate121inter8));
  nand2 gate1452(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1453(.a(s_129), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1454(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1455(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1456(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate715(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate716(.a(gate126inter0), .b(s_24), .O(gate126inter1));
  and2  gate717(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate718(.a(s_24), .O(gate126inter3));
  inv1  gate719(.a(s_25), .O(gate126inter4));
  nand2 gate720(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate721(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate722(.a(G404), .O(gate126inter7));
  inv1  gate723(.a(G405), .O(gate126inter8));
  nand2 gate724(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate725(.a(s_25), .b(gate126inter3), .O(gate126inter10));
  nor2  gate726(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate727(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate728(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1681(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1682(.a(gate132inter0), .b(s_162), .O(gate132inter1));
  and2  gate1683(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1684(.a(s_162), .O(gate132inter3));
  inv1  gate1685(.a(s_163), .O(gate132inter4));
  nand2 gate1686(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1687(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1688(.a(G416), .O(gate132inter7));
  inv1  gate1689(.a(G417), .O(gate132inter8));
  nand2 gate1690(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1691(.a(s_163), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1692(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1693(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1694(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1261(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1262(.a(gate135inter0), .b(s_102), .O(gate135inter1));
  and2  gate1263(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1264(.a(s_102), .O(gate135inter3));
  inv1  gate1265(.a(s_103), .O(gate135inter4));
  nand2 gate1266(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1267(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1268(.a(G422), .O(gate135inter7));
  inv1  gate1269(.a(G423), .O(gate135inter8));
  nand2 gate1270(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1271(.a(s_103), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1272(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1273(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1274(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate827(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate828(.a(gate144inter0), .b(s_40), .O(gate144inter1));
  and2  gate829(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate830(.a(s_40), .O(gate144inter3));
  inv1  gate831(.a(s_41), .O(gate144inter4));
  nand2 gate832(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate833(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate834(.a(G468), .O(gate144inter7));
  inv1  gate835(.a(G471), .O(gate144inter8));
  nand2 gate836(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate837(.a(s_41), .b(gate144inter3), .O(gate144inter10));
  nor2  gate838(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate839(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate840(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1583(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1584(.a(gate147inter0), .b(s_148), .O(gate147inter1));
  and2  gate1585(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1586(.a(s_148), .O(gate147inter3));
  inv1  gate1587(.a(s_149), .O(gate147inter4));
  nand2 gate1588(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1589(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1590(.a(G486), .O(gate147inter7));
  inv1  gate1591(.a(G489), .O(gate147inter8));
  nand2 gate1592(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1593(.a(s_149), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1594(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1595(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1596(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate757(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate758(.a(gate148inter0), .b(s_30), .O(gate148inter1));
  and2  gate759(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate760(.a(s_30), .O(gate148inter3));
  inv1  gate761(.a(s_31), .O(gate148inter4));
  nand2 gate762(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate763(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate764(.a(G492), .O(gate148inter7));
  inv1  gate765(.a(G495), .O(gate148inter8));
  nand2 gate766(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate767(.a(s_31), .b(gate148inter3), .O(gate148inter10));
  nor2  gate768(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate769(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate770(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate1639(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1640(.a(gate149inter0), .b(s_156), .O(gate149inter1));
  and2  gate1641(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1642(.a(s_156), .O(gate149inter3));
  inv1  gate1643(.a(s_157), .O(gate149inter4));
  nand2 gate1644(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1645(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1646(.a(G498), .O(gate149inter7));
  inv1  gate1647(.a(G501), .O(gate149inter8));
  nand2 gate1648(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1649(.a(s_157), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1650(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1651(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1652(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1317(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1318(.a(gate154inter0), .b(s_110), .O(gate154inter1));
  and2  gate1319(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1320(.a(s_110), .O(gate154inter3));
  inv1  gate1321(.a(s_111), .O(gate154inter4));
  nand2 gate1322(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1323(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1324(.a(G429), .O(gate154inter7));
  inv1  gate1325(.a(G522), .O(gate154inter8));
  nand2 gate1326(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1327(.a(s_111), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1328(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1329(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1330(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate659(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate660(.a(gate155inter0), .b(s_16), .O(gate155inter1));
  and2  gate661(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate662(.a(s_16), .O(gate155inter3));
  inv1  gate663(.a(s_17), .O(gate155inter4));
  nand2 gate664(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate665(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate666(.a(G432), .O(gate155inter7));
  inv1  gate667(.a(G525), .O(gate155inter8));
  nand2 gate668(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate669(.a(s_17), .b(gate155inter3), .O(gate155inter10));
  nor2  gate670(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate671(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate672(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate701(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate702(.a(gate157inter0), .b(s_22), .O(gate157inter1));
  and2  gate703(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate704(.a(s_22), .O(gate157inter3));
  inv1  gate705(.a(s_23), .O(gate157inter4));
  nand2 gate706(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate707(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate708(.a(G438), .O(gate157inter7));
  inv1  gate709(.a(G528), .O(gate157inter8));
  nand2 gate710(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate711(.a(s_23), .b(gate157inter3), .O(gate157inter10));
  nor2  gate712(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate713(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate714(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1667(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1668(.a(gate160inter0), .b(s_160), .O(gate160inter1));
  and2  gate1669(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1670(.a(s_160), .O(gate160inter3));
  inv1  gate1671(.a(s_161), .O(gate160inter4));
  nand2 gate1672(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1673(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1674(.a(G447), .O(gate160inter7));
  inv1  gate1675(.a(G531), .O(gate160inter8));
  nand2 gate1676(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1677(.a(s_161), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1678(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1679(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1680(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1037(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1038(.a(gate162inter0), .b(s_70), .O(gate162inter1));
  and2  gate1039(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1040(.a(s_70), .O(gate162inter3));
  inv1  gate1041(.a(s_71), .O(gate162inter4));
  nand2 gate1042(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1043(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1044(.a(G453), .O(gate162inter7));
  inv1  gate1045(.a(G534), .O(gate162inter8));
  nand2 gate1046(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1047(.a(s_71), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1048(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1049(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1050(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate645(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate646(.a(gate164inter0), .b(s_14), .O(gate164inter1));
  and2  gate647(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate648(.a(s_14), .O(gate164inter3));
  inv1  gate649(.a(s_15), .O(gate164inter4));
  nand2 gate650(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate651(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate652(.a(G459), .O(gate164inter7));
  inv1  gate653(.a(G537), .O(gate164inter8));
  nand2 gate654(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate655(.a(s_15), .b(gate164inter3), .O(gate164inter10));
  nor2  gate656(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate657(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate658(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate841(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate842(.a(gate165inter0), .b(s_42), .O(gate165inter1));
  and2  gate843(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate844(.a(s_42), .O(gate165inter3));
  inv1  gate845(.a(s_43), .O(gate165inter4));
  nand2 gate846(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate847(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate848(.a(G462), .O(gate165inter7));
  inv1  gate849(.a(G540), .O(gate165inter8));
  nand2 gate850(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate851(.a(s_43), .b(gate165inter3), .O(gate165inter10));
  nor2  gate852(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate853(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate854(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1359(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1360(.a(gate171inter0), .b(s_116), .O(gate171inter1));
  and2  gate1361(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1362(.a(s_116), .O(gate171inter3));
  inv1  gate1363(.a(s_117), .O(gate171inter4));
  nand2 gate1364(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1365(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1366(.a(G480), .O(gate171inter7));
  inv1  gate1367(.a(G549), .O(gate171inter8));
  nand2 gate1368(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1369(.a(s_117), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1370(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1371(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1372(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1233(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1234(.a(gate172inter0), .b(s_98), .O(gate172inter1));
  and2  gate1235(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1236(.a(s_98), .O(gate172inter3));
  inv1  gate1237(.a(s_99), .O(gate172inter4));
  nand2 gate1238(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1239(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1240(.a(G483), .O(gate172inter7));
  inv1  gate1241(.a(G549), .O(gate172inter8));
  nand2 gate1242(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1243(.a(s_99), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1244(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1245(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1246(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1527(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1528(.a(gate184inter0), .b(s_140), .O(gate184inter1));
  and2  gate1529(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1530(.a(s_140), .O(gate184inter3));
  inv1  gate1531(.a(s_141), .O(gate184inter4));
  nand2 gate1532(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1533(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1534(.a(G519), .O(gate184inter7));
  inv1  gate1535(.a(G567), .O(gate184inter8));
  nand2 gate1536(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1537(.a(s_141), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1538(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1539(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1540(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate995(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate996(.a(gate222inter0), .b(s_64), .O(gate222inter1));
  and2  gate997(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate998(.a(s_64), .O(gate222inter3));
  inv1  gate999(.a(s_65), .O(gate222inter4));
  nand2 gate1000(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1001(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1002(.a(G632), .O(gate222inter7));
  inv1  gate1003(.a(G684), .O(gate222inter8));
  nand2 gate1004(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1005(.a(s_65), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1006(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1007(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1008(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1275(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1276(.a(gate225inter0), .b(s_104), .O(gate225inter1));
  and2  gate1277(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1278(.a(s_104), .O(gate225inter3));
  inv1  gate1279(.a(s_105), .O(gate225inter4));
  nand2 gate1280(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1281(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1282(.a(G690), .O(gate225inter7));
  inv1  gate1283(.a(G691), .O(gate225inter8));
  nand2 gate1284(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1285(.a(s_105), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1286(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1287(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1288(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate603(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate604(.a(gate227inter0), .b(s_8), .O(gate227inter1));
  and2  gate605(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate606(.a(s_8), .O(gate227inter3));
  inv1  gate607(.a(s_9), .O(gate227inter4));
  nand2 gate608(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate609(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate610(.a(G694), .O(gate227inter7));
  inv1  gate611(.a(G695), .O(gate227inter8));
  nand2 gate612(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate613(.a(s_9), .b(gate227inter3), .O(gate227inter10));
  nor2  gate614(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate615(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate616(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate561(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate562(.a(gate233inter0), .b(s_2), .O(gate233inter1));
  and2  gate563(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate564(.a(s_2), .O(gate233inter3));
  inv1  gate565(.a(s_3), .O(gate233inter4));
  nand2 gate566(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate567(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate568(.a(G242), .O(gate233inter7));
  inv1  gate569(.a(G718), .O(gate233inter8));
  nand2 gate570(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate571(.a(s_3), .b(gate233inter3), .O(gate233inter10));
  nor2  gate572(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate573(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate574(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1387(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1388(.a(gate236inter0), .b(s_120), .O(gate236inter1));
  and2  gate1389(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1390(.a(s_120), .O(gate236inter3));
  inv1  gate1391(.a(s_121), .O(gate236inter4));
  nand2 gate1392(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1393(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1394(.a(G251), .O(gate236inter7));
  inv1  gate1395(.a(G727), .O(gate236inter8));
  nand2 gate1396(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1397(.a(s_121), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1398(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1399(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1400(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1051(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1052(.a(gate239inter0), .b(s_72), .O(gate239inter1));
  and2  gate1053(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1054(.a(s_72), .O(gate239inter3));
  inv1  gate1055(.a(s_73), .O(gate239inter4));
  nand2 gate1056(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1057(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1058(.a(G260), .O(gate239inter7));
  inv1  gate1059(.a(G712), .O(gate239inter8));
  nand2 gate1060(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1061(.a(s_73), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1062(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1063(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1064(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate911(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate912(.a(gate241inter0), .b(s_52), .O(gate241inter1));
  and2  gate913(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate914(.a(s_52), .O(gate241inter3));
  inv1  gate915(.a(s_53), .O(gate241inter4));
  nand2 gate916(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate917(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate918(.a(G242), .O(gate241inter7));
  inv1  gate919(.a(G730), .O(gate241inter8));
  nand2 gate920(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate921(.a(s_53), .b(gate241inter3), .O(gate241inter10));
  nor2  gate922(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate923(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate924(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1485(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1486(.a(gate242inter0), .b(s_134), .O(gate242inter1));
  and2  gate1487(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1488(.a(s_134), .O(gate242inter3));
  inv1  gate1489(.a(s_135), .O(gate242inter4));
  nand2 gate1490(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1491(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1492(.a(G718), .O(gate242inter7));
  inv1  gate1493(.a(G730), .O(gate242inter8));
  nand2 gate1494(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1495(.a(s_135), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1496(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1497(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1498(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate869(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate870(.a(gate250inter0), .b(s_46), .O(gate250inter1));
  and2  gate871(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate872(.a(s_46), .O(gate250inter3));
  inv1  gate873(.a(s_47), .O(gate250inter4));
  nand2 gate874(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate875(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate876(.a(G706), .O(gate250inter7));
  inv1  gate877(.a(G742), .O(gate250inter8));
  nand2 gate878(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate879(.a(s_47), .b(gate250inter3), .O(gate250inter10));
  nor2  gate880(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate881(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate882(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1737(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1738(.a(gate251inter0), .b(s_170), .O(gate251inter1));
  and2  gate1739(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1740(.a(s_170), .O(gate251inter3));
  inv1  gate1741(.a(s_171), .O(gate251inter4));
  nand2 gate1742(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1743(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1744(.a(G257), .O(gate251inter7));
  inv1  gate1745(.a(G745), .O(gate251inter8));
  nand2 gate1746(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1747(.a(s_171), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1748(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1749(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1750(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1401(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1402(.a(gate254inter0), .b(s_122), .O(gate254inter1));
  and2  gate1403(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1404(.a(s_122), .O(gate254inter3));
  inv1  gate1405(.a(s_123), .O(gate254inter4));
  nand2 gate1406(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1407(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1408(.a(G712), .O(gate254inter7));
  inv1  gate1409(.a(G748), .O(gate254inter8));
  nand2 gate1410(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1411(.a(s_123), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1412(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1413(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1414(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1331(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1332(.a(gate256inter0), .b(s_112), .O(gate256inter1));
  and2  gate1333(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1334(.a(s_112), .O(gate256inter3));
  inv1  gate1335(.a(s_113), .O(gate256inter4));
  nand2 gate1336(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1337(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1338(.a(G715), .O(gate256inter7));
  inv1  gate1339(.a(G751), .O(gate256inter8));
  nand2 gate1340(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1341(.a(s_113), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1342(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1343(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1344(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate953(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate954(.a(gate262inter0), .b(s_58), .O(gate262inter1));
  and2  gate955(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate956(.a(s_58), .O(gate262inter3));
  inv1  gate957(.a(s_59), .O(gate262inter4));
  nand2 gate958(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate959(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate960(.a(G764), .O(gate262inter7));
  inv1  gate961(.a(G765), .O(gate262inter8));
  nand2 gate962(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate963(.a(s_59), .b(gate262inter3), .O(gate262inter10));
  nor2  gate964(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate965(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate966(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate617(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate618(.a(gate266inter0), .b(s_10), .O(gate266inter1));
  and2  gate619(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate620(.a(s_10), .O(gate266inter3));
  inv1  gate621(.a(s_11), .O(gate266inter4));
  nand2 gate622(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate623(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate624(.a(G645), .O(gate266inter7));
  inv1  gate625(.a(G773), .O(gate266inter8));
  nand2 gate626(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate627(.a(s_11), .b(gate266inter3), .O(gate266inter10));
  nor2  gate628(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate629(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate630(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1555(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1556(.a(gate268inter0), .b(s_144), .O(gate268inter1));
  and2  gate1557(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1558(.a(s_144), .O(gate268inter3));
  inv1  gate1559(.a(s_145), .O(gate268inter4));
  nand2 gate1560(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1561(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1562(.a(G651), .O(gate268inter7));
  inv1  gate1563(.a(G779), .O(gate268inter8));
  nand2 gate1564(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1565(.a(s_145), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1566(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1567(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1568(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1121(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1122(.a(gate269inter0), .b(s_82), .O(gate269inter1));
  and2  gate1123(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1124(.a(s_82), .O(gate269inter3));
  inv1  gate1125(.a(s_83), .O(gate269inter4));
  nand2 gate1126(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1127(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1128(.a(G654), .O(gate269inter7));
  inv1  gate1129(.a(G782), .O(gate269inter8));
  nand2 gate1130(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1131(.a(s_83), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1132(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1133(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1134(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate883(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate884(.a(gate275inter0), .b(s_48), .O(gate275inter1));
  and2  gate885(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate886(.a(s_48), .O(gate275inter3));
  inv1  gate887(.a(s_49), .O(gate275inter4));
  nand2 gate888(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate889(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate890(.a(G645), .O(gate275inter7));
  inv1  gate891(.a(G797), .O(gate275inter8));
  nand2 gate892(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate893(.a(s_49), .b(gate275inter3), .O(gate275inter10));
  nor2  gate894(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate895(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate896(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1723(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1724(.a(gate277inter0), .b(s_168), .O(gate277inter1));
  and2  gate1725(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1726(.a(s_168), .O(gate277inter3));
  inv1  gate1727(.a(s_169), .O(gate277inter4));
  nand2 gate1728(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1729(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1730(.a(G648), .O(gate277inter7));
  inv1  gate1731(.a(G800), .O(gate277inter8));
  nand2 gate1732(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1733(.a(s_169), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1734(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1735(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1736(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate743(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate744(.a(gate279inter0), .b(s_28), .O(gate279inter1));
  and2  gate745(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate746(.a(s_28), .O(gate279inter3));
  inv1  gate747(.a(s_29), .O(gate279inter4));
  nand2 gate748(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate749(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate750(.a(G651), .O(gate279inter7));
  inv1  gate751(.a(G803), .O(gate279inter8));
  nand2 gate752(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate753(.a(s_29), .b(gate279inter3), .O(gate279inter10));
  nor2  gate754(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate755(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate756(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate799(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate800(.a(gate282inter0), .b(s_36), .O(gate282inter1));
  and2  gate801(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate802(.a(s_36), .O(gate282inter3));
  inv1  gate803(.a(s_37), .O(gate282inter4));
  nand2 gate804(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate805(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate806(.a(G782), .O(gate282inter7));
  inv1  gate807(.a(G806), .O(gate282inter8));
  nand2 gate808(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate809(.a(s_37), .b(gate282inter3), .O(gate282inter10));
  nor2  gate810(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate811(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate812(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1807(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1808(.a(gate285inter0), .b(s_180), .O(gate285inter1));
  and2  gate1809(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1810(.a(s_180), .O(gate285inter3));
  inv1  gate1811(.a(s_181), .O(gate285inter4));
  nand2 gate1812(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1813(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1814(.a(G660), .O(gate285inter7));
  inv1  gate1815(.a(G812), .O(gate285inter8));
  nand2 gate1816(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1817(.a(s_181), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1818(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1819(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1820(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate785(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate786(.a(gate287inter0), .b(s_34), .O(gate287inter1));
  and2  gate787(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate788(.a(s_34), .O(gate287inter3));
  inv1  gate789(.a(s_35), .O(gate287inter4));
  nand2 gate790(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate791(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate792(.a(G663), .O(gate287inter7));
  inv1  gate793(.a(G815), .O(gate287inter8));
  nand2 gate794(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate795(.a(s_35), .b(gate287inter3), .O(gate287inter10));
  nor2  gate796(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate797(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate798(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1303(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1304(.a(gate387inter0), .b(s_108), .O(gate387inter1));
  and2  gate1305(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1306(.a(s_108), .O(gate387inter3));
  inv1  gate1307(.a(s_109), .O(gate387inter4));
  nand2 gate1308(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1309(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1310(.a(G1), .O(gate387inter7));
  inv1  gate1311(.a(G1036), .O(gate387inter8));
  nand2 gate1312(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1313(.a(s_109), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1314(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1315(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1316(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1149(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1150(.a(gate394inter0), .b(s_86), .O(gate394inter1));
  and2  gate1151(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1152(.a(s_86), .O(gate394inter3));
  inv1  gate1153(.a(s_87), .O(gate394inter4));
  nand2 gate1154(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1155(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1156(.a(G8), .O(gate394inter7));
  inv1  gate1157(.a(G1057), .O(gate394inter8));
  nand2 gate1158(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1159(.a(s_87), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1160(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1161(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1162(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate813(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate814(.a(gate396inter0), .b(s_38), .O(gate396inter1));
  and2  gate815(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate816(.a(s_38), .O(gate396inter3));
  inv1  gate817(.a(s_39), .O(gate396inter4));
  nand2 gate818(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate819(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate820(.a(G10), .O(gate396inter7));
  inv1  gate821(.a(G1063), .O(gate396inter8));
  nand2 gate822(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate823(.a(s_39), .b(gate396inter3), .O(gate396inter10));
  nor2  gate824(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate825(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate826(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1765(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1766(.a(gate399inter0), .b(s_174), .O(gate399inter1));
  and2  gate1767(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1768(.a(s_174), .O(gate399inter3));
  inv1  gate1769(.a(s_175), .O(gate399inter4));
  nand2 gate1770(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1771(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1772(.a(G13), .O(gate399inter7));
  inv1  gate1773(.a(G1072), .O(gate399inter8));
  nand2 gate1774(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1775(.a(s_175), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1776(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1777(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1778(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate547(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate548(.a(gate402inter0), .b(s_0), .O(gate402inter1));
  and2  gate549(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate550(.a(s_0), .O(gate402inter3));
  inv1  gate551(.a(s_1), .O(gate402inter4));
  nand2 gate552(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate553(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate554(.a(G16), .O(gate402inter7));
  inv1  gate555(.a(G1081), .O(gate402inter8));
  nand2 gate556(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate557(.a(s_1), .b(gate402inter3), .O(gate402inter10));
  nor2  gate558(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate559(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate560(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate967(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate968(.a(gate404inter0), .b(s_60), .O(gate404inter1));
  and2  gate969(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate970(.a(s_60), .O(gate404inter3));
  inv1  gate971(.a(s_61), .O(gate404inter4));
  nand2 gate972(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate973(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate974(.a(G18), .O(gate404inter7));
  inv1  gate975(.a(G1087), .O(gate404inter8));
  nand2 gate976(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate977(.a(s_61), .b(gate404inter3), .O(gate404inter10));
  nor2  gate978(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate979(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate980(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1849(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1850(.a(gate411inter0), .b(s_186), .O(gate411inter1));
  and2  gate1851(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1852(.a(s_186), .O(gate411inter3));
  inv1  gate1853(.a(s_187), .O(gate411inter4));
  nand2 gate1854(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1855(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1856(.a(G25), .O(gate411inter7));
  inv1  gate1857(.a(G1108), .O(gate411inter8));
  nand2 gate1858(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1859(.a(s_187), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1860(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1861(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1862(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1065(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1066(.a(gate422inter0), .b(s_74), .O(gate422inter1));
  and2  gate1067(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1068(.a(s_74), .O(gate422inter3));
  inv1  gate1069(.a(s_75), .O(gate422inter4));
  nand2 gate1070(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1071(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1072(.a(G1039), .O(gate422inter7));
  inv1  gate1073(.a(G1135), .O(gate422inter8));
  nand2 gate1074(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1075(.a(s_75), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1076(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1077(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1078(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1205(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1206(.a(gate425inter0), .b(s_94), .O(gate425inter1));
  and2  gate1207(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1208(.a(s_94), .O(gate425inter3));
  inv1  gate1209(.a(s_95), .O(gate425inter4));
  nand2 gate1210(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1211(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1212(.a(G4), .O(gate425inter7));
  inv1  gate1213(.a(G1141), .O(gate425inter8));
  nand2 gate1214(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1215(.a(s_95), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1216(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1217(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1218(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1835(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1836(.a(gate426inter0), .b(s_184), .O(gate426inter1));
  and2  gate1837(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1838(.a(s_184), .O(gate426inter3));
  inv1  gate1839(.a(s_185), .O(gate426inter4));
  nand2 gate1840(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1841(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1842(.a(G1045), .O(gate426inter7));
  inv1  gate1843(.a(G1141), .O(gate426inter8));
  nand2 gate1844(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1845(.a(s_185), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1846(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1847(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1848(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate673(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate674(.a(gate436inter0), .b(s_18), .O(gate436inter1));
  and2  gate675(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate676(.a(s_18), .O(gate436inter3));
  inv1  gate677(.a(s_19), .O(gate436inter4));
  nand2 gate678(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate679(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate680(.a(G1060), .O(gate436inter7));
  inv1  gate681(.a(G1156), .O(gate436inter8));
  nand2 gate682(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate683(.a(s_19), .b(gate436inter3), .O(gate436inter10));
  nor2  gate684(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate685(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate686(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1457(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1458(.a(gate439inter0), .b(s_130), .O(gate439inter1));
  and2  gate1459(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1460(.a(s_130), .O(gate439inter3));
  inv1  gate1461(.a(s_131), .O(gate439inter4));
  nand2 gate1462(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1463(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1464(.a(G11), .O(gate439inter7));
  inv1  gate1465(.a(G1162), .O(gate439inter8));
  nand2 gate1466(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1467(.a(s_131), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1468(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1469(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1470(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1709(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1710(.a(gate440inter0), .b(s_166), .O(gate440inter1));
  and2  gate1711(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1712(.a(s_166), .O(gate440inter3));
  inv1  gate1713(.a(s_167), .O(gate440inter4));
  nand2 gate1714(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1715(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1716(.a(G1066), .O(gate440inter7));
  inv1  gate1717(.a(G1162), .O(gate440inter8));
  nand2 gate1718(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1719(.a(s_167), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1720(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1721(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1722(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1821(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1822(.a(gate441inter0), .b(s_182), .O(gate441inter1));
  and2  gate1823(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1824(.a(s_182), .O(gate441inter3));
  inv1  gate1825(.a(s_183), .O(gate441inter4));
  nand2 gate1826(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1827(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1828(.a(G12), .O(gate441inter7));
  inv1  gate1829(.a(G1165), .O(gate441inter8));
  nand2 gate1830(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1831(.a(s_183), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1832(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1833(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1834(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate589(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate590(.a(gate446inter0), .b(s_6), .O(gate446inter1));
  and2  gate591(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate592(.a(s_6), .O(gate446inter3));
  inv1  gate593(.a(s_7), .O(gate446inter4));
  nand2 gate594(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate595(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate596(.a(G1075), .O(gate446inter7));
  inv1  gate597(.a(G1171), .O(gate446inter8));
  nand2 gate598(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate599(.a(s_7), .b(gate446inter3), .O(gate446inter10));
  nor2  gate600(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate601(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate602(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1093(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1094(.a(gate454inter0), .b(s_78), .O(gate454inter1));
  and2  gate1095(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1096(.a(s_78), .O(gate454inter3));
  inv1  gate1097(.a(s_79), .O(gate454inter4));
  nand2 gate1098(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1099(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1100(.a(G1087), .O(gate454inter7));
  inv1  gate1101(.a(G1183), .O(gate454inter8));
  nand2 gate1102(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1103(.a(s_79), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1104(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1105(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1106(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate575(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate576(.a(gate456inter0), .b(s_4), .O(gate456inter1));
  and2  gate577(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate578(.a(s_4), .O(gate456inter3));
  inv1  gate579(.a(s_5), .O(gate456inter4));
  nand2 gate580(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate581(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate582(.a(G1090), .O(gate456inter7));
  inv1  gate583(.a(G1186), .O(gate456inter8));
  nand2 gate584(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate585(.a(s_5), .b(gate456inter3), .O(gate456inter10));
  nor2  gate586(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate587(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate588(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1345(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1346(.a(gate459inter0), .b(s_114), .O(gate459inter1));
  and2  gate1347(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1348(.a(s_114), .O(gate459inter3));
  inv1  gate1349(.a(s_115), .O(gate459inter4));
  nand2 gate1350(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1351(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1352(.a(G21), .O(gate459inter7));
  inv1  gate1353(.a(G1192), .O(gate459inter8));
  nand2 gate1354(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1355(.a(s_115), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1356(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1357(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1358(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1499(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1500(.a(gate462inter0), .b(s_136), .O(gate462inter1));
  and2  gate1501(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1502(.a(s_136), .O(gate462inter3));
  inv1  gate1503(.a(s_137), .O(gate462inter4));
  nand2 gate1504(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1505(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1506(.a(G1099), .O(gate462inter7));
  inv1  gate1507(.a(G1195), .O(gate462inter8));
  nand2 gate1508(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1509(.a(s_137), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1510(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1511(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1512(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate729(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate730(.a(gate464inter0), .b(s_26), .O(gate464inter1));
  and2  gate731(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate732(.a(s_26), .O(gate464inter3));
  inv1  gate733(.a(s_27), .O(gate464inter4));
  nand2 gate734(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate735(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate736(.a(G1102), .O(gate464inter7));
  inv1  gate737(.a(G1198), .O(gate464inter8));
  nand2 gate738(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate739(.a(s_27), .b(gate464inter3), .O(gate464inter10));
  nor2  gate740(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate741(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate742(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate855(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate856(.a(gate465inter0), .b(s_44), .O(gate465inter1));
  and2  gate857(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate858(.a(s_44), .O(gate465inter3));
  inv1  gate859(.a(s_45), .O(gate465inter4));
  nand2 gate860(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate861(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate862(.a(G24), .O(gate465inter7));
  inv1  gate863(.a(G1201), .O(gate465inter8));
  nand2 gate864(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate865(.a(s_45), .b(gate465inter3), .O(gate465inter10));
  nor2  gate866(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate867(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate868(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1373(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1374(.a(gate466inter0), .b(s_118), .O(gate466inter1));
  and2  gate1375(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1376(.a(s_118), .O(gate466inter3));
  inv1  gate1377(.a(s_119), .O(gate466inter4));
  nand2 gate1378(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1379(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1380(.a(G1105), .O(gate466inter7));
  inv1  gate1381(.a(G1201), .O(gate466inter8));
  nand2 gate1382(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1383(.a(s_119), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1384(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1385(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1386(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate925(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate926(.a(gate470inter0), .b(s_54), .O(gate470inter1));
  and2  gate927(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate928(.a(s_54), .O(gate470inter3));
  inv1  gate929(.a(s_55), .O(gate470inter4));
  nand2 gate930(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate931(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate932(.a(G1111), .O(gate470inter7));
  inv1  gate933(.a(G1207), .O(gate470inter8));
  nand2 gate934(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate935(.a(s_55), .b(gate470inter3), .O(gate470inter10));
  nor2  gate936(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate937(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate938(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1751(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1752(.a(gate473inter0), .b(s_172), .O(gate473inter1));
  and2  gate1753(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1754(.a(s_172), .O(gate473inter3));
  inv1  gate1755(.a(s_173), .O(gate473inter4));
  nand2 gate1756(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1757(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1758(.a(G28), .O(gate473inter7));
  inv1  gate1759(.a(G1213), .O(gate473inter8));
  nand2 gate1760(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1761(.a(s_173), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1762(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1763(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1764(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1191(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1192(.a(gate479inter0), .b(s_92), .O(gate479inter1));
  and2  gate1193(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1194(.a(s_92), .O(gate479inter3));
  inv1  gate1195(.a(s_93), .O(gate479inter4));
  nand2 gate1196(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1197(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1198(.a(G31), .O(gate479inter7));
  inv1  gate1199(.a(G1222), .O(gate479inter8));
  nand2 gate1200(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1201(.a(s_93), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1202(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1203(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1204(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1415(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1416(.a(gate497inter0), .b(s_124), .O(gate497inter1));
  and2  gate1417(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1418(.a(s_124), .O(gate497inter3));
  inv1  gate1419(.a(s_125), .O(gate497inter4));
  nand2 gate1420(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1421(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1422(.a(G1256), .O(gate497inter7));
  inv1  gate1423(.a(G1257), .O(gate497inter8));
  nand2 gate1424(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1425(.a(s_125), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1426(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1427(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1428(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate897(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate898(.a(gate507inter0), .b(s_50), .O(gate507inter1));
  and2  gate899(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate900(.a(s_50), .O(gate507inter3));
  inv1  gate901(.a(s_51), .O(gate507inter4));
  nand2 gate902(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate903(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate904(.a(G1276), .O(gate507inter7));
  inv1  gate905(.a(G1277), .O(gate507inter8));
  nand2 gate906(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate907(.a(s_51), .b(gate507inter3), .O(gate507inter10));
  nor2  gate908(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate909(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate910(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1793(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1794(.a(gate508inter0), .b(s_178), .O(gate508inter1));
  and2  gate1795(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1796(.a(s_178), .O(gate508inter3));
  inv1  gate1797(.a(s_179), .O(gate508inter4));
  nand2 gate1798(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1799(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1800(.a(G1278), .O(gate508inter7));
  inv1  gate1801(.a(G1279), .O(gate508inter8));
  nand2 gate1802(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1803(.a(s_179), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1804(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1805(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1806(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1695(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1696(.a(gate509inter0), .b(s_164), .O(gate509inter1));
  and2  gate1697(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1698(.a(s_164), .O(gate509inter3));
  inv1  gate1699(.a(s_165), .O(gate509inter4));
  nand2 gate1700(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1701(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1702(.a(G1280), .O(gate509inter7));
  inv1  gate1703(.a(G1281), .O(gate509inter8));
  nand2 gate1704(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1705(.a(s_165), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1706(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1707(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1708(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1079(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1080(.a(gate514inter0), .b(s_76), .O(gate514inter1));
  and2  gate1081(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1082(.a(s_76), .O(gate514inter3));
  inv1  gate1083(.a(s_77), .O(gate514inter4));
  nand2 gate1084(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1085(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1086(.a(G1290), .O(gate514inter7));
  inv1  gate1087(.a(G1291), .O(gate514inter8));
  nand2 gate1088(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1089(.a(s_77), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1090(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1091(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1092(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule