module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );

  xor2  gate175(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate176(.a(gate20inter0), .b(s_2), .O(gate20inter1));
  and2  gate177(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate178(.a(s_2), .O(gate20inter3));
  inv1  gate179(.a(s_3), .O(gate20inter4));
  nand2 gate180(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate181(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate182(.a(N8), .O(gate20inter7));
  inv1  gate183(.a(N119), .O(gate20inter8));
  nand2 gate184(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate185(.a(s_3), .b(gate20inter3), .O(gate20inter10));
  nor2  gate186(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate187(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate188(.a(gate20inter12), .b(gate20inter1), .O(N157));

  xor2  gate483(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate484(.a(gate21inter0), .b(s_46), .O(gate21inter1));
  and2  gate485(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate486(.a(s_46), .O(gate21inter3));
  inv1  gate487(.a(s_47), .O(gate21inter4));
  nand2 gate488(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate489(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate490(.a(N14), .O(gate21inter7));
  inv1  gate491(.a(N119), .O(gate21inter8));
  nand2 gate492(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate493(.a(s_47), .b(gate21inter3), .O(gate21inter10));
  nor2  gate494(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate495(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate496(.a(gate21inter12), .b(gate21inter1), .O(N158));
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate161(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate162(.a(gate29inter0), .b(s_0), .O(gate29inter1));
  and2  gate163(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate164(.a(s_0), .O(gate29inter3));
  inv1  gate165(.a(s_1), .O(gate29inter4));
  nand2 gate166(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate167(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate168(.a(N150), .O(gate29inter7));
  inv1  gate169(.a(N108), .O(gate29inter8));
  nand2 gate170(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate171(.a(s_1), .b(gate29inter3), .O(gate29inter10));
  nor2  gate172(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate173(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate174(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );

  xor2  gate441(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate442(.a(gate31inter0), .b(s_40), .O(gate31inter1));
  and2  gate443(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate444(.a(s_40), .O(gate31inter3));
  inv1  gate445(.a(s_41), .O(gate31inter4));
  nand2 gate446(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate447(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate448(.a(N27), .O(gate31inter7));
  inv1  gate449(.a(N123), .O(gate31inter8));
  nand2 gate450(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate451(.a(s_41), .b(gate31inter3), .O(gate31inter10));
  nor2  gate452(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate453(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate454(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );

  xor2  gate511(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate512(.a(gate39inter0), .b(s_50), .O(gate39inter1));
  and2  gate513(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate514(.a(s_50), .O(gate39inter3));
  inv1  gate515(.a(s_51), .O(gate39inter4));
  nand2 gate516(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate517(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate518(.a(N79), .O(gate39inter7));
  inv1  gate519(.a(N139), .O(gate39inter8));
  nand2 gate520(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate521(.a(s_51), .b(gate39inter3), .O(gate39inter10));
  nor2  gate522(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate523(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate524(.a(gate39inter12), .b(gate39inter1), .O(N192));

  xor2  gate287(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate288(.a(gate40inter0), .b(s_18), .O(gate40inter1));
  and2  gate289(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate290(.a(s_18), .O(gate40inter3));
  inv1  gate291(.a(s_19), .O(gate40inter4));
  nand2 gate292(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate293(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate294(.a(N86), .O(gate40inter7));
  inv1  gate295(.a(N143), .O(gate40inter8));
  nand2 gate296(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate297(.a(s_19), .b(gate40inter3), .O(gate40inter10));
  nor2  gate298(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate299(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate300(.a(gate40inter12), .b(gate40inter1), .O(N193));
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );

  xor2  gate413(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate414(.a(gate58inter0), .b(s_36), .O(gate58inter1));
  and2  gate415(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate416(.a(s_36), .O(gate58inter3));
  inv1  gate417(.a(s_37), .O(gate58inter4));
  nand2 gate418(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate419(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate420(.a(N213), .O(gate58inter7));
  inv1  gate421(.a(N11), .O(gate58inter8));
  nand2 gate422(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate423(.a(s_37), .b(gate58inter3), .O(gate58inter10));
  nor2  gate424(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate425(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate426(.a(gate58inter12), .b(gate58inter1), .O(N246));

  xor2  gate399(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate400(.a(gate59inter0), .b(s_34), .O(gate59inter1));
  and2  gate401(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate402(.a(s_34), .O(gate59inter3));
  inv1  gate403(.a(s_35), .O(gate59inter4));
  nand2 gate404(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate405(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate406(.a(N203), .O(gate59inter7));
  inv1  gate407(.a(N177), .O(gate59inter8));
  nand2 gate408(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate409(.a(s_35), .b(gate59inter3), .O(gate59inter10));
  nor2  gate410(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate411(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate412(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate371(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate372(.a(gate70inter0), .b(s_30), .O(gate70inter1));
  and2  gate373(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate374(.a(s_30), .O(gate70inter3));
  inv1  gate375(.a(s_31), .O(gate70inter4));
  nand2 gate376(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate377(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate378(.a(N227), .O(gate70inter7));
  inv1  gate379(.a(N183), .O(gate70inter8));
  nand2 gate380(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate381(.a(s_31), .b(gate70inter3), .O(gate70inter10));
  nor2  gate382(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate383(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate384(.a(gate70inter12), .b(gate70inter1), .O(N264));

  xor2  gate329(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate330(.a(gate71inter0), .b(s_24), .O(gate71inter1));
  and2  gate331(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate332(.a(s_24), .O(gate71inter3));
  inv1  gate333(.a(s_25), .O(gate71inter4));
  nand2 gate334(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate335(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate336(.a(N230), .O(gate71inter7));
  inv1  gate337(.a(N185), .O(gate71inter8));
  nand2 gate338(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate339(.a(s_25), .b(gate71inter3), .O(gate71inter10));
  nor2  gate340(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate341(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate342(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate357(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate358(.a(gate73inter0), .b(s_28), .O(gate73inter1));
  and2  gate359(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate360(.a(s_28), .O(gate73inter3));
  inv1  gate361(.a(s_29), .O(gate73inter4));
  nand2 gate362(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate363(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate364(.a(N236), .O(gate73inter7));
  inv1  gate365(.a(N189), .O(gate73inter8));
  nand2 gate366(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate367(.a(s_29), .b(gate73inter3), .O(gate73inter10));
  nor2  gate368(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate369(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate370(.a(gate73inter12), .b(gate73inter1), .O(N273));

  xor2  gate385(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate386(.a(gate74inter0), .b(s_32), .O(gate74inter1));
  and2  gate387(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate388(.a(s_32), .O(gate74inter3));
  inv1  gate389(.a(s_33), .O(gate74inter4));
  nand2 gate390(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate391(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate392(.a(N239), .O(gate74inter7));
  inv1  gate393(.a(N191), .O(gate74inter8));
  nand2 gate394(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate395(.a(s_33), .b(gate74inter3), .O(gate74inter10));
  nor2  gate396(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate397(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate398(.a(gate74inter12), .b(gate74inter1), .O(N276));
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate273(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate274(.a(gate78inter0), .b(s_16), .O(gate78inter1));
  and2  gate275(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate276(.a(s_16), .O(gate78inter3));
  inv1  gate277(.a(s_17), .O(gate78inter4));
  nand2 gate278(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate279(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate280(.a(N227), .O(gate78inter7));
  inv1  gate281(.a(N184), .O(gate78inter8));
  nand2 gate282(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate283(.a(s_17), .b(gate78inter3), .O(gate78inter10));
  nor2  gate284(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate285(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate286(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );

  xor2  gate203(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate204(.a(gate81inter0), .b(s_6), .O(gate81inter1));
  and2  gate205(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate206(.a(s_6), .O(gate81inter3));
  inv1  gate207(.a(s_7), .O(gate81inter4));
  nand2 gate208(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate209(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate210(.a(N236), .O(gate81inter7));
  inv1  gate211(.a(N190), .O(gate81inter8));
  nand2 gate212(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate213(.a(s_7), .b(gate81inter3), .O(gate81inter10));
  nor2  gate214(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate215(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate216(.a(gate81inter12), .b(gate81inter1), .O(N291));
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );

  xor2  gate343(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate344(.a(gate85inter0), .b(s_26), .O(gate85inter1));
  and2  gate345(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate346(.a(s_26), .O(gate85inter3));
  inv1  gate347(.a(s_27), .O(gate85inter4));
  nand2 gate348(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate349(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate350(.a(N251), .O(gate85inter7));
  inv1  gate351(.a(N198), .O(gate85inter8));
  nand2 gate352(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate353(.a(s_27), .b(gate85inter3), .O(gate85inter10));
  nor2  gate354(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate355(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate356(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate245(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate246(.a(gate99inter0), .b(s_12), .O(gate99inter1));
  and2  gate247(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate248(.a(s_12), .O(gate99inter3));
  inv1  gate249(.a(s_13), .O(gate99inter4));
  nand2 gate250(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate251(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate252(.a(N309), .O(gate99inter7));
  inv1  gate253(.a(N260), .O(gate99inter8));
  nand2 gate254(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate255(.a(s_13), .b(gate99inter3), .O(gate99inter10));
  nor2  gate256(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate257(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate258(.a(gate99inter12), .b(gate99inter1), .O(N330));
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );

  xor2  gate189(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate190(.a(gate106inter0), .b(s_4), .O(gate106inter1));
  and2  gate191(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate192(.a(s_4), .O(gate106inter3));
  inv1  gate193(.a(s_5), .O(gate106inter4));
  nand2 gate194(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate195(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate196(.a(N309), .O(gate106inter7));
  inv1  gate197(.a(N276), .O(gate106inter8));
  nand2 gate198(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate199(.a(s_5), .b(gate106inter3), .O(gate106inter10));
  nor2  gate200(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate201(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate202(.a(gate106inter12), .b(gate106inter1), .O(N337));

  xor2  gate315(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate316(.a(gate107inter0), .b(s_22), .O(gate107inter1));
  and2  gate317(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate318(.a(s_22), .O(gate107inter3));
  inv1  gate319(.a(s_23), .O(gate107inter4));
  nand2 gate320(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate321(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate322(.a(N319), .O(gate107inter7));
  inv1  gate323(.a(N34), .O(gate107inter8));
  nand2 gate324(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate325(.a(s_23), .b(gate107inter3), .O(gate107inter10));
  nor2  gate326(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate327(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate328(.a(gate107inter12), .b(gate107inter1), .O(N338));

  xor2  gate469(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate470(.a(gate108inter0), .b(s_44), .O(gate108inter1));
  and2  gate471(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate472(.a(s_44), .O(gate108inter3));
  inv1  gate473(.a(s_45), .O(gate108inter4));
  nand2 gate474(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate475(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate476(.a(N309), .O(gate108inter7));
  inv1  gate477(.a(N279), .O(gate108inter8));
  nand2 gate478(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate479(.a(s_45), .b(gate108inter3), .O(gate108inter10));
  nor2  gate480(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate481(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate482(.a(gate108inter12), .b(gate108inter1), .O(N339));
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate217(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate218(.a(gate111inter0), .b(s_8), .O(gate111inter1));
  and2  gate219(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate220(.a(s_8), .O(gate111inter3));
  inv1  gate221(.a(s_9), .O(gate111inter4));
  nand2 gate222(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate223(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate224(.a(N319), .O(gate111inter7));
  inv1  gate225(.a(N60), .O(gate111inter8));
  nand2 gate226(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate227(.a(s_9), .b(gate111inter3), .O(gate111inter10));
  nor2  gate228(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate229(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate230(.a(gate111inter12), .b(gate111inter1), .O(N342));

  xor2  gate259(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate260(.a(gate112inter0), .b(s_14), .O(gate112inter1));
  and2  gate261(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate262(.a(s_14), .O(gate112inter3));
  inv1  gate263(.a(s_15), .O(gate112inter4));
  nand2 gate264(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate265(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate266(.a(N309), .O(gate112inter7));
  inv1  gate267(.a(N285), .O(gate112inter8));
  nand2 gate268(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate269(.a(s_15), .b(gate112inter3), .O(gate112inter10));
  nor2  gate270(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate271(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate272(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );

  xor2  gate231(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate232(.a(gate114inter0), .b(s_10), .O(gate114inter1));
  and2  gate233(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate234(.a(s_10), .O(gate114inter3));
  inv1  gate235(.a(s_11), .O(gate114inter4));
  nand2 gate236(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate237(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate238(.a(N319), .O(gate114inter7));
  inv1  gate239(.a(N86), .O(gate114inter8));
  nand2 gate240(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate241(.a(s_11), .b(gate114inter3), .O(gate114inter10));
  nor2  gate242(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate243(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate244(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate301(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate302(.a(gate121inter0), .b(s_20), .O(gate121inter1));
  and2  gate303(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate304(.a(s_20), .O(gate121inter3));
  inv1  gate305(.a(s_21), .O(gate121inter4));
  nand2 gate306(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate307(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate308(.a(N335), .O(gate121inter7));
  inv1  gate309(.a(N304), .O(gate121inter8));
  nand2 gate310(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate311(.a(s_21), .b(gate121inter3), .O(gate121inter10));
  nor2  gate312(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate313(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate314(.a(gate121inter12), .b(gate121inter1), .O(N352));

  xor2  gate497(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate498(.a(gate122inter0), .b(s_48), .O(gate122inter1));
  and2  gate499(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate500(.a(s_48), .O(gate122inter3));
  inv1  gate501(.a(s_49), .O(gate122inter4));
  nand2 gate502(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate503(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate504(.a(N337), .O(gate122inter7));
  inv1  gate505(.a(N305), .O(gate122inter8));
  nand2 gate506(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate507(.a(s_49), .b(gate122inter3), .O(gate122inter10));
  nor2  gate508(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate509(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate510(.a(gate122inter12), .b(gate122inter1), .O(N353));
nand2 gate123( .a(N339), .b(N306), .O(N354) );

  xor2  gate455(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate456(.a(gate124inter0), .b(s_42), .O(gate124inter1));
  and2  gate457(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate458(.a(s_42), .O(gate124inter3));
  inv1  gate459(.a(s_43), .O(gate124inter4));
  nand2 gate460(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate461(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate462(.a(N341), .O(gate124inter7));
  inv1  gate463(.a(N307), .O(gate124inter8));
  nand2 gate464(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate465(.a(s_43), .b(gate124inter3), .O(gate124inter10));
  nor2  gate466(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate467(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate468(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );

  xor2  gate427(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate428(.a(gate133inter0), .b(s_38), .O(gate133inter1));
  and2  gate429(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate430(.a(s_38), .O(gate133inter3));
  inv1  gate431(.a(s_39), .O(gate133inter4));
  nand2 gate432(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate433(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate434(.a(N360), .O(gate133inter7));
  inv1  gate435(.a(N66), .O(gate133inter8));
  nand2 gate436(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate437(.a(s_39), .b(gate133inter3), .O(gate133inter10));
  nor2  gate438(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate439(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate440(.a(gate133inter12), .b(gate133inter1), .O(N375));
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule