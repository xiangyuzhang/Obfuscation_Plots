module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1415(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1416(.a(gate11inter0), .b(s_124), .O(gate11inter1));
  and2  gate1417(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1418(.a(s_124), .O(gate11inter3));
  inv1  gate1419(.a(s_125), .O(gate11inter4));
  nand2 gate1420(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1421(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1422(.a(G5), .O(gate11inter7));
  inv1  gate1423(.a(G6), .O(gate11inter8));
  nand2 gate1424(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1425(.a(s_125), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1426(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1427(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1428(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1695(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1696(.a(gate14inter0), .b(s_164), .O(gate14inter1));
  and2  gate1697(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1698(.a(s_164), .O(gate14inter3));
  inv1  gate1699(.a(s_165), .O(gate14inter4));
  nand2 gate1700(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1701(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1702(.a(G11), .O(gate14inter7));
  inv1  gate1703(.a(G12), .O(gate14inter8));
  nand2 gate1704(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1705(.a(s_165), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1706(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1707(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1708(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate2479(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2480(.a(gate15inter0), .b(s_276), .O(gate15inter1));
  and2  gate2481(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2482(.a(s_276), .O(gate15inter3));
  inv1  gate2483(.a(s_277), .O(gate15inter4));
  nand2 gate2484(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2485(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2486(.a(G13), .O(gate15inter7));
  inv1  gate2487(.a(G14), .O(gate15inter8));
  nand2 gate2488(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2489(.a(s_277), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2490(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2491(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2492(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1443(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1444(.a(gate17inter0), .b(s_128), .O(gate17inter1));
  and2  gate1445(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1446(.a(s_128), .O(gate17inter3));
  inv1  gate1447(.a(s_129), .O(gate17inter4));
  nand2 gate1448(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1449(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1450(.a(G17), .O(gate17inter7));
  inv1  gate1451(.a(G18), .O(gate17inter8));
  nand2 gate1452(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1453(.a(s_129), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1454(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1455(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1456(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2241(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2242(.a(gate19inter0), .b(s_242), .O(gate19inter1));
  and2  gate2243(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2244(.a(s_242), .O(gate19inter3));
  inv1  gate2245(.a(s_243), .O(gate19inter4));
  nand2 gate2246(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2247(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2248(.a(G21), .O(gate19inter7));
  inv1  gate2249(.a(G22), .O(gate19inter8));
  nand2 gate2250(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2251(.a(s_243), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2252(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2253(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2254(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1863(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1864(.a(gate28inter0), .b(s_188), .O(gate28inter1));
  and2  gate1865(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1866(.a(s_188), .O(gate28inter3));
  inv1  gate1867(.a(s_189), .O(gate28inter4));
  nand2 gate1868(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1869(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1870(.a(G10), .O(gate28inter7));
  inv1  gate1871(.a(G14), .O(gate28inter8));
  nand2 gate1872(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1873(.a(s_189), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1874(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1875(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1876(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1219(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1220(.a(gate33inter0), .b(s_96), .O(gate33inter1));
  and2  gate1221(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1222(.a(s_96), .O(gate33inter3));
  inv1  gate1223(.a(s_97), .O(gate33inter4));
  nand2 gate1224(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1225(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1226(.a(G17), .O(gate33inter7));
  inv1  gate1227(.a(G21), .O(gate33inter8));
  nand2 gate1228(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1229(.a(s_97), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1230(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1231(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1232(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2423(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2424(.a(gate34inter0), .b(s_268), .O(gate34inter1));
  and2  gate2425(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2426(.a(s_268), .O(gate34inter3));
  inv1  gate2427(.a(s_269), .O(gate34inter4));
  nand2 gate2428(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2429(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2430(.a(G25), .O(gate34inter7));
  inv1  gate2431(.a(G29), .O(gate34inter8));
  nand2 gate2432(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2433(.a(s_269), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2434(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2435(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2436(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1499(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1500(.a(gate36inter0), .b(s_136), .O(gate36inter1));
  and2  gate1501(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1502(.a(s_136), .O(gate36inter3));
  inv1  gate1503(.a(s_137), .O(gate36inter4));
  nand2 gate1504(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1505(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1506(.a(G26), .O(gate36inter7));
  inv1  gate1507(.a(G30), .O(gate36inter8));
  nand2 gate1508(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1509(.a(s_137), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1510(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1511(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1512(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate617(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate618(.a(gate39inter0), .b(s_10), .O(gate39inter1));
  and2  gate619(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate620(.a(s_10), .O(gate39inter3));
  inv1  gate621(.a(s_11), .O(gate39inter4));
  nand2 gate622(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate623(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate624(.a(G20), .O(gate39inter7));
  inv1  gate625(.a(G24), .O(gate39inter8));
  nand2 gate626(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate627(.a(s_11), .b(gate39inter3), .O(gate39inter10));
  nor2  gate628(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate629(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate630(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2087(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2088(.a(gate41inter0), .b(s_220), .O(gate41inter1));
  and2  gate2089(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2090(.a(s_220), .O(gate41inter3));
  inv1  gate2091(.a(s_221), .O(gate41inter4));
  nand2 gate2092(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2093(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2094(.a(G1), .O(gate41inter7));
  inv1  gate2095(.a(G266), .O(gate41inter8));
  nand2 gate2096(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2097(.a(s_221), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2098(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2099(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2100(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1429(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1430(.a(gate42inter0), .b(s_126), .O(gate42inter1));
  and2  gate1431(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1432(.a(s_126), .O(gate42inter3));
  inv1  gate1433(.a(s_127), .O(gate42inter4));
  nand2 gate1434(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1435(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1436(.a(G2), .O(gate42inter7));
  inv1  gate1437(.a(G266), .O(gate42inter8));
  nand2 gate1438(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1439(.a(s_127), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1440(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1441(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1442(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1233(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1234(.a(gate43inter0), .b(s_98), .O(gate43inter1));
  and2  gate1235(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1236(.a(s_98), .O(gate43inter3));
  inv1  gate1237(.a(s_99), .O(gate43inter4));
  nand2 gate1238(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1239(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1240(.a(G3), .O(gate43inter7));
  inv1  gate1241(.a(G269), .O(gate43inter8));
  nand2 gate1242(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1243(.a(s_99), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1244(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1245(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1246(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2507(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2508(.a(gate44inter0), .b(s_280), .O(gate44inter1));
  and2  gate2509(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2510(.a(s_280), .O(gate44inter3));
  inv1  gate2511(.a(s_281), .O(gate44inter4));
  nand2 gate2512(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2513(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2514(.a(G4), .O(gate44inter7));
  inv1  gate2515(.a(G269), .O(gate44inter8));
  nand2 gate2516(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2517(.a(s_281), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2518(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2519(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2520(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1107(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1108(.a(gate45inter0), .b(s_80), .O(gate45inter1));
  and2  gate1109(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1110(.a(s_80), .O(gate45inter3));
  inv1  gate1111(.a(s_81), .O(gate45inter4));
  nand2 gate1112(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1113(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1114(.a(G5), .O(gate45inter7));
  inv1  gate1115(.a(G272), .O(gate45inter8));
  nand2 gate1116(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1117(.a(s_81), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1118(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1119(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1120(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate841(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate842(.a(gate47inter0), .b(s_42), .O(gate47inter1));
  and2  gate843(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate844(.a(s_42), .O(gate47inter3));
  inv1  gate845(.a(s_43), .O(gate47inter4));
  nand2 gate846(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate847(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate848(.a(G7), .O(gate47inter7));
  inv1  gate849(.a(G275), .O(gate47inter8));
  nand2 gate850(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate851(.a(s_43), .b(gate47inter3), .O(gate47inter10));
  nor2  gate852(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate853(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate854(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate813(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate814(.a(gate51inter0), .b(s_38), .O(gate51inter1));
  and2  gate815(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate816(.a(s_38), .O(gate51inter3));
  inv1  gate817(.a(s_39), .O(gate51inter4));
  nand2 gate818(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate819(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate820(.a(G11), .O(gate51inter7));
  inv1  gate821(.a(G281), .O(gate51inter8));
  nand2 gate822(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate823(.a(s_39), .b(gate51inter3), .O(gate51inter10));
  nor2  gate824(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate825(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate826(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate645(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate646(.a(gate52inter0), .b(s_14), .O(gate52inter1));
  and2  gate647(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate648(.a(s_14), .O(gate52inter3));
  inv1  gate649(.a(s_15), .O(gate52inter4));
  nand2 gate650(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate651(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate652(.a(G12), .O(gate52inter7));
  inv1  gate653(.a(G281), .O(gate52inter8));
  nand2 gate654(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate655(.a(s_15), .b(gate52inter3), .O(gate52inter10));
  nor2  gate656(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate657(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate658(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1359(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1360(.a(gate57inter0), .b(s_116), .O(gate57inter1));
  and2  gate1361(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1362(.a(s_116), .O(gate57inter3));
  inv1  gate1363(.a(s_117), .O(gate57inter4));
  nand2 gate1364(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1365(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1366(.a(G17), .O(gate57inter7));
  inv1  gate1367(.a(G290), .O(gate57inter8));
  nand2 gate1368(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1369(.a(s_117), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1370(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1371(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1372(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1667(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1668(.a(gate58inter0), .b(s_160), .O(gate58inter1));
  and2  gate1669(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1670(.a(s_160), .O(gate58inter3));
  inv1  gate1671(.a(s_161), .O(gate58inter4));
  nand2 gate1672(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1673(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1674(.a(G18), .O(gate58inter7));
  inv1  gate1675(.a(G290), .O(gate58inter8));
  nand2 gate1676(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1677(.a(s_161), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1678(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1679(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1680(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate589(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate590(.a(gate59inter0), .b(s_6), .O(gate59inter1));
  and2  gate591(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate592(.a(s_6), .O(gate59inter3));
  inv1  gate593(.a(s_7), .O(gate59inter4));
  nand2 gate594(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate595(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate596(.a(G19), .O(gate59inter7));
  inv1  gate597(.a(G293), .O(gate59inter8));
  nand2 gate598(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate599(.a(s_7), .b(gate59inter3), .O(gate59inter10));
  nor2  gate600(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate601(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate602(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate981(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate982(.a(gate60inter0), .b(s_62), .O(gate60inter1));
  and2  gate983(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate984(.a(s_62), .O(gate60inter3));
  inv1  gate985(.a(s_63), .O(gate60inter4));
  nand2 gate986(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate987(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate988(.a(G20), .O(gate60inter7));
  inv1  gate989(.a(G293), .O(gate60inter8));
  nand2 gate990(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate991(.a(s_63), .b(gate60inter3), .O(gate60inter10));
  nor2  gate992(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate993(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate994(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1877(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1878(.a(gate61inter0), .b(s_190), .O(gate61inter1));
  and2  gate1879(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1880(.a(s_190), .O(gate61inter3));
  inv1  gate1881(.a(s_191), .O(gate61inter4));
  nand2 gate1882(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1883(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1884(.a(G21), .O(gate61inter7));
  inv1  gate1885(.a(G296), .O(gate61inter8));
  nand2 gate1886(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1887(.a(s_191), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1888(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1889(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1890(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1569(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1570(.a(gate63inter0), .b(s_146), .O(gate63inter1));
  and2  gate1571(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1572(.a(s_146), .O(gate63inter3));
  inv1  gate1573(.a(s_147), .O(gate63inter4));
  nand2 gate1574(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1575(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1576(.a(G23), .O(gate63inter7));
  inv1  gate1577(.a(G299), .O(gate63inter8));
  nand2 gate1578(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1579(.a(s_147), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1580(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1581(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1582(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1541(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1542(.a(gate67inter0), .b(s_142), .O(gate67inter1));
  and2  gate1543(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1544(.a(s_142), .O(gate67inter3));
  inv1  gate1545(.a(s_143), .O(gate67inter4));
  nand2 gate1546(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1547(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1548(.a(G27), .O(gate67inter7));
  inv1  gate1549(.a(G305), .O(gate67inter8));
  nand2 gate1550(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1551(.a(s_143), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1552(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1553(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1554(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1891(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1892(.a(gate70inter0), .b(s_192), .O(gate70inter1));
  and2  gate1893(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1894(.a(s_192), .O(gate70inter3));
  inv1  gate1895(.a(s_193), .O(gate70inter4));
  nand2 gate1896(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1897(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1898(.a(G30), .O(gate70inter7));
  inv1  gate1899(.a(G308), .O(gate70inter8));
  nand2 gate1900(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1901(.a(s_193), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1902(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1903(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1904(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2297(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2298(.a(gate72inter0), .b(s_250), .O(gate72inter1));
  and2  gate2299(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2300(.a(s_250), .O(gate72inter3));
  inv1  gate2301(.a(s_251), .O(gate72inter4));
  nand2 gate2302(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2303(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2304(.a(G32), .O(gate72inter7));
  inv1  gate2305(.a(G311), .O(gate72inter8));
  nand2 gate2306(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2307(.a(s_251), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2308(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2309(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2310(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1009(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1010(.a(gate74inter0), .b(s_66), .O(gate74inter1));
  and2  gate1011(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1012(.a(s_66), .O(gate74inter3));
  inv1  gate1013(.a(s_67), .O(gate74inter4));
  nand2 gate1014(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1015(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1016(.a(G5), .O(gate74inter7));
  inv1  gate1017(.a(G314), .O(gate74inter8));
  nand2 gate1018(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1019(.a(s_67), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1020(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1021(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1022(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2157(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2158(.a(gate76inter0), .b(s_230), .O(gate76inter1));
  and2  gate2159(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2160(.a(s_230), .O(gate76inter3));
  inv1  gate2161(.a(s_231), .O(gate76inter4));
  nand2 gate2162(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2163(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2164(.a(G13), .O(gate76inter7));
  inv1  gate2165(.a(G317), .O(gate76inter8));
  nand2 gate2166(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2167(.a(s_231), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2168(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2169(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2170(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1555(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1556(.a(gate78inter0), .b(s_144), .O(gate78inter1));
  and2  gate1557(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1558(.a(s_144), .O(gate78inter3));
  inv1  gate1559(.a(s_145), .O(gate78inter4));
  nand2 gate1560(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1561(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1562(.a(G6), .O(gate78inter7));
  inv1  gate1563(.a(G320), .O(gate78inter8));
  nand2 gate1564(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1565(.a(s_145), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1566(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1567(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1568(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2003(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2004(.a(gate80inter0), .b(s_208), .O(gate80inter1));
  and2  gate2005(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2006(.a(s_208), .O(gate80inter3));
  inv1  gate2007(.a(s_209), .O(gate80inter4));
  nand2 gate2008(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2009(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2010(.a(G14), .O(gate80inter7));
  inv1  gate2011(.a(G323), .O(gate80inter8));
  nand2 gate2012(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2013(.a(s_209), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2014(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2015(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2016(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1331(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1332(.a(gate81inter0), .b(s_112), .O(gate81inter1));
  and2  gate1333(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1334(.a(s_112), .O(gate81inter3));
  inv1  gate1335(.a(s_113), .O(gate81inter4));
  nand2 gate1336(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1337(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1338(.a(G3), .O(gate81inter7));
  inv1  gate1339(.a(G326), .O(gate81inter8));
  nand2 gate1340(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1341(.a(s_113), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1342(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1343(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1344(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2101(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2102(.a(gate84inter0), .b(s_222), .O(gate84inter1));
  and2  gate2103(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2104(.a(s_222), .O(gate84inter3));
  inv1  gate2105(.a(s_223), .O(gate84inter4));
  nand2 gate2106(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2107(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2108(.a(G15), .O(gate84inter7));
  inv1  gate2109(.a(G329), .O(gate84inter8));
  nand2 gate2110(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2111(.a(s_223), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2112(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2113(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2114(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1373(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1374(.a(gate88inter0), .b(s_118), .O(gate88inter1));
  and2  gate1375(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1376(.a(s_118), .O(gate88inter3));
  inv1  gate1377(.a(s_119), .O(gate88inter4));
  nand2 gate1378(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1379(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1380(.a(G16), .O(gate88inter7));
  inv1  gate1381(.a(G335), .O(gate88inter8));
  nand2 gate1382(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1383(.a(s_119), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1384(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1385(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1386(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1625(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1626(.a(gate90inter0), .b(s_154), .O(gate90inter1));
  and2  gate1627(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1628(.a(s_154), .O(gate90inter3));
  inv1  gate1629(.a(s_155), .O(gate90inter4));
  nand2 gate1630(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1631(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1632(.a(G21), .O(gate90inter7));
  inv1  gate1633(.a(G338), .O(gate90inter8));
  nand2 gate1634(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1635(.a(s_155), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1636(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1637(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1638(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1751(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1752(.a(gate91inter0), .b(s_172), .O(gate91inter1));
  and2  gate1753(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1754(.a(s_172), .O(gate91inter3));
  inv1  gate1755(.a(s_173), .O(gate91inter4));
  nand2 gate1756(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1757(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1758(.a(G25), .O(gate91inter7));
  inv1  gate1759(.a(G341), .O(gate91inter8));
  nand2 gate1760(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1761(.a(s_173), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1762(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1763(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1764(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2367(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2368(.a(gate92inter0), .b(s_260), .O(gate92inter1));
  and2  gate2369(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2370(.a(s_260), .O(gate92inter3));
  inv1  gate2371(.a(s_261), .O(gate92inter4));
  nand2 gate2372(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2373(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2374(.a(G29), .O(gate92inter7));
  inv1  gate2375(.a(G341), .O(gate92inter8));
  nand2 gate2376(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2377(.a(s_261), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2378(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2379(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2380(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1821(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1822(.a(gate96inter0), .b(s_182), .O(gate96inter1));
  and2  gate1823(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1824(.a(s_182), .O(gate96inter3));
  inv1  gate1825(.a(s_183), .O(gate96inter4));
  nand2 gate1826(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1827(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1828(.a(G30), .O(gate96inter7));
  inv1  gate1829(.a(G347), .O(gate96inter8));
  nand2 gate1830(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1831(.a(s_183), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1832(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1833(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1834(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2451(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2452(.a(gate100inter0), .b(s_272), .O(gate100inter1));
  and2  gate2453(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2454(.a(s_272), .O(gate100inter3));
  inv1  gate2455(.a(s_273), .O(gate100inter4));
  nand2 gate2456(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2457(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2458(.a(G31), .O(gate100inter7));
  inv1  gate2459(.a(G353), .O(gate100inter8));
  nand2 gate2460(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2461(.a(s_273), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2462(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2463(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2464(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate925(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate926(.a(gate102inter0), .b(s_54), .O(gate102inter1));
  and2  gate927(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate928(.a(s_54), .O(gate102inter3));
  inv1  gate929(.a(s_55), .O(gate102inter4));
  nand2 gate930(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate931(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate932(.a(G24), .O(gate102inter7));
  inv1  gate933(.a(G356), .O(gate102inter8));
  nand2 gate934(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate935(.a(s_55), .b(gate102inter3), .O(gate102inter10));
  nor2  gate936(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate937(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate938(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate2255(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2256(.a(gate103inter0), .b(s_244), .O(gate103inter1));
  and2  gate2257(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2258(.a(s_244), .O(gate103inter3));
  inv1  gate2259(.a(s_245), .O(gate103inter4));
  nand2 gate2260(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2261(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2262(.a(G28), .O(gate103inter7));
  inv1  gate2263(.a(G359), .O(gate103inter8));
  nand2 gate2264(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2265(.a(s_245), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2266(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2267(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2268(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2073(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2074(.a(gate104inter0), .b(s_218), .O(gate104inter1));
  and2  gate2075(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2076(.a(s_218), .O(gate104inter3));
  inv1  gate2077(.a(s_219), .O(gate104inter4));
  nand2 gate2078(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2079(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2080(.a(G32), .O(gate104inter7));
  inv1  gate2081(.a(G359), .O(gate104inter8));
  nand2 gate2082(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2083(.a(s_219), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2084(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2085(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2086(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate869(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate870(.a(gate106inter0), .b(s_46), .O(gate106inter1));
  and2  gate871(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate872(.a(s_46), .O(gate106inter3));
  inv1  gate873(.a(s_47), .O(gate106inter4));
  nand2 gate874(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate875(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate876(.a(G364), .O(gate106inter7));
  inv1  gate877(.a(G365), .O(gate106inter8));
  nand2 gate878(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate879(.a(s_47), .b(gate106inter3), .O(gate106inter10));
  nor2  gate880(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate881(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate882(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1037(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1038(.a(gate109inter0), .b(s_70), .O(gate109inter1));
  and2  gate1039(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1040(.a(s_70), .O(gate109inter3));
  inv1  gate1041(.a(s_71), .O(gate109inter4));
  nand2 gate1042(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1043(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1044(.a(G370), .O(gate109inter7));
  inv1  gate1045(.a(G371), .O(gate109inter8));
  nand2 gate1046(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1047(.a(s_71), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1048(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1049(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1050(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2199(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2200(.a(gate114inter0), .b(s_236), .O(gate114inter1));
  and2  gate2201(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2202(.a(s_236), .O(gate114inter3));
  inv1  gate2203(.a(s_237), .O(gate114inter4));
  nand2 gate2204(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2205(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2206(.a(G380), .O(gate114inter7));
  inv1  gate2207(.a(G381), .O(gate114inter8));
  nand2 gate2208(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2209(.a(s_237), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2210(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2211(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2212(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate897(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate898(.a(gate117inter0), .b(s_50), .O(gate117inter1));
  and2  gate899(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate900(.a(s_50), .O(gate117inter3));
  inv1  gate901(.a(s_51), .O(gate117inter4));
  nand2 gate902(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate903(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate904(.a(G386), .O(gate117inter7));
  inv1  gate905(.a(G387), .O(gate117inter8));
  nand2 gate906(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate907(.a(s_51), .b(gate117inter3), .O(gate117inter10));
  nor2  gate908(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate909(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate910(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate729(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate730(.a(gate122inter0), .b(s_26), .O(gate122inter1));
  and2  gate731(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate732(.a(s_26), .O(gate122inter3));
  inv1  gate733(.a(s_27), .O(gate122inter4));
  nand2 gate734(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate735(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate736(.a(G396), .O(gate122inter7));
  inv1  gate737(.a(G397), .O(gate122inter8));
  nand2 gate738(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate739(.a(s_27), .b(gate122inter3), .O(gate122inter10));
  nor2  gate740(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate741(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate742(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1191(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1192(.a(gate123inter0), .b(s_92), .O(gate123inter1));
  and2  gate1193(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1194(.a(s_92), .O(gate123inter3));
  inv1  gate1195(.a(s_93), .O(gate123inter4));
  nand2 gate1196(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1197(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1198(.a(G398), .O(gate123inter7));
  inv1  gate1199(.a(G399), .O(gate123inter8));
  nand2 gate1200(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1201(.a(s_93), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1202(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1203(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1204(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1933(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1934(.a(gate124inter0), .b(s_198), .O(gate124inter1));
  and2  gate1935(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1936(.a(s_198), .O(gate124inter3));
  inv1  gate1937(.a(s_199), .O(gate124inter4));
  nand2 gate1938(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1939(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1940(.a(G400), .O(gate124inter7));
  inv1  gate1941(.a(G401), .O(gate124inter8));
  nand2 gate1942(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1943(.a(s_199), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1944(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1945(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1946(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate883(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate884(.a(gate127inter0), .b(s_48), .O(gate127inter1));
  and2  gate885(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate886(.a(s_48), .O(gate127inter3));
  inv1  gate887(.a(s_49), .O(gate127inter4));
  nand2 gate888(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate889(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate890(.a(G406), .O(gate127inter7));
  inv1  gate891(.a(G407), .O(gate127inter8));
  nand2 gate892(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate893(.a(s_49), .b(gate127inter3), .O(gate127inter10));
  nor2  gate894(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate895(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate896(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1583(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1584(.a(gate132inter0), .b(s_148), .O(gate132inter1));
  and2  gate1585(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1586(.a(s_148), .O(gate132inter3));
  inv1  gate1587(.a(s_149), .O(gate132inter4));
  nand2 gate1588(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1589(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1590(.a(G416), .O(gate132inter7));
  inv1  gate1591(.a(G417), .O(gate132inter8));
  nand2 gate1592(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1593(.a(s_149), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1594(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1595(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1596(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1051(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1052(.a(gate133inter0), .b(s_72), .O(gate133inter1));
  and2  gate1053(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1054(.a(s_72), .O(gate133inter3));
  inv1  gate1055(.a(s_73), .O(gate133inter4));
  nand2 gate1056(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1057(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1058(.a(G418), .O(gate133inter7));
  inv1  gate1059(.a(G419), .O(gate133inter8));
  nand2 gate1060(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1061(.a(s_73), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1062(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1063(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1064(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2227(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2228(.a(gate136inter0), .b(s_240), .O(gate136inter1));
  and2  gate2229(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2230(.a(s_240), .O(gate136inter3));
  inv1  gate2231(.a(s_241), .O(gate136inter4));
  nand2 gate2232(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2233(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2234(.a(G424), .O(gate136inter7));
  inv1  gate2235(.a(G425), .O(gate136inter8));
  nand2 gate2236(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2237(.a(s_241), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2238(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2239(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2240(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate911(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate912(.a(gate137inter0), .b(s_52), .O(gate137inter1));
  and2  gate913(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate914(.a(s_52), .O(gate137inter3));
  inv1  gate915(.a(s_53), .O(gate137inter4));
  nand2 gate916(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate917(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate918(.a(G426), .O(gate137inter7));
  inv1  gate919(.a(G429), .O(gate137inter8));
  nand2 gate920(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate921(.a(s_53), .b(gate137inter3), .O(gate137inter10));
  nor2  gate922(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate923(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate924(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate967(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate968(.a(gate140inter0), .b(s_60), .O(gate140inter1));
  and2  gate969(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate970(.a(s_60), .O(gate140inter3));
  inv1  gate971(.a(s_61), .O(gate140inter4));
  nand2 gate972(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate973(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate974(.a(G444), .O(gate140inter7));
  inv1  gate975(.a(G447), .O(gate140inter8));
  nand2 gate976(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate977(.a(s_61), .b(gate140inter3), .O(gate140inter10));
  nor2  gate978(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate979(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate980(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1919(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1920(.a(gate145inter0), .b(s_196), .O(gate145inter1));
  and2  gate1921(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1922(.a(s_196), .O(gate145inter3));
  inv1  gate1923(.a(s_197), .O(gate145inter4));
  nand2 gate1924(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1925(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1926(.a(G474), .O(gate145inter7));
  inv1  gate1927(.a(G477), .O(gate145inter8));
  nand2 gate1928(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1929(.a(s_197), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1930(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1931(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1932(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2059(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2060(.a(gate147inter0), .b(s_216), .O(gate147inter1));
  and2  gate2061(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2062(.a(s_216), .O(gate147inter3));
  inv1  gate2063(.a(s_217), .O(gate147inter4));
  nand2 gate2064(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2065(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2066(.a(G486), .O(gate147inter7));
  inv1  gate2067(.a(G489), .O(gate147inter8));
  nand2 gate2068(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2069(.a(s_217), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2070(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2071(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2072(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate785(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate786(.a(gate149inter0), .b(s_34), .O(gate149inter1));
  and2  gate787(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate788(.a(s_34), .O(gate149inter3));
  inv1  gate789(.a(s_35), .O(gate149inter4));
  nand2 gate790(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate791(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate792(.a(G498), .O(gate149inter7));
  inv1  gate793(.a(G501), .O(gate149inter8));
  nand2 gate794(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate795(.a(s_35), .b(gate149inter3), .O(gate149inter10));
  nor2  gate796(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate797(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate798(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2493(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2494(.a(gate153inter0), .b(s_278), .O(gate153inter1));
  and2  gate2495(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2496(.a(s_278), .O(gate153inter3));
  inv1  gate2497(.a(s_279), .O(gate153inter4));
  nand2 gate2498(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2499(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2500(.a(G426), .O(gate153inter7));
  inv1  gate2501(.a(G522), .O(gate153inter8));
  nand2 gate2502(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2503(.a(s_279), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2504(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2505(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2506(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2381(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2382(.a(gate154inter0), .b(s_262), .O(gate154inter1));
  and2  gate2383(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2384(.a(s_262), .O(gate154inter3));
  inv1  gate2385(.a(s_263), .O(gate154inter4));
  nand2 gate2386(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2387(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2388(.a(G429), .O(gate154inter7));
  inv1  gate2389(.a(G522), .O(gate154inter8));
  nand2 gate2390(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2391(.a(s_263), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2392(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2393(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2394(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate687(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate688(.a(gate157inter0), .b(s_20), .O(gate157inter1));
  and2  gate689(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate690(.a(s_20), .O(gate157inter3));
  inv1  gate691(.a(s_21), .O(gate157inter4));
  nand2 gate692(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate693(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate694(.a(G438), .O(gate157inter7));
  inv1  gate695(.a(G528), .O(gate157inter8));
  nand2 gate696(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate697(.a(s_21), .b(gate157inter3), .O(gate157inter10));
  nor2  gate698(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate699(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate700(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate757(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate758(.a(gate162inter0), .b(s_30), .O(gate162inter1));
  and2  gate759(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate760(.a(s_30), .O(gate162inter3));
  inv1  gate761(.a(s_31), .O(gate162inter4));
  nand2 gate762(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate763(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate764(.a(G453), .O(gate162inter7));
  inv1  gate765(.a(G534), .O(gate162inter8));
  nand2 gate766(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate767(.a(s_31), .b(gate162inter3), .O(gate162inter10));
  nor2  gate768(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate769(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate770(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1835(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1836(.a(gate164inter0), .b(s_184), .O(gate164inter1));
  and2  gate1837(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1838(.a(s_184), .O(gate164inter3));
  inv1  gate1839(.a(s_185), .O(gate164inter4));
  nand2 gate1840(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1841(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1842(.a(G459), .O(gate164inter7));
  inv1  gate1843(.a(G537), .O(gate164inter8));
  nand2 gate1844(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1845(.a(s_185), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1846(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1847(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1848(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate575(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate576(.a(gate166inter0), .b(s_4), .O(gate166inter1));
  and2  gate577(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate578(.a(s_4), .O(gate166inter3));
  inv1  gate579(.a(s_5), .O(gate166inter4));
  nand2 gate580(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate581(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate582(.a(G465), .O(gate166inter7));
  inv1  gate583(.a(G540), .O(gate166inter8));
  nand2 gate584(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate585(.a(s_5), .b(gate166inter3), .O(gate166inter10));
  nor2  gate586(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate587(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate588(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2437(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2438(.a(gate172inter0), .b(s_270), .O(gate172inter1));
  and2  gate2439(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2440(.a(s_270), .O(gate172inter3));
  inv1  gate2441(.a(s_271), .O(gate172inter4));
  nand2 gate2442(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2443(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2444(.a(G483), .O(gate172inter7));
  inv1  gate2445(.a(G549), .O(gate172inter8));
  nand2 gate2446(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2447(.a(s_271), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2448(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2449(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2450(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1289(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1290(.a(gate174inter0), .b(s_106), .O(gate174inter1));
  and2  gate1291(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1292(.a(s_106), .O(gate174inter3));
  inv1  gate1293(.a(s_107), .O(gate174inter4));
  nand2 gate1294(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1295(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1296(.a(G489), .O(gate174inter7));
  inv1  gate1297(.a(G552), .O(gate174inter8));
  nand2 gate1298(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1299(.a(s_107), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1300(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1301(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1302(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1905(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1906(.a(gate175inter0), .b(s_194), .O(gate175inter1));
  and2  gate1907(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1908(.a(s_194), .O(gate175inter3));
  inv1  gate1909(.a(s_195), .O(gate175inter4));
  nand2 gate1910(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1911(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1912(.a(G492), .O(gate175inter7));
  inv1  gate1913(.a(G555), .O(gate175inter8));
  nand2 gate1914(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1915(.a(s_195), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1916(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1917(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1918(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1723(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1724(.a(gate176inter0), .b(s_168), .O(gate176inter1));
  and2  gate1725(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1726(.a(s_168), .O(gate176inter3));
  inv1  gate1727(.a(s_169), .O(gate176inter4));
  nand2 gate1728(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1729(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1730(.a(G495), .O(gate176inter7));
  inv1  gate1731(.a(G555), .O(gate176inter8));
  nand2 gate1732(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1733(.a(s_169), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1734(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1735(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1736(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate701(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate702(.a(gate178inter0), .b(s_22), .O(gate178inter1));
  and2  gate703(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate704(.a(s_22), .O(gate178inter3));
  inv1  gate705(.a(s_23), .O(gate178inter4));
  nand2 gate706(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate707(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate708(.a(G501), .O(gate178inter7));
  inv1  gate709(.a(G558), .O(gate178inter8));
  nand2 gate710(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate711(.a(s_23), .b(gate178inter3), .O(gate178inter10));
  nor2  gate712(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate713(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate714(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1401(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1402(.a(gate182inter0), .b(s_122), .O(gate182inter1));
  and2  gate1403(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1404(.a(s_122), .O(gate182inter3));
  inv1  gate1405(.a(s_123), .O(gate182inter4));
  nand2 gate1406(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1407(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1408(.a(G513), .O(gate182inter7));
  inv1  gate1409(.a(G564), .O(gate182inter8));
  nand2 gate1410(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1411(.a(s_123), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1412(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1413(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1414(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2325(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2326(.a(gate190inter0), .b(s_254), .O(gate190inter1));
  and2  gate2327(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2328(.a(s_254), .O(gate190inter3));
  inv1  gate2329(.a(s_255), .O(gate190inter4));
  nand2 gate2330(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2331(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2332(.a(G580), .O(gate190inter7));
  inv1  gate2333(.a(G581), .O(gate190inter8));
  nand2 gate2334(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2335(.a(s_255), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2336(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2337(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2338(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1163(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1164(.a(gate192inter0), .b(s_88), .O(gate192inter1));
  and2  gate1165(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1166(.a(s_88), .O(gate192inter3));
  inv1  gate1167(.a(s_89), .O(gate192inter4));
  nand2 gate1168(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1169(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1170(.a(G584), .O(gate192inter7));
  inv1  gate1171(.a(G585), .O(gate192inter8));
  nand2 gate1172(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1173(.a(s_89), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1174(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1175(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1176(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate2213(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2214(.a(gate199inter0), .b(s_238), .O(gate199inter1));
  and2  gate2215(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2216(.a(s_238), .O(gate199inter3));
  inv1  gate2217(.a(s_239), .O(gate199inter4));
  nand2 gate2218(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2219(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2220(.a(G598), .O(gate199inter7));
  inv1  gate2221(.a(G599), .O(gate199inter8));
  nand2 gate2222(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2223(.a(s_239), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2224(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2225(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2226(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1387(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1388(.a(gate200inter0), .b(s_120), .O(gate200inter1));
  and2  gate1389(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1390(.a(s_120), .O(gate200inter3));
  inv1  gate1391(.a(s_121), .O(gate200inter4));
  nand2 gate1392(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1393(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1394(.a(G600), .O(gate200inter7));
  inv1  gate1395(.a(G601), .O(gate200inter8));
  nand2 gate1396(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1397(.a(s_121), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1398(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1399(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1400(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1205(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1206(.a(gate207inter0), .b(s_94), .O(gate207inter1));
  and2  gate1207(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1208(.a(s_94), .O(gate207inter3));
  inv1  gate1209(.a(s_95), .O(gate207inter4));
  nand2 gate1210(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1211(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1212(.a(G622), .O(gate207inter7));
  inv1  gate1213(.a(G632), .O(gate207inter8));
  nand2 gate1214(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1215(.a(s_95), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1216(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1217(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1218(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2465(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2466(.a(gate216inter0), .b(s_274), .O(gate216inter1));
  and2  gate2467(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2468(.a(s_274), .O(gate216inter3));
  inv1  gate2469(.a(s_275), .O(gate216inter4));
  nand2 gate2470(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2471(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2472(.a(G617), .O(gate216inter7));
  inv1  gate2473(.a(G675), .O(gate216inter8));
  nand2 gate2474(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2475(.a(s_275), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2476(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2477(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2478(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1345(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1346(.a(gate217inter0), .b(s_114), .O(gate217inter1));
  and2  gate1347(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1348(.a(s_114), .O(gate217inter3));
  inv1  gate1349(.a(s_115), .O(gate217inter4));
  nand2 gate1350(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1351(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1352(.a(G622), .O(gate217inter7));
  inv1  gate1353(.a(G678), .O(gate217inter8));
  nand2 gate1354(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1355(.a(s_115), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1356(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1357(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1358(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate995(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate996(.a(gate219inter0), .b(s_64), .O(gate219inter1));
  and2  gate997(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate998(.a(s_64), .O(gate219inter3));
  inv1  gate999(.a(s_65), .O(gate219inter4));
  nand2 gate1000(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1001(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1002(.a(G632), .O(gate219inter7));
  inv1  gate1003(.a(G681), .O(gate219inter8));
  nand2 gate1004(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1005(.a(s_65), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1006(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1007(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1008(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1261(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1262(.a(gate221inter0), .b(s_102), .O(gate221inter1));
  and2  gate1263(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1264(.a(s_102), .O(gate221inter3));
  inv1  gate1265(.a(s_103), .O(gate221inter4));
  nand2 gate1266(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1267(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1268(.a(G622), .O(gate221inter7));
  inv1  gate1269(.a(G684), .O(gate221inter8));
  nand2 gate1270(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1271(.a(s_103), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1272(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1273(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1274(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1765(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1766(.a(gate222inter0), .b(s_174), .O(gate222inter1));
  and2  gate1767(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1768(.a(s_174), .O(gate222inter3));
  inv1  gate1769(.a(s_175), .O(gate222inter4));
  nand2 gate1770(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1771(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1772(.a(G632), .O(gate222inter7));
  inv1  gate1773(.a(G684), .O(gate222inter8));
  nand2 gate1774(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1775(.a(s_175), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1776(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1777(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1778(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1975(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1976(.a(gate224inter0), .b(s_204), .O(gate224inter1));
  and2  gate1977(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1978(.a(s_204), .O(gate224inter3));
  inv1  gate1979(.a(s_205), .O(gate224inter4));
  nand2 gate1980(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1981(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1982(.a(G637), .O(gate224inter7));
  inv1  gate1983(.a(G687), .O(gate224inter8));
  nand2 gate1984(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1985(.a(s_205), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1986(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1987(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1988(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate673(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate674(.a(gate226inter0), .b(s_18), .O(gate226inter1));
  and2  gate675(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate676(.a(s_18), .O(gate226inter3));
  inv1  gate677(.a(s_19), .O(gate226inter4));
  nand2 gate678(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate679(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate680(.a(G692), .O(gate226inter7));
  inv1  gate681(.a(G693), .O(gate226inter8));
  nand2 gate682(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate683(.a(s_19), .b(gate226inter3), .O(gate226inter10));
  nor2  gate684(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate685(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate686(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate547(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate548(.a(gate228inter0), .b(s_0), .O(gate228inter1));
  and2  gate549(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate550(.a(s_0), .O(gate228inter3));
  inv1  gate551(.a(s_1), .O(gate228inter4));
  nand2 gate552(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate553(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate554(.a(G696), .O(gate228inter7));
  inv1  gate555(.a(G697), .O(gate228inter8));
  nand2 gate556(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate557(.a(s_1), .b(gate228inter3), .O(gate228inter10));
  nor2  gate558(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate559(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate560(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2045(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2046(.a(gate233inter0), .b(s_214), .O(gate233inter1));
  and2  gate2047(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2048(.a(s_214), .O(gate233inter3));
  inv1  gate2049(.a(s_215), .O(gate233inter4));
  nand2 gate2050(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2051(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2052(.a(G242), .O(gate233inter7));
  inv1  gate2053(.a(G718), .O(gate233inter8));
  nand2 gate2054(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2055(.a(s_215), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2056(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2057(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2058(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2339(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2340(.a(gate237inter0), .b(s_256), .O(gate237inter1));
  and2  gate2341(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2342(.a(s_256), .O(gate237inter3));
  inv1  gate2343(.a(s_257), .O(gate237inter4));
  nand2 gate2344(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2345(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2346(.a(G254), .O(gate237inter7));
  inv1  gate2347(.a(G706), .O(gate237inter8));
  nand2 gate2348(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2349(.a(s_257), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2350(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2351(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2352(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate771(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate772(.a(gate239inter0), .b(s_32), .O(gate239inter1));
  and2  gate773(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate774(.a(s_32), .O(gate239inter3));
  inv1  gate775(.a(s_33), .O(gate239inter4));
  nand2 gate776(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate777(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate778(.a(G260), .O(gate239inter7));
  inv1  gate779(.a(G712), .O(gate239inter8));
  nand2 gate780(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate781(.a(s_33), .b(gate239inter3), .O(gate239inter10));
  nor2  gate782(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate783(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate784(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate2185(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2186(.a(gate240inter0), .b(s_234), .O(gate240inter1));
  and2  gate2187(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2188(.a(s_234), .O(gate240inter3));
  inv1  gate2189(.a(s_235), .O(gate240inter4));
  nand2 gate2190(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2191(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2192(.a(G263), .O(gate240inter7));
  inv1  gate2193(.a(G715), .O(gate240inter8));
  nand2 gate2194(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2195(.a(s_235), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2196(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2197(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2198(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate855(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate856(.a(gate241inter0), .b(s_44), .O(gate241inter1));
  and2  gate857(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate858(.a(s_44), .O(gate241inter3));
  inv1  gate859(.a(s_45), .O(gate241inter4));
  nand2 gate860(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate861(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate862(.a(G242), .O(gate241inter7));
  inv1  gate863(.a(G730), .O(gate241inter8));
  nand2 gate864(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate865(.a(s_45), .b(gate241inter3), .O(gate241inter10));
  nor2  gate866(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate867(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate868(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1023(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1024(.a(gate243inter0), .b(s_68), .O(gate243inter1));
  and2  gate1025(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1026(.a(s_68), .O(gate243inter3));
  inv1  gate1027(.a(s_69), .O(gate243inter4));
  nand2 gate1028(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1029(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1030(.a(G245), .O(gate243inter7));
  inv1  gate1031(.a(G733), .O(gate243inter8));
  nand2 gate1032(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1033(.a(s_69), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1034(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1035(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1036(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1737(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1738(.a(gate251inter0), .b(s_170), .O(gate251inter1));
  and2  gate1739(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1740(.a(s_170), .O(gate251inter3));
  inv1  gate1741(.a(s_171), .O(gate251inter4));
  nand2 gate1742(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1743(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1744(.a(G257), .O(gate251inter7));
  inv1  gate1745(.a(G745), .O(gate251inter8));
  nand2 gate1746(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1747(.a(s_171), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1748(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1749(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1750(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1709(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1710(.a(gate253inter0), .b(s_166), .O(gate253inter1));
  and2  gate1711(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1712(.a(s_166), .O(gate253inter3));
  inv1  gate1713(.a(s_167), .O(gate253inter4));
  nand2 gate1714(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1715(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1716(.a(G260), .O(gate253inter7));
  inv1  gate1717(.a(G748), .O(gate253inter8));
  nand2 gate1718(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1719(.a(s_167), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1720(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1721(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1722(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate743(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate744(.a(gate254inter0), .b(s_28), .O(gate254inter1));
  and2  gate745(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate746(.a(s_28), .O(gate254inter3));
  inv1  gate747(.a(s_29), .O(gate254inter4));
  nand2 gate748(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate749(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate750(.a(G712), .O(gate254inter7));
  inv1  gate751(.a(G748), .O(gate254inter8));
  nand2 gate752(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate753(.a(s_29), .b(gate254inter3), .O(gate254inter10));
  nor2  gate754(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate755(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate756(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1079(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1080(.a(gate257inter0), .b(s_76), .O(gate257inter1));
  and2  gate1081(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1082(.a(s_76), .O(gate257inter3));
  inv1  gate1083(.a(s_77), .O(gate257inter4));
  nand2 gate1084(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1085(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1086(.a(G754), .O(gate257inter7));
  inv1  gate1087(.a(G755), .O(gate257inter8));
  nand2 gate1088(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1089(.a(s_77), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1090(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1091(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1092(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1177(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1178(.a(gate258inter0), .b(s_90), .O(gate258inter1));
  and2  gate1179(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1180(.a(s_90), .O(gate258inter3));
  inv1  gate1181(.a(s_91), .O(gate258inter4));
  nand2 gate1182(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1183(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1184(.a(G756), .O(gate258inter7));
  inv1  gate1185(.a(G757), .O(gate258inter8));
  nand2 gate1186(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1187(.a(s_91), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1188(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1189(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1190(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1485(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1486(.a(gate260inter0), .b(s_134), .O(gate260inter1));
  and2  gate1487(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1488(.a(s_134), .O(gate260inter3));
  inv1  gate1489(.a(s_135), .O(gate260inter4));
  nand2 gate1490(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1491(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1492(.a(G760), .O(gate260inter7));
  inv1  gate1493(.a(G761), .O(gate260inter8));
  nand2 gate1494(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1495(.a(s_135), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1496(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1497(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1498(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2311(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2312(.a(gate263inter0), .b(s_252), .O(gate263inter1));
  and2  gate2313(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2314(.a(s_252), .O(gate263inter3));
  inv1  gate2315(.a(s_253), .O(gate263inter4));
  nand2 gate2316(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2317(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2318(.a(G766), .O(gate263inter7));
  inv1  gate2319(.a(G767), .O(gate263inter8));
  nand2 gate2320(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2321(.a(s_253), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2322(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2323(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2324(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate2283(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2284(.a(gate266inter0), .b(s_248), .O(gate266inter1));
  and2  gate2285(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2286(.a(s_248), .O(gate266inter3));
  inv1  gate2287(.a(s_249), .O(gate266inter4));
  nand2 gate2288(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2289(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2290(.a(G645), .O(gate266inter7));
  inv1  gate2291(.a(G773), .O(gate266inter8));
  nand2 gate2292(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2293(.a(s_249), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2294(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2295(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2296(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate827(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate828(.a(gate267inter0), .b(s_40), .O(gate267inter1));
  and2  gate829(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate830(.a(s_40), .O(gate267inter3));
  inv1  gate831(.a(s_41), .O(gate267inter4));
  nand2 gate832(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate833(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate834(.a(G648), .O(gate267inter7));
  inv1  gate835(.a(G776), .O(gate267inter8));
  nand2 gate836(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate837(.a(s_41), .b(gate267inter3), .O(gate267inter10));
  nor2  gate838(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate839(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate840(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate953(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate954(.a(gate268inter0), .b(s_58), .O(gate268inter1));
  and2  gate955(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate956(.a(s_58), .O(gate268inter3));
  inv1  gate957(.a(s_59), .O(gate268inter4));
  nand2 gate958(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate959(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate960(.a(G651), .O(gate268inter7));
  inv1  gate961(.a(G779), .O(gate268inter8));
  nand2 gate962(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate963(.a(s_59), .b(gate268inter3), .O(gate268inter10));
  nor2  gate964(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate965(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate966(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1121(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1122(.a(gate270inter0), .b(s_82), .O(gate270inter1));
  and2  gate1123(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1124(.a(s_82), .O(gate270inter3));
  inv1  gate1125(.a(s_83), .O(gate270inter4));
  nand2 gate1126(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1127(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1128(.a(G657), .O(gate270inter7));
  inv1  gate1129(.a(G785), .O(gate270inter8));
  nand2 gate1130(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1131(.a(s_83), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1132(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1133(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1134(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2353(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2354(.a(gate274inter0), .b(s_258), .O(gate274inter1));
  and2  gate2355(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2356(.a(s_258), .O(gate274inter3));
  inv1  gate2357(.a(s_259), .O(gate274inter4));
  nand2 gate2358(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2359(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2360(.a(G770), .O(gate274inter7));
  inv1  gate2361(.a(G794), .O(gate274inter8));
  nand2 gate2362(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2363(.a(s_259), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2364(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2365(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2366(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2031(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2032(.a(gate275inter0), .b(s_212), .O(gate275inter1));
  and2  gate2033(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2034(.a(s_212), .O(gate275inter3));
  inv1  gate2035(.a(s_213), .O(gate275inter4));
  nand2 gate2036(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2037(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2038(.a(G645), .O(gate275inter7));
  inv1  gate2039(.a(G797), .O(gate275inter8));
  nand2 gate2040(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2041(.a(s_213), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2042(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2043(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2044(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1681(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1682(.a(gate277inter0), .b(s_162), .O(gate277inter1));
  and2  gate1683(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1684(.a(s_162), .O(gate277inter3));
  inv1  gate1685(.a(s_163), .O(gate277inter4));
  nand2 gate1686(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1687(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1688(.a(G648), .O(gate277inter7));
  inv1  gate1689(.a(G800), .O(gate277inter8));
  nand2 gate1690(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1691(.a(s_163), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1692(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1693(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1694(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2115(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2116(.a(gate280inter0), .b(s_224), .O(gate280inter1));
  and2  gate2117(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2118(.a(s_224), .O(gate280inter3));
  inv1  gate2119(.a(s_225), .O(gate280inter4));
  nand2 gate2120(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2121(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2122(.a(G779), .O(gate280inter7));
  inv1  gate2123(.a(G803), .O(gate280inter8));
  nand2 gate2124(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2125(.a(s_225), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2126(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2127(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2128(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1793(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1794(.a(gate283inter0), .b(s_178), .O(gate283inter1));
  and2  gate1795(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1796(.a(s_178), .O(gate283inter3));
  inv1  gate1797(.a(s_179), .O(gate283inter4));
  nand2 gate1798(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1799(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1800(.a(G657), .O(gate283inter7));
  inv1  gate1801(.a(G809), .O(gate283inter8));
  nand2 gate1802(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1803(.a(s_179), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1804(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1805(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1806(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate2017(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2018(.a(gate284inter0), .b(s_210), .O(gate284inter1));
  and2  gate2019(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2020(.a(s_210), .O(gate284inter3));
  inv1  gate2021(.a(s_211), .O(gate284inter4));
  nand2 gate2022(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2023(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2024(.a(G785), .O(gate284inter7));
  inv1  gate2025(.a(G809), .O(gate284inter8));
  nand2 gate2026(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2027(.a(s_211), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2028(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2029(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2030(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate939(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate940(.a(gate286inter0), .b(s_56), .O(gate286inter1));
  and2  gate941(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate942(.a(s_56), .O(gate286inter3));
  inv1  gate943(.a(s_57), .O(gate286inter4));
  nand2 gate944(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate945(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate946(.a(G788), .O(gate286inter7));
  inv1  gate947(.a(G812), .O(gate286inter8));
  nand2 gate948(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate949(.a(s_57), .b(gate286inter3), .O(gate286inter10));
  nor2  gate950(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate951(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate952(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1275(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1276(.a(gate289inter0), .b(s_104), .O(gate289inter1));
  and2  gate1277(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1278(.a(s_104), .O(gate289inter3));
  inv1  gate1279(.a(s_105), .O(gate289inter4));
  nand2 gate1280(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1281(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1282(.a(G818), .O(gate289inter7));
  inv1  gate1283(.a(G819), .O(gate289inter8));
  nand2 gate1284(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1285(.a(s_105), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1286(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1287(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1288(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1471(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1472(.a(gate291inter0), .b(s_132), .O(gate291inter1));
  and2  gate1473(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1474(.a(s_132), .O(gate291inter3));
  inv1  gate1475(.a(s_133), .O(gate291inter4));
  nand2 gate1476(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1477(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1478(.a(G822), .O(gate291inter7));
  inv1  gate1479(.a(G823), .O(gate291inter8));
  nand2 gate1480(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1481(.a(s_133), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1482(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1483(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1484(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1611(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1612(.a(gate295inter0), .b(s_152), .O(gate295inter1));
  and2  gate1613(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1614(.a(s_152), .O(gate295inter3));
  inv1  gate1615(.a(s_153), .O(gate295inter4));
  nand2 gate1616(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1617(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1618(.a(G830), .O(gate295inter7));
  inv1  gate1619(.a(G831), .O(gate295inter8));
  nand2 gate1620(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1621(.a(s_153), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1622(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1623(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1624(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1639(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1640(.a(gate296inter0), .b(s_156), .O(gate296inter1));
  and2  gate1641(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1642(.a(s_156), .O(gate296inter3));
  inv1  gate1643(.a(s_157), .O(gate296inter4));
  nand2 gate1644(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1645(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1646(.a(G826), .O(gate296inter7));
  inv1  gate1647(.a(G827), .O(gate296inter8));
  nand2 gate1648(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1649(.a(s_157), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1650(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1651(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1652(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2395(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2396(.a(gate388inter0), .b(s_264), .O(gate388inter1));
  and2  gate2397(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2398(.a(s_264), .O(gate388inter3));
  inv1  gate2399(.a(s_265), .O(gate388inter4));
  nand2 gate2400(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2401(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2402(.a(G2), .O(gate388inter7));
  inv1  gate2403(.a(G1039), .O(gate388inter8));
  nand2 gate2404(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2405(.a(s_265), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2406(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2407(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2408(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1247(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1248(.a(gate389inter0), .b(s_100), .O(gate389inter1));
  and2  gate1249(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1250(.a(s_100), .O(gate389inter3));
  inv1  gate1251(.a(s_101), .O(gate389inter4));
  nand2 gate1252(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1253(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1254(.a(G3), .O(gate389inter7));
  inv1  gate1255(.a(G1042), .O(gate389inter8));
  nand2 gate1256(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1257(.a(s_101), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1258(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1259(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1260(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1317(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1318(.a(gate391inter0), .b(s_110), .O(gate391inter1));
  and2  gate1319(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1320(.a(s_110), .O(gate391inter3));
  inv1  gate1321(.a(s_111), .O(gate391inter4));
  nand2 gate1322(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1323(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1324(.a(G5), .O(gate391inter7));
  inv1  gate1325(.a(G1048), .O(gate391inter8));
  nand2 gate1326(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1327(.a(s_111), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1328(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1329(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1330(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1513(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1514(.a(gate399inter0), .b(s_138), .O(gate399inter1));
  and2  gate1515(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1516(.a(s_138), .O(gate399inter3));
  inv1  gate1517(.a(s_139), .O(gate399inter4));
  nand2 gate1518(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1519(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1520(.a(G13), .O(gate399inter7));
  inv1  gate1521(.a(G1072), .O(gate399inter8));
  nand2 gate1522(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1523(.a(s_139), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1524(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1525(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1526(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1653(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1654(.a(gate401inter0), .b(s_158), .O(gate401inter1));
  and2  gate1655(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1656(.a(s_158), .O(gate401inter3));
  inv1  gate1657(.a(s_159), .O(gate401inter4));
  nand2 gate1658(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1659(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1660(.a(G15), .O(gate401inter7));
  inv1  gate1661(.a(G1078), .O(gate401inter8));
  nand2 gate1662(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1663(.a(s_159), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1664(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1665(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1666(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1849(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1850(.a(gate402inter0), .b(s_186), .O(gate402inter1));
  and2  gate1851(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1852(.a(s_186), .O(gate402inter3));
  inv1  gate1853(.a(s_187), .O(gate402inter4));
  nand2 gate1854(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1855(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1856(.a(G16), .O(gate402inter7));
  inv1  gate1857(.a(G1081), .O(gate402inter8));
  nand2 gate1858(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1859(.a(s_187), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1860(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1861(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1862(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate715(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate716(.a(gate409inter0), .b(s_24), .O(gate409inter1));
  and2  gate717(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate718(.a(s_24), .O(gate409inter3));
  inv1  gate719(.a(s_25), .O(gate409inter4));
  nand2 gate720(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate721(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate722(.a(G23), .O(gate409inter7));
  inv1  gate723(.a(G1102), .O(gate409inter8));
  nand2 gate724(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate725(.a(s_25), .b(gate409inter3), .O(gate409inter10));
  nor2  gate726(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate727(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate728(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1135(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1136(.a(gate420inter0), .b(s_84), .O(gate420inter1));
  and2  gate1137(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1138(.a(s_84), .O(gate420inter3));
  inv1  gate1139(.a(s_85), .O(gate420inter4));
  nand2 gate1140(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1141(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1142(.a(G1036), .O(gate420inter7));
  inv1  gate1143(.a(G1132), .O(gate420inter8));
  nand2 gate1144(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1145(.a(s_85), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1146(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1147(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1148(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1093(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1094(.a(gate423inter0), .b(s_78), .O(gate423inter1));
  and2  gate1095(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1096(.a(s_78), .O(gate423inter3));
  inv1  gate1097(.a(s_79), .O(gate423inter4));
  nand2 gate1098(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1099(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1100(.a(G3), .O(gate423inter7));
  inv1  gate1101(.a(G1138), .O(gate423inter8));
  nand2 gate1102(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1103(.a(s_79), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1104(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1105(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1106(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1149(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1150(.a(gate428inter0), .b(s_86), .O(gate428inter1));
  and2  gate1151(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1152(.a(s_86), .O(gate428inter3));
  inv1  gate1153(.a(s_87), .O(gate428inter4));
  nand2 gate1154(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1155(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1156(.a(G1048), .O(gate428inter7));
  inv1  gate1157(.a(G1144), .O(gate428inter8));
  nand2 gate1158(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1159(.a(s_87), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1160(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1161(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1162(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2269(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2270(.a(gate438inter0), .b(s_246), .O(gate438inter1));
  and2  gate2271(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2272(.a(s_246), .O(gate438inter3));
  inv1  gate2273(.a(s_247), .O(gate438inter4));
  nand2 gate2274(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2275(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2276(.a(G1063), .O(gate438inter7));
  inv1  gate2277(.a(G1159), .O(gate438inter8));
  nand2 gate2278(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2279(.a(s_247), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2280(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2281(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2282(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate2129(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2130(.a(gate439inter0), .b(s_226), .O(gate439inter1));
  and2  gate2131(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2132(.a(s_226), .O(gate439inter3));
  inv1  gate2133(.a(s_227), .O(gate439inter4));
  nand2 gate2134(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2135(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2136(.a(G11), .O(gate439inter7));
  inv1  gate2137(.a(G1162), .O(gate439inter8));
  nand2 gate2138(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2139(.a(s_227), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2140(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2141(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2142(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate799(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate800(.a(gate440inter0), .b(s_36), .O(gate440inter1));
  and2  gate801(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate802(.a(s_36), .O(gate440inter3));
  inv1  gate803(.a(s_37), .O(gate440inter4));
  nand2 gate804(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate805(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate806(.a(G1066), .O(gate440inter7));
  inv1  gate807(.a(G1162), .O(gate440inter8));
  nand2 gate808(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate809(.a(s_37), .b(gate440inter3), .O(gate440inter10));
  nor2  gate810(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate811(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate812(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1065(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1066(.a(gate441inter0), .b(s_74), .O(gate441inter1));
  and2  gate1067(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1068(.a(s_74), .O(gate441inter3));
  inv1  gate1069(.a(s_75), .O(gate441inter4));
  nand2 gate1070(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1071(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1072(.a(G12), .O(gate441inter7));
  inv1  gate1073(.a(G1165), .O(gate441inter8));
  nand2 gate1074(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1075(.a(s_75), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1076(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1077(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1078(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate631(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate632(.a(gate444inter0), .b(s_12), .O(gate444inter1));
  and2  gate633(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate634(.a(s_12), .O(gate444inter3));
  inv1  gate635(.a(s_13), .O(gate444inter4));
  nand2 gate636(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate637(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate638(.a(G1072), .O(gate444inter7));
  inv1  gate639(.a(G1168), .O(gate444inter8));
  nand2 gate640(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate641(.a(s_13), .b(gate444inter3), .O(gate444inter10));
  nor2  gate642(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate643(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate644(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate659(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate660(.a(gate449inter0), .b(s_16), .O(gate449inter1));
  and2  gate661(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate662(.a(s_16), .O(gate449inter3));
  inv1  gate663(.a(s_17), .O(gate449inter4));
  nand2 gate664(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate665(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate666(.a(G16), .O(gate449inter7));
  inv1  gate667(.a(G1177), .O(gate449inter8));
  nand2 gate668(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate669(.a(s_17), .b(gate449inter3), .O(gate449inter10));
  nor2  gate670(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate671(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate672(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate561(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate562(.a(gate450inter0), .b(s_2), .O(gate450inter1));
  and2  gate563(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate564(.a(s_2), .O(gate450inter3));
  inv1  gate565(.a(s_3), .O(gate450inter4));
  nand2 gate566(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate567(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate568(.a(G1081), .O(gate450inter7));
  inv1  gate569(.a(G1177), .O(gate450inter8));
  nand2 gate570(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate571(.a(s_3), .b(gate450inter3), .O(gate450inter10));
  nor2  gate572(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate573(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate574(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1961(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1962(.a(gate451inter0), .b(s_202), .O(gate451inter1));
  and2  gate1963(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1964(.a(s_202), .O(gate451inter3));
  inv1  gate1965(.a(s_203), .O(gate451inter4));
  nand2 gate1966(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1967(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1968(.a(G17), .O(gate451inter7));
  inv1  gate1969(.a(G1180), .O(gate451inter8));
  nand2 gate1970(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1971(.a(s_203), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1972(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1973(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1974(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1457(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1458(.a(gate453inter0), .b(s_130), .O(gate453inter1));
  and2  gate1459(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1460(.a(s_130), .O(gate453inter3));
  inv1  gate1461(.a(s_131), .O(gate453inter4));
  nand2 gate1462(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1463(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1464(.a(G18), .O(gate453inter7));
  inv1  gate1465(.a(G1183), .O(gate453inter8));
  nand2 gate1466(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1467(.a(s_131), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1468(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1469(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1470(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1779(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1780(.a(gate454inter0), .b(s_176), .O(gate454inter1));
  and2  gate1781(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1782(.a(s_176), .O(gate454inter3));
  inv1  gate1783(.a(s_177), .O(gate454inter4));
  nand2 gate1784(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1785(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1786(.a(G1087), .O(gate454inter7));
  inv1  gate1787(.a(G1183), .O(gate454inter8));
  nand2 gate1788(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1789(.a(s_177), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1790(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1791(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1792(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1597(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1598(.a(gate462inter0), .b(s_150), .O(gate462inter1));
  and2  gate1599(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1600(.a(s_150), .O(gate462inter3));
  inv1  gate1601(.a(s_151), .O(gate462inter4));
  nand2 gate1602(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1603(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1604(.a(G1099), .O(gate462inter7));
  inv1  gate1605(.a(G1195), .O(gate462inter8));
  nand2 gate1606(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1607(.a(s_151), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1608(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1609(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1610(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1989(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1990(.a(gate468inter0), .b(s_206), .O(gate468inter1));
  and2  gate1991(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1992(.a(s_206), .O(gate468inter3));
  inv1  gate1993(.a(s_207), .O(gate468inter4));
  nand2 gate1994(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1995(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1996(.a(G1108), .O(gate468inter7));
  inv1  gate1997(.a(G1204), .O(gate468inter8));
  nand2 gate1998(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1999(.a(s_207), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2000(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2001(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2002(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2143(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2144(.a(gate471inter0), .b(s_228), .O(gate471inter1));
  and2  gate2145(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2146(.a(s_228), .O(gate471inter3));
  inv1  gate2147(.a(s_229), .O(gate471inter4));
  nand2 gate2148(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2149(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2150(.a(G27), .O(gate471inter7));
  inv1  gate2151(.a(G1210), .O(gate471inter8));
  nand2 gate2152(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2153(.a(s_229), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2154(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2155(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2156(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1807(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1808(.a(gate475inter0), .b(s_180), .O(gate475inter1));
  and2  gate1809(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1810(.a(s_180), .O(gate475inter3));
  inv1  gate1811(.a(s_181), .O(gate475inter4));
  nand2 gate1812(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1813(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1814(.a(G29), .O(gate475inter7));
  inv1  gate1815(.a(G1216), .O(gate475inter8));
  nand2 gate1816(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1817(.a(s_181), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1818(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1819(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1820(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1303(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1304(.a(gate484inter0), .b(s_108), .O(gate484inter1));
  and2  gate1305(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1306(.a(s_108), .O(gate484inter3));
  inv1  gate1307(.a(s_109), .O(gate484inter4));
  nand2 gate1308(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1309(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1310(.a(G1230), .O(gate484inter7));
  inv1  gate1311(.a(G1231), .O(gate484inter8));
  nand2 gate1312(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1313(.a(s_109), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1314(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1315(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1316(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate603(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate604(.a(gate487inter0), .b(s_8), .O(gate487inter1));
  and2  gate605(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate606(.a(s_8), .O(gate487inter3));
  inv1  gate607(.a(s_9), .O(gate487inter4));
  nand2 gate608(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate609(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate610(.a(G1236), .O(gate487inter7));
  inv1  gate611(.a(G1237), .O(gate487inter8));
  nand2 gate612(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate613(.a(s_9), .b(gate487inter3), .O(gate487inter10));
  nor2  gate614(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate615(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate616(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1947(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1948(.a(gate494inter0), .b(s_200), .O(gate494inter1));
  and2  gate1949(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1950(.a(s_200), .O(gate494inter3));
  inv1  gate1951(.a(s_201), .O(gate494inter4));
  nand2 gate1952(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1953(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1954(.a(G1250), .O(gate494inter7));
  inv1  gate1955(.a(G1251), .O(gate494inter8));
  nand2 gate1956(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1957(.a(s_201), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1958(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1959(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1960(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2171(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2172(.a(gate500inter0), .b(s_232), .O(gate500inter1));
  and2  gate2173(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2174(.a(s_232), .O(gate500inter3));
  inv1  gate2175(.a(s_233), .O(gate500inter4));
  nand2 gate2176(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2177(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2178(.a(G1262), .O(gate500inter7));
  inv1  gate2179(.a(G1263), .O(gate500inter8));
  nand2 gate2180(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2181(.a(s_233), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2182(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2183(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2184(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1527(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1528(.a(gate505inter0), .b(s_140), .O(gate505inter1));
  and2  gate1529(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1530(.a(s_140), .O(gate505inter3));
  inv1  gate1531(.a(s_141), .O(gate505inter4));
  nand2 gate1532(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1533(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1534(.a(G1272), .O(gate505inter7));
  inv1  gate1535(.a(G1273), .O(gate505inter8));
  nand2 gate1536(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1537(.a(s_141), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1538(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1539(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1540(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate2409(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2410(.a(gate506inter0), .b(s_266), .O(gate506inter1));
  and2  gate2411(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2412(.a(s_266), .O(gate506inter3));
  inv1  gate2413(.a(s_267), .O(gate506inter4));
  nand2 gate2414(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2415(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2416(.a(G1274), .O(gate506inter7));
  inv1  gate2417(.a(G1275), .O(gate506inter8));
  nand2 gate2418(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2419(.a(s_267), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2420(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2421(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2422(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule