module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381, s_382, s_383, s_384, s_385, s_386, s_387, s_388, s_389, s_390, s_391;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1457(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1458(.a(gate9inter0), .b(s_130), .O(gate9inter1));
  and2  gate1459(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1460(.a(s_130), .O(gate9inter3));
  inv1  gate1461(.a(s_131), .O(gate9inter4));
  nand2 gate1462(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1463(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1464(.a(G1), .O(gate9inter7));
  inv1  gate1465(.a(G2), .O(gate9inter8));
  nand2 gate1466(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1467(.a(s_131), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1468(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1469(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1470(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1023(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1024(.a(gate10inter0), .b(s_68), .O(gate10inter1));
  and2  gate1025(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1026(.a(s_68), .O(gate10inter3));
  inv1  gate1027(.a(s_69), .O(gate10inter4));
  nand2 gate1028(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1029(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1030(.a(G3), .O(gate10inter7));
  inv1  gate1031(.a(G4), .O(gate10inter8));
  nand2 gate1032(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1033(.a(s_69), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1034(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1035(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1036(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate3179(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate3180(.a(gate13inter0), .b(s_376), .O(gate13inter1));
  and2  gate3181(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate3182(.a(s_376), .O(gate13inter3));
  inv1  gate3183(.a(s_377), .O(gate13inter4));
  nand2 gate3184(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate3185(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate3186(.a(G9), .O(gate13inter7));
  inv1  gate3187(.a(G10), .O(gate13inter8));
  nand2 gate3188(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate3189(.a(s_377), .b(gate13inter3), .O(gate13inter10));
  nor2  gate3190(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate3191(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate3192(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2017(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2018(.a(gate15inter0), .b(s_210), .O(gate15inter1));
  and2  gate2019(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2020(.a(s_210), .O(gate15inter3));
  inv1  gate2021(.a(s_211), .O(gate15inter4));
  nand2 gate2022(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2023(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2024(.a(G13), .O(gate15inter7));
  inv1  gate2025(.a(G14), .O(gate15inter8));
  nand2 gate2026(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2027(.a(s_211), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2028(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2029(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2030(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2353(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2354(.a(gate16inter0), .b(s_258), .O(gate16inter1));
  and2  gate2355(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2356(.a(s_258), .O(gate16inter3));
  inv1  gate2357(.a(s_259), .O(gate16inter4));
  nand2 gate2358(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2359(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2360(.a(G15), .O(gate16inter7));
  inv1  gate2361(.a(G16), .O(gate16inter8));
  nand2 gate2362(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2363(.a(s_259), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2364(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2365(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2366(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1317(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1318(.a(gate17inter0), .b(s_110), .O(gate17inter1));
  and2  gate1319(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1320(.a(s_110), .O(gate17inter3));
  inv1  gate1321(.a(s_111), .O(gate17inter4));
  nand2 gate1322(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1323(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1324(.a(G17), .O(gate17inter7));
  inv1  gate1325(.a(G18), .O(gate17inter8));
  nand2 gate1326(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1327(.a(s_111), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1328(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1329(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1330(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate841(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate842(.a(gate19inter0), .b(s_42), .O(gate19inter1));
  and2  gate843(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate844(.a(s_42), .O(gate19inter3));
  inv1  gate845(.a(s_43), .O(gate19inter4));
  nand2 gate846(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate847(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate848(.a(G21), .O(gate19inter7));
  inv1  gate849(.a(G22), .O(gate19inter8));
  nand2 gate850(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate851(.a(s_43), .b(gate19inter3), .O(gate19inter10));
  nor2  gate852(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate853(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate854(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1835(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1836(.a(gate20inter0), .b(s_184), .O(gate20inter1));
  and2  gate1837(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1838(.a(s_184), .O(gate20inter3));
  inv1  gate1839(.a(s_185), .O(gate20inter4));
  nand2 gate1840(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1841(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1842(.a(G23), .O(gate20inter7));
  inv1  gate1843(.a(G24), .O(gate20inter8));
  nand2 gate1844(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1845(.a(s_185), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1846(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1847(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1848(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1303(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1304(.a(gate22inter0), .b(s_108), .O(gate22inter1));
  and2  gate1305(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1306(.a(s_108), .O(gate22inter3));
  inv1  gate1307(.a(s_109), .O(gate22inter4));
  nand2 gate1308(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1309(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1310(.a(G27), .O(gate22inter7));
  inv1  gate1311(.a(G28), .O(gate22inter8));
  nand2 gate1312(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1313(.a(s_109), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1314(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1315(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1316(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2969(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2970(.a(gate23inter0), .b(s_346), .O(gate23inter1));
  and2  gate2971(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2972(.a(s_346), .O(gate23inter3));
  inv1  gate2973(.a(s_347), .O(gate23inter4));
  nand2 gate2974(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2975(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2976(.a(G29), .O(gate23inter7));
  inv1  gate2977(.a(G30), .O(gate23inter8));
  nand2 gate2978(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2979(.a(s_347), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2980(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2981(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2982(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1695(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1696(.a(gate25inter0), .b(s_164), .O(gate25inter1));
  and2  gate1697(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1698(.a(s_164), .O(gate25inter3));
  inv1  gate1699(.a(s_165), .O(gate25inter4));
  nand2 gate1700(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1701(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1702(.a(G1), .O(gate25inter7));
  inv1  gate1703(.a(G5), .O(gate25inter8));
  nand2 gate1704(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1705(.a(s_165), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1706(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1707(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1708(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2913(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2914(.a(gate28inter0), .b(s_338), .O(gate28inter1));
  and2  gate2915(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2916(.a(s_338), .O(gate28inter3));
  inv1  gate2917(.a(s_339), .O(gate28inter4));
  nand2 gate2918(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2919(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2920(.a(G10), .O(gate28inter7));
  inv1  gate2921(.a(G14), .O(gate28inter8));
  nand2 gate2922(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2923(.a(s_339), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2924(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2925(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2926(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate3151(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate3152(.a(gate30inter0), .b(s_372), .O(gate30inter1));
  and2  gate3153(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate3154(.a(s_372), .O(gate30inter3));
  inv1  gate3155(.a(s_373), .O(gate30inter4));
  nand2 gate3156(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate3157(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate3158(.a(G11), .O(gate30inter7));
  inv1  gate3159(.a(G15), .O(gate30inter8));
  nand2 gate3160(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate3161(.a(s_373), .b(gate30inter3), .O(gate30inter10));
  nor2  gate3162(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate3163(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate3164(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2199(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2200(.a(gate32inter0), .b(s_236), .O(gate32inter1));
  and2  gate2201(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2202(.a(s_236), .O(gate32inter3));
  inv1  gate2203(.a(s_237), .O(gate32inter4));
  nand2 gate2204(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2205(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2206(.a(G12), .O(gate32inter7));
  inv1  gate2207(.a(G16), .O(gate32inter8));
  nand2 gate2208(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2209(.a(s_237), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2210(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2211(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2212(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate561(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate562(.a(gate34inter0), .b(s_2), .O(gate34inter1));
  and2  gate563(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate564(.a(s_2), .O(gate34inter3));
  inv1  gate565(.a(s_3), .O(gate34inter4));
  nand2 gate566(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate567(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate568(.a(G25), .O(gate34inter7));
  inv1  gate569(.a(G29), .O(gate34inter8));
  nand2 gate570(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate571(.a(s_3), .b(gate34inter3), .O(gate34inter10));
  nor2  gate572(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate573(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate574(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1779(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1780(.a(gate35inter0), .b(s_176), .O(gate35inter1));
  and2  gate1781(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1782(.a(s_176), .O(gate35inter3));
  inv1  gate1783(.a(s_177), .O(gate35inter4));
  nand2 gate1784(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1785(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1786(.a(G18), .O(gate35inter7));
  inv1  gate1787(.a(G22), .O(gate35inter8));
  nand2 gate1788(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1789(.a(s_177), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1790(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1791(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1792(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate2815(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2816(.a(gate36inter0), .b(s_324), .O(gate36inter1));
  and2  gate2817(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2818(.a(s_324), .O(gate36inter3));
  inv1  gate2819(.a(s_325), .O(gate36inter4));
  nand2 gate2820(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2821(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2822(.a(G26), .O(gate36inter7));
  inv1  gate2823(.a(G30), .O(gate36inter8));
  nand2 gate2824(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2825(.a(s_325), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2826(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2827(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2828(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1499(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1500(.a(gate38inter0), .b(s_136), .O(gate38inter1));
  and2  gate1501(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1502(.a(s_136), .O(gate38inter3));
  inv1  gate1503(.a(s_137), .O(gate38inter4));
  nand2 gate1504(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1505(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1506(.a(G27), .O(gate38inter7));
  inv1  gate1507(.a(G31), .O(gate38inter8));
  nand2 gate1508(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1509(.a(s_137), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1510(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1511(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1512(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate2787(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2788(.a(gate39inter0), .b(s_320), .O(gate39inter1));
  and2  gate2789(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2790(.a(s_320), .O(gate39inter3));
  inv1  gate2791(.a(s_321), .O(gate39inter4));
  nand2 gate2792(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2793(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2794(.a(G20), .O(gate39inter7));
  inv1  gate2795(.a(G24), .O(gate39inter8));
  nand2 gate2796(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2797(.a(s_321), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2798(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2799(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2800(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2409(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2410(.a(gate43inter0), .b(s_266), .O(gate43inter1));
  and2  gate2411(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2412(.a(s_266), .O(gate43inter3));
  inv1  gate2413(.a(s_267), .O(gate43inter4));
  nand2 gate2414(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2415(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2416(.a(G3), .O(gate43inter7));
  inv1  gate2417(.a(G269), .O(gate43inter8));
  nand2 gate2418(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2419(.a(s_267), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2420(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2421(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2422(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate3221(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate3222(.a(gate46inter0), .b(s_382), .O(gate46inter1));
  and2  gate3223(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate3224(.a(s_382), .O(gate46inter3));
  inv1  gate3225(.a(s_383), .O(gate46inter4));
  nand2 gate3226(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate3227(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate3228(.a(G6), .O(gate46inter7));
  inv1  gate3229(.a(G272), .O(gate46inter8));
  nand2 gate3230(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate3231(.a(s_383), .b(gate46inter3), .O(gate46inter10));
  nor2  gate3232(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate3233(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate3234(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1443(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1444(.a(gate54inter0), .b(s_128), .O(gate54inter1));
  and2  gate1445(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1446(.a(s_128), .O(gate54inter3));
  inv1  gate1447(.a(s_129), .O(gate54inter4));
  nand2 gate1448(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1449(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1450(.a(G14), .O(gate54inter7));
  inv1  gate1451(.a(G284), .O(gate54inter8));
  nand2 gate1452(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1453(.a(s_129), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1454(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1455(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1456(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate631(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate632(.a(gate57inter0), .b(s_12), .O(gate57inter1));
  and2  gate633(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate634(.a(s_12), .O(gate57inter3));
  inv1  gate635(.a(s_13), .O(gate57inter4));
  nand2 gate636(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate637(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate638(.a(G17), .O(gate57inter7));
  inv1  gate639(.a(G290), .O(gate57inter8));
  nand2 gate640(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate641(.a(s_13), .b(gate57inter3), .O(gate57inter10));
  nor2  gate642(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate643(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate644(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate2745(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2746(.a(gate58inter0), .b(s_314), .O(gate58inter1));
  and2  gate2747(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2748(.a(s_314), .O(gate58inter3));
  inv1  gate2749(.a(s_315), .O(gate58inter4));
  nand2 gate2750(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2751(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2752(.a(G18), .O(gate58inter7));
  inv1  gate2753(.a(G290), .O(gate58inter8));
  nand2 gate2754(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2755(.a(s_315), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2756(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2757(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2758(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2689(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2690(.a(gate64inter0), .b(s_306), .O(gate64inter1));
  and2  gate2691(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2692(.a(s_306), .O(gate64inter3));
  inv1  gate2693(.a(s_307), .O(gate64inter4));
  nand2 gate2694(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2695(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2696(.a(G24), .O(gate64inter7));
  inv1  gate2697(.a(G299), .O(gate64inter8));
  nand2 gate2698(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2699(.a(s_307), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2700(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2701(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2702(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1751(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1752(.a(gate67inter0), .b(s_172), .O(gate67inter1));
  and2  gate1753(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1754(.a(s_172), .O(gate67inter3));
  inv1  gate1755(.a(s_173), .O(gate67inter4));
  nand2 gate1756(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1757(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1758(.a(G27), .O(gate67inter7));
  inv1  gate1759(.a(G305), .O(gate67inter8));
  nand2 gate1760(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1761(.a(s_173), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1762(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1763(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1764(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate3249(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate3250(.a(gate68inter0), .b(s_386), .O(gate68inter1));
  and2  gate3251(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate3252(.a(s_386), .O(gate68inter3));
  inv1  gate3253(.a(s_387), .O(gate68inter4));
  nand2 gate3254(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate3255(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate3256(.a(G28), .O(gate68inter7));
  inv1  gate3257(.a(G305), .O(gate68inter8));
  nand2 gate3258(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate3259(.a(s_387), .b(gate68inter3), .O(gate68inter10));
  nor2  gate3260(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate3261(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate3262(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate2731(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2732(.a(gate69inter0), .b(s_312), .O(gate69inter1));
  and2  gate2733(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2734(.a(s_312), .O(gate69inter3));
  inv1  gate2735(.a(s_313), .O(gate69inter4));
  nand2 gate2736(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2737(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2738(.a(G29), .O(gate69inter7));
  inv1  gate2739(.a(G308), .O(gate69inter8));
  nand2 gate2740(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2741(.a(s_313), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2742(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2743(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2744(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate3039(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate3040(.a(gate70inter0), .b(s_356), .O(gate70inter1));
  and2  gate3041(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate3042(.a(s_356), .O(gate70inter3));
  inv1  gate3043(.a(s_357), .O(gate70inter4));
  nand2 gate3044(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate3045(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate3046(.a(G30), .O(gate70inter7));
  inv1  gate3047(.a(G308), .O(gate70inter8));
  nand2 gate3048(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate3049(.a(s_357), .b(gate70inter3), .O(gate70inter10));
  nor2  gate3050(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate3051(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate3052(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2675(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2676(.a(gate74inter0), .b(s_304), .O(gate74inter1));
  and2  gate2677(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2678(.a(s_304), .O(gate74inter3));
  inv1  gate2679(.a(s_305), .O(gate74inter4));
  nand2 gate2680(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2681(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2682(.a(G5), .O(gate74inter7));
  inv1  gate2683(.a(G314), .O(gate74inter8));
  nand2 gate2684(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2685(.a(s_305), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2686(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2687(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2688(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2059(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2060(.a(gate76inter0), .b(s_216), .O(gate76inter1));
  and2  gate2061(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2062(.a(s_216), .O(gate76inter3));
  inv1  gate2063(.a(s_217), .O(gate76inter4));
  nand2 gate2064(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2065(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2066(.a(G13), .O(gate76inter7));
  inv1  gate2067(.a(G317), .O(gate76inter8));
  nand2 gate2068(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2069(.a(s_217), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2070(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2071(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2072(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1625(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1626(.a(gate77inter0), .b(s_154), .O(gate77inter1));
  and2  gate1627(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1628(.a(s_154), .O(gate77inter3));
  inv1  gate1629(.a(s_155), .O(gate77inter4));
  nand2 gate1630(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1631(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1632(.a(G2), .O(gate77inter7));
  inv1  gate1633(.a(G320), .O(gate77inter8));
  nand2 gate1634(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1635(.a(s_155), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1636(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1637(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1638(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate939(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate940(.a(gate78inter0), .b(s_56), .O(gate78inter1));
  and2  gate941(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate942(.a(s_56), .O(gate78inter3));
  inv1  gate943(.a(s_57), .O(gate78inter4));
  nand2 gate944(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate945(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate946(.a(G6), .O(gate78inter7));
  inv1  gate947(.a(G320), .O(gate78inter8));
  nand2 gate948(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate949(.a(s_57), .b(gate78inter3), .O(gate78inter10));
  nor2  gate950(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate951(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate952(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2437(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2438(.a(gate80inter0), .b(s_270), .O(gate80inter1));
  and2  gate2439(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2440(.a(s_270), .O(gate80inter3));
  inv1  gate2441(.a(s_271), .O(gate80inter4));
  nand2 gate2442(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2443(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2444(.a(G14), .O(gate80inter7));
  inv1  gate2445(.a(G323), .O(gate80inter8));
  nand2 gate2446(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2447(.a(s_271), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2448(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2449(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2450(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate715(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate716(.a(gate82inter0), .b(s_24), .O(gate82inter1));
  and2  gate717(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate718(.a(s_24), .O(gate82inter3));
  inv1  gate719(.a(s_25), .O(gate82inter4));
  nand2 gate720(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate721(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate722(.a(G7), .O(gate82inter7));
  inv1  gate723(.a(G326), .O(gate82inter8));
  nand2 gate724(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate725(.a(s_25), .b(gate82inter3), .O(gate82inter10));
  nor2  gate726(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate727(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate728(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1807(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1808(.a(gate88inter0), .b(s_180), .O(gate88inter1));
  and2  gate1809(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1810(.a(s_180), .O(gate88inter3));
  inv1  gate1811(.a(s_181), .O(gate88inter4));
  nand2 gate1812(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1813(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1814(.a(G16), .O(gate88inter7));
  inv1  gate1815(.a(G335), .O(gate88inter8));
  nand2 gate1816(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1817(.a(s_181), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1818(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1819(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1820(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2423(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2424(.a(gate90inter0), .b(s_268), .O(gate90inter1));
  and2  gate2425(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2426(.a(s_268), .O(gate90inter3));
  inv1  gate2427(.a(s_269), .O(gate90inter4));
  nand2 gate2428(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2429(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2430(.a(G21), .O(gate90inter7));
  inv1  gate2431(.a(G338), .O(gate90inter8));
  nand2 gate2432(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2433(.a(s_269), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2434(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2435(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2436(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1471(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1472(.a(gate91inter0), .b(s_132), .O(gate91inter1));
  and2  gate1473(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1474(.a(s_132), .O(gate91inter3));
  inv1  gate1475(.a(s_133), .O(gate91inter4));
  nand2 gate1476(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1477(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1478(.a(G25), .O(gate91inter7));
  inv1  gate1479(.a(G341), .O(gate91inter8));
  nand2 gate1480(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1481(.a(s_133), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1482(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1483(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1484(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1079(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1080(.a(gate99inter0), .b(s_76), .O(gate99inter1));
  and2  gate1081(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1082(.a(s_76), .O(gate99inter3));
  inv1  gate1083(.a(s_77), .O(gate99inter4));
  nand2 gate1084(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1085(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1086(.a(G27), .O(gate99inter7));
  inv1  gate1087(.a(G353), .O(gate99inter8));
  nand2 gate1088(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1089(.a(s_77), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1090(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1091(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1092(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate2227(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2228(.a(gate100inter0), .b(s_240), .O(gate100inter1));
  and2  gate2229(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2230(.a(s_240), .O(gate100inter3));
  inv1  gate2231(.a(s_241), .O(gate100inter4));
  nand2 gate2232(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2233(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2234(.a(G31), .O(gate100inter7));
  inv1  gate2235(.a(G353), .O(gate100inter8));
  nand2 gate2236(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2237(.a(s_241), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2238(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2239(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2240(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate743(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate744(.a(gate101inter0), .b(s_28), .O(gate101inter1));
  and2  gate745(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate746(.a(s_28), .O(gate101inter3));
  inv1  gate747(.a(s_29), .O(gate101inter4));
  nand2 gate748(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate749(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate750(.a(G20), .O(gate101inter7));
  inv1  gate751(.a(G356), .O(gate101inter8));
  nand2 gate752(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate753(.a(s_29), .b(gate101inter3), .O(gate101inter10));
  nor2  gate754(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate755(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate756(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2941(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2942(.a(gate102inter0), .b(s_342), .O(gate102inter1));
  and2  gate2943(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2944(.a(s_342), .O(gate102inter3));
  inv1  gate2945(.a(s_343), .O(gate102inter4));
  nand2 gate2946(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2947(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2948(.a(G24), .O(gate102inter7));
  inv1  gate2949(.a(G356), .O(gate102inter8));
  nand2 gate2950(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2951(.a(s_343), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2952(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2953(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2954(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1205(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1206(.a(gate103inter0), .b(s_94), .O(gate103inter1));
  and2  gate1207(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1208(.a(s_94), .O(gate103inter3));
  inv1  gate1209(.a(s_95), .O(gate103inter4));
  nand2 gate1210(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1211(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1212(.a(G28), .O(gate103inter7));
  inv1  gate1213(.a(G359), .O(gate103inter8));
  nand2 gate1214(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1215(.a(s_95), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1216(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1217(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1218(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1429(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1430(.a(gate105inter0), .b(s_126), .O(gate105inter1));
  and2  gate1431(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1432(.a(s_126), .O(gate105inter3));
  inv1  gate1433(.a(s_127), .O(gate105inter4));
  nand2 gate1434(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1435(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1436(.a(G362), .O(gate105inter7));
  inv1  gate1437(.a(G363), .O(gate105inter8));
  nand2 gate1438(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1439(.a(s_127), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1440(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1441(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1442(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1723(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1724(.a(gate108inter0), .b(s_168), .O(gate108inter1));
  and2  gate1725(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1726(.a(s_168), .O(gate108inter3));
  inv1  gate1727(.a(s_169), .O(gate108inter4));
  nand2 gate1728(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1729(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1730(.a(G368), .O(gate108inter7));
  inv1  gate1731(.a(G369), .O(gate108inter8));
  nand2 gate1732(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1733(.a(s_169), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1734(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1735(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1736(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate2213(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2214(.a(gate109inter0), .b(s_238), .O(gate109inter1));
  and2  gate2215(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2216(.a(s_238), .O(gate109inter3));
  inv1  gate2217(.a(s_239), .O(gate109inter4));
  nand2 gate2218(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2219(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2220(.a(G370), .O(gate109inter7));
  inv1  gate2221(.a(G371), .O(gate109inter8));
  nand2 gate2222(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2223(.a(s_239), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2224(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2225(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2226(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1009(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1010(.a(gate112inter0), .b(s_66), .O(gate112inter1));
  and2  gate1011(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1012(.a(s_66), .O(gate112inter3));
  inv1  gate1013(.a(s_67), .O(gate112inter4));
  nand2 gate1014(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1015(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1016(.a(G376), .O(gate112inter7));
  inv1  gate1017(.a(G377), .O(gate112inter8));
  nand2 gate1018(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1019(.a(s_67), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1020(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1021(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1022(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate2283(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2284(.a(gate113inter0), .b(s_248), .O(gate113inter1));
  and2  gate2285(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2286(.a(s_248), .O(gate113inter3));
  inv1  gate2287(.a(s_249), .O(gate113inter4));
  nand2 gate2288(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2289(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2290(.a(G378), .O(gate113inter7));
  inv1  gate2291(.a(G379), .O(gate113inter8));
  nand2 gate2292(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2293(.a(s_249), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2294(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2295(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2296(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate1583(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1584(.a(gate114inter0), .b(s_148), .O(gate114inter1));
  and2  gate1585(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1586(.a(s_148), .O(gate114inter3));
  inv1  gate1587(.a(s_149), .O(gate114inter4));
  nand2 gate1588(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1589(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1590(.a(G380), .O(gate114inter7));
  inv1  gate1591(.a(G381), .O(gate114inter8));
  nand2 gate1592(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1593(.a(s_149), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1594(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1595(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1596(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate2843(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2844(.a(gate115inter0), .b(s_328), .O(gate115inter1));
  and2  gate2845(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2846(.a(s_328), .O(gate115inter3));
  inv1  gate2847(.a(s_329), .O(gate115inter4));
  nand2 gate2848(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2849(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2850(.a(G382), .O(gate115inter7));
  inv1  gate2851(.a(G383), .O(gate115inter8));
  nand2 gate2852(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2853(.a(s_329), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2854(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2855(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2856(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate2311(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2312(.a(gate116inter0), .b(s_252), .O(gate116inter1));
  and2  gate2313(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2314(.a(s_252), .O(gate116inter3));
  inv1  gate2315(.a(s_253), .O(gate116inter4));
  nand2 gate2316(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2317(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2318(.a(G384), .O(gate116inter7));
  inv1  gate2319(.a(G385), .O(gate116inter8));
  nand2 gate2320(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2321(.a(s_253), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2322(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2323(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2324(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1737(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1738(.a(gate117inter0), .b(s_170), .O(gate117inter1));
  and2  gate1739(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1740(.a(s_170), .O(gate117inter3));
  inv1  gate1741(.a(s_171), .O(gate117inter4));
  nand2 gate1742(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1743(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1744(.a(G386), .O(gate117inter7));
  inv1  gate1745(.a(G387), .O(gate117inter8));
  nand2 gate1746(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1747(.a(s_171), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1748(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1749(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1750(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1527(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1528(.a(gate119inter0), .b(s_140), .O(gate119inter1));
  and2  gate1529(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1530(.a(s_140), .O(gate119inter3));
  inv1  gate1531(.a(s_141), .O(gate119inter4));
  nand2 gate1532(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1533(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1534(.a(G390), .O(gate119inter7));
  inv1  gate1535(.a(G391), .O(gate119inter8));
  nand2 gate1536(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1537(.a(s_141), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1538(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1539(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1540(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1821(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1822(.a(gate130inter0), .b(s_182), .O(gate130inter1));
  and2  gate1823(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1824(.a(s_182), .O(gate130inter3));
  inv1  gate1825(.a(s_183), .O(gate130inter4));
  nand2 gate1826(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1827(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1828(.a(G412), .O(gate130inter7));
  inv1  gate1829(.a(G413), .O(gate130inter8));
  nand2 gate1830(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1831(.a(s_183), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1832(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1833(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1834(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate3011(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate3012(.a(gate132inter0), .b(s_352), .O(gate132inter1));
  and2  gate3013(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate3014(.a(s_352), .O(gate132inter3));
  inv1  gate3015(.a(s_353), .O(gate132inter4));
  nand2 gate3016(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate3017(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate3018(.a(G416), .O(gate132inter7));
  inv1  gate3019(.a(G417), .O(gate132inter8));
  nand2 gate3020(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate3021(.a(s_353), .b(gate132inter3), .O(gate132inter10));
  nor2  gate3022(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate3023(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate3024(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1667(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1668(.a(gate134inter0), .b(s_160), .O(gate134inter1));
  and2  gate1669(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1670(.a(s_160), .O(gate134inter3));
  inv1  gate1671(.a(s_161), .O(gate134inter4));
  nand2 gate1672(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1673(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1674(.a(G420), .O(gate134inter7));
  inv1  gate1675(.a(G421), .O(gate134inter8));
  nand2 gate1676(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1677(.a(s_161), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1678(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1679(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1680(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2591(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2592(.a(gate135inter0), .b(s_292), .O(gate135inter1));
  and2  gate2593(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2594(.a(s_292), .O(gate135inter3));
  inv1  gate2595(.a(s_293), .O(gate135inter4));
  nand2 gate2596(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2597(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2598(.a(G422), .O(gate135inter7));
  inv1  gate2599(.a(G423), .O(gate135inter8));
  nand2 gate2600(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2601(.a(s_293), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2602(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2603(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2604(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate2619(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2620(.a(gate136inter0), .b(s_296), .O(gate136inter1));
  and2  gate2621(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2622(.a(s_296), .O(gate136inter3));
  inv1  gate2623(.a(s_297), .O(gate136inter4));
  nand2 gate2624(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2625(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2626(.a(G424), .O(gate136inter7));
  inv1  gate2627(.a(G425), .O(gate136inter8));
  nand2 gate2628(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2629(.a(s_297), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2630(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2631(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2632(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate3053(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate3054(.a(gate138inter0), .b(s_358), .O(gate138inter1));
  and2  gate3055(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate3056(.a(s_358), .O(gate138inter3));
  inv1  gate3057(.a(s_359), .O(gate138inter4));
  nand2 gate3058(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate3059(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate3060(.a(G432), .O(gate138inter7));
  inv1  gate3061(.a(G435), .O(gate138inter8));
  nand2 gate3062(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate3063(.a(s_359), .b(gate138inter3), .O(gate138inter10));
  nor2  gate3064(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate3065(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate3066(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate799(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate800(.a(gate139inter0), .b(s_36), .O(gate139inter1));
  and2  gate801(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate802(.a(s_36), .O(gate139inter3));
  inv1  gate803(.a(s_37), .O(gate139inter4));
  nand2 gate804(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate805(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate806(.a(G438), .O(gate139inter7));
  inv1  gate807(.a(G441), .O(gate139inter8));
  nand2 gate808(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate809(.a(s_37), .b(gate139inter3), .O(gate139inter10));
  nor2  gate810(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate811(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate812(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate2143(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2144(.a(gate140inter0), .b(s_228), .O(gate140inter1));
  and2  gate2145(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2146(.a(s_228), .O(gate140inter3));
  inv1  gate2147(.a(s_229), .O(gate140inter4));
  nand2 gate2148(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2149(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2150(.a(G444), .O(gate140inter7));
  inv1  gate2151(.a(G447), .O(gate140inter8));
  nand2 gate2152(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2153(.a(s_229), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2154(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2155(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2156(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1275(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1276(.a(gate142inter0), .b(s_104), .O(gate142inter1));
  and2  gate1277(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1278(.a(s_104), .O(gate142inter3));
  inv1  gate1279(.a(s_105), .O(gate142inter4));
  nand2 gate1280(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1281(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1282(.a(G456), .O(gate142inter7));
  inv1  gate1283(.a(G459), .O(gate142inter8));
  nand2 gate1284(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1285(.a(s_105), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1286(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1287(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1288(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1177(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1178(.a(gate143inter0), .b(s_90), .O(gate143inter1));
  and2  gate1179(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1180(.a(s_90), .O(gate143inter3));
  inv1  gate1181(.a(s_91), .O(gate143inter4));
  nand2 gate1182(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1183(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1184(.a(G462), .O(gate143inter7));
  inv1  gate1185(.a(G465), .O(gate143inter8));
  nand2 gate1186(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1187(.a(s_91), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1188(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1189(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1190(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate575(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate576(.a(gate145inter0), .b(s_4), .O(gate145inter1));
  and2  gate577(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate578(.a(s_4), .O(gate145inter3));
  inv1  gate579(.a(s_5), .O(gate145inter4));
  nand2 gate580(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate581(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate582(.a(G474), .O(gate145inter7));
  inv1  gate583(.a(G477), .O(gate145inter8));
  nand2 gate584(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate585(.a(s_5), .b(gate145inter3), .O(gate145inter10));
  nor2  gate586(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate587(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate588(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1121(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1122(.a(gate146inter0), .b(s_82), .O(gate146inter1));
  and2  gate1123(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1124(.a(s_82), .O(gate146inter3));
  inv1  gate1125(.a(s_83), .O(gate146inter4));
  nand2 gate1126(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1127(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1128(.a(G480), .O(gate146inter7));
  inv1  gate1129(.a(G483), .O(gate146inter8));
  nand2 gate1130(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1131(.a(s_83), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1132(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1133(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1134(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1289(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1290(.a(gate147inter0), .b(s_106), .O(gate147inter1));
  and2  gate1291(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1292(.a(s_106), .O(gate147inter3));
  inv1  gate1293(.a(s_107), .O(gate147inter4));
  nand2 gate1294(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1295(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1296(.a(G486), .O(gate147inter7));
  inv1  gate1297(.a(G489), .O(gate147inter8));
  nand2 gate1298(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1299(.a(s_107), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1300(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1301(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1302(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1331(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1332(.a(gate151inter0), .b(s_112), .O(gate151inter1));
  and2  gate1333(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1334(.a(s_112), .O(gate151inter3));
  inv1  gate1335(.a(s_113), .O(gate151inter4));
  nand2 gate1336(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1337(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1338(.a(G510), .O(gate151inter7));
  inv1  gate1339(.a(G513), .O(gate151inter8));
  nand2 gate1340(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1341(.a(s_113), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1342(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1343(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1344(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate729(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate730(.a(gate152inter0), .b(s_26), .O(gate152inter1));
  and2  gate731(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate732(.a(s_26), .O(gate152inter3));
  inv1  gate733(.a(s_27), .O(gate152inter4));
  nand2 gate734(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate735(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate736(.a(G516), .O(gate152inter7));
  inv1  gate737(.a(G519), .O(gate152inter8));
  nand2 gate738(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate739(.a(s_27), .b(gate152inter3), .O(gate152inter10));
  nor2  gate740(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate741(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate742(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2521(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2522(.a(gate157inter0), .b(s_282), .O(gate157inter1));
  and2  gate2523(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2524(.a(s_282), .O(gate157inter3));
  inv1  gate2525(.a(s_283), .O(gate157inter4));
  nand2 gate2526(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2527(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2528(.a(G438), .O(gate157inter7));
  inv1  gate2529(.a(G528), .O(gate157inter8));
  nand2 gate2530(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2531(.a(s_283), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2532(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2533(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2534(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1359(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1360(.a(gate158inter0), .b(s_116), .O(gate158inter1));
  and2  gate1361(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1362(.a(s_116), .O(gate158inter3));
  inv1  gate1363(.a(s_117), .O(gate158inter4));
  nand2 gate1364(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1365(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1366(.a(G441), .O(gate158inter7));
  inv1  gate1367(.a(G528), .O(gate158inter8));
  nand2 gate1368(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1369(.a(s_117), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1370(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1371(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1372(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2759(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2760(.a(gate161inter0), .b(s_316), .O(gate161inter1));
  and2  gate2761(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2762(.a(s_316), .O(gate161inter3));
  inv1  gate2763(.a(s_317), .O(gate161inter4));
  nand2 gate2764(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2765(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2766(.a(G450), .O(gate161inter7));
  inv1  gate2767(.a(G534), .O(gate161inter8));
  nand2 gate2768(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2769(.a(s_317), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2770(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2771(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2772(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate589(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate590(.a(gate163inter0), .b(s_6), .O(gate163inter1));
  and2  gate591(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate592(.a(s_6), .O(gate163inter3));
  inv1  gate593(.a(s_7), .O(gate163inter4));
  nand2 gate594(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate595(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate596(.a(G456), .O(gate163inter7));
  inv1  gate597(.a(G537), .O(gate163inter8));
  nand2 gate598(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate599(.a(s_7), .b(gate163inter3), .O(gate163inter10));
  nor2  gate600(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate601(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate602(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1877(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1878(.a(gate165inter0), .b(s_190), .O(gate165inter1));
  and2  gate1879(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1880(.a(s_190), .O(gate165inter3));
  inv1  gate1881(.a(s_191), .O(gate165inter4));
  nand2 gate1882(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1883(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1884(.a(G462), .O(gate165inter7));
  inv1  gate1885(.a(G540), .O(gate165inter8));
  nand2 gate1886(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1887(.a(s_191), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1888(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1889(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1890(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate953(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate954(.a(gate167inter0), .b(s_58), .O(gate167inter1));
  and2  gate955(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate956(.a(s_58), .O(gate167inter3));
  inv1  gate957(.a(s_59), .O(gate167inter4));
  nand2 gate958(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate959(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate960(.a(G468), .O(gate167inter7));
  inv1  gate961(.a(G543), .O(gate167inter8));
  nand2 gate962(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate963(.a(s_59), .b(gate167inter3), .O(gate167inter10));
  nor2  gate964(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate965(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate966(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate3123(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate3124(.a(gate170inter0), .b(s_368), .O(gate170inter1));
  and2  gate3125(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate3126(.a(s_368), .O(gate170inter3));
  inv1  gate3127(.a(s_369), .O(gate170inter4));
  nand2 gate3128(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate3129(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate3130(.a(G477), .O(gate170inter7));
  inv1  gate3131(.a(G546), .O(gate170inter8));
  nand2 gate3132(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate3133(.a(s_369), .b(gate170inter3), .O(gate170inter10));
  nor2  gate3134(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate3135(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate3136(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2157(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2158(.a(gate175inter0), .b(s_230), .O(gate175inter1));
  and2  gate2159(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2160(.a(s_230), .O(gate175inter3));
  inv1  gate2161(.a(s_231), .O(gate175inter4));
  nand2 gate2162(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2163(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2164(.a(G492), .O(gate175inter7));
  inv1  gate2165(.a(G555), .O(gate175inter8));
  nand2 gate2166(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2167(.a(s_231), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2168(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2169(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2170(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate2507(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2508(.a(gate176inter0), .b(s_280), .O(gate176inter1));
  and2  gate2509(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2510(.a(s_280), .O(gate176inter3));
  inv1  gate2511(.a(s_281), .O(gate176inter4));
  nand2 gate2512(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2513(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2514(.a(G495), .O(gate176inter7));
  inv1  gate2515(.a(G555), .O(gate176inter8));
  nand2 gate2516(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2517(.a(s_281), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2518(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2519(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2520(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate2367(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2368(.a(gate178inter0), .b(s_260), .O(gate178inter1));
  and2  gate2369(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2370(.a(s_260), .O(gate178inter3));
  inv1  gate2371(.a(s_261), .O(gate178inter4));
  nand2 gate2372(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2373(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2374(.a(G501), .O(gate178inter7));
  inv1  gate2375(.a(G558), .O(gate178inter8));
  nand2 gate2376(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2377(.a(s_261), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2378(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2379(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2380(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate3207(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate3208(.a(gate181inter0), .b(s_380), .O(gate181inter1));
  and2  gate3209(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate3210(.a(s_380), .O(gate181inter3));
  inv1  gate3211(.a(s_381), .O(gate181inter4));
  nand2 gate3212(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate3213(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate3214(.a(G510), .O(gate181inter7));
  inv1  gate3215(.a(G564), .O(gate181inter8));
  nand2 gate3216(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate3217(.a(s_381), .b(gate181inter3), .O(gate181inter10));
  nor2  gate3218(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate3219(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate3220(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate3067(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate3068(.a(gate182inter0), .b(s_360), .O(gate182inter1));
  and2  gate3069(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate3070(.a(s_360), .O(gate182inter3));
  inv1  gate3071(.a(s_361), .O(gate182inter4));
  nand2 gate3072(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate3073(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate3074(.a(G513), .O(gate182inter7));
  inv1  gate3075(.a(G564), .O(gate182inter8));
  nand2 gate3076(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate3077(.a(s_361), .b(gate182inter3), .O(gate182inter10));
  nor2  gate3078(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate3079(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate3080(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1247(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1248(.a(gate183inter0), .b(s_100), .O(gate183inter1));
  and2  gate1249(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1250(.a(s_100), .O(gate183inter3));
  inv1  gate1251(.a(s_101), .O(gate183inter4));
  nand2 gate1252(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1253(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1254(.a(G516), .O(gate183inter7));
  inv1  gate1255(.a(G567), .O(gate183inter8));
  nand2 gate1256(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1257(.a(s_101), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1258(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1259(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1260(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1541(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1542(.a(gate186inter0), .b(s_142), .O(gate186inter1));
  and2  gate1543(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1544(.a(s_142), .O(gate186inter3));
  inv1  gate1545(.a(s_143), .O(gate186inter4));
  nand2 gate1546(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1547(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1548(.a(G572), .O(gate186inter7));
  inv1  gate1549(.a(G573), .O(gate186inter8));
  nand2 gate1550(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1551(.a(s_143), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1552(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1553(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1554(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate2563(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2564(.a(gate187inter0), .b(s_288), .O(gate187inter1));
  and2  gate2565(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2566(.a(s_288), .O(gate187inter3));
  inv1  gate2567(.a(s_289), .O(gate187inter4));
  nand2 gate2568(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2569(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2570(.a(G574), .O(gate187inter7));
  inv1  gate2571(.a(G575), .O(gate187inter8));
  nand2 gate2572(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2573(.a(s_289), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2574(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2575(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2576(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate603(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate604(.a(gate188inter0), .b(s_8), .O(gate188inter1));
  and2  gate605(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate606(.a(s_8), .O(gate188inter3));
  inv1  gate607(.a(s_9), .O(gate188inter4));
  nand2 gate608(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate609(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate610(.a(G576), .O(gate188inter7));
  inv1  gate611(.a(G577), .O(gate188inter8));
  nand2 gate612(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate613(.a(s_9), .b(gate188inter3), .O(gate188inter10));
  nor2  gate614(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate615(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate616(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate645(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate646(.a(gate189inter0), .b(s_14), .O(gate189inter1));
  and2  gate647(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate648(.a(s_14), .O(gate189inter3));
  inv1  gate649(.a(s_15), .O(gate189inter4));
  nand2 gate650(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate651(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate652(.a(G578), .O(gate189inter7));
  inv1  gate653(.a(G579), .O(gate189inter8));
  nand2 gate654(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate655(.a(s_15), .b(gate189inter3), .O(gate189inter10));
  nor2  gate656(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate657(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate658(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1933(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1934(.a(gate196inter0), .b(s_198), .O(gate196inter1));
  and2  gate1935(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1936(.a(s_198), .O(gate196inter3));
  inv1  gate1937(.a(s_199), .O(gate196inter4));
  nand2 gate1938(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1939(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1940(.a(G592), .O(gate196inter7));
  inv1  gate1941(.a(G593), .O(gate196inter8));
  nand2 gate1942(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1943(.a(s_199), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1944(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1945(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1946(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1975(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1976(.a(gate197inter0), .b(s_204), .O(gate197inter1));
  and2  gate1977(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1978(.a(s_204), .O(gate197inter3));
  inv1  gate1979(.a(s_205), .O(gate197inter4));
  nand2 gate1980(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1981(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1982(.a(G594), .O(gate197inter7));
  inv1  gate1983(.a(G595), .O(gate197inter8));
  nand2 gate1984(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1985(.a(s_205), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1986(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1987(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1988(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2087(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2088(.a(gate201inter0), .b(s_220), .O(gate201inter1));
  and2  gate2089(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2090(.a(s_220), .O(gate201inter3));
  inv1  gate2091(.a(s_221), .O(gate201inter4));
  nand2 gate2092(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2093(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2094(.a(G602), .O(gate201inter7));
  inv1  gate2095(.a(G607), .O(gate201inter8));
  nand2 gate2096(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2097(.a(s_221), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2098(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2099(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2100(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1261(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1262(.a(gate202inter0), .b(s_102), .O(gate202inter1));
  and2  gate1263(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1264(.a(s_102), .O(gate202inter3));
  inv1  gate1265(.a(s_103), .O(gate202inter4));
  nand2 gate1266(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1267(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1268(.a(G612), .O(gate202inter7));
  inv1  gate1269(.a(G617), .O(gate202inter8));
  nand2 gate1270(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1271(.a(s_103), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1272(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1273(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1274(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate2269(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2270(.a(gate203inter0), .b(s_246), .O(gate203inter1));
  and2  gate2271(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2272(.a(s_246), .O(gate203inter3));
  inv1  gate2273(.a(s_247), .O(gate203inter4));
  nand2 gate2274(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2275(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2276(.a(G602), .O(gate203inter7));
  inv1  gate2277(.a(G612), .O(gate203inter8));
  nand2 gate2278(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2279(.a(s_247), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2280(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2281(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2282(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate3235(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate3236(.a(gate212inter0), .b(s_384), .O(gate212inter1));
  and2  gate3237(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate3238(.a(s_384), .O(gate212inter3));
  inv1  gate3239(.a(s_385), .O(gate212inter4));
  nand2 gate3240(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate3241(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate3242(.a(G617), .O(gate212inter7));
  inv1  gate3243(.a(G669), .O(gate212inter8));
  nand2 gate3244(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate3245(.a(s_385), .b(gate212inter3), .O(gate212inter10));
  nor2  gate3246(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate3247(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate3248(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate2255(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2256(.a(gate213inter0), .b(s_244), .O(gate213inter1));
  and2  gate2257(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2258(.a(s_244), .O(gate213inter3));
  inv1  gate2259(.a(s_245), .O(gate213inter4));
  nand2 gate2260(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2261(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2262(.a(G602), .O(gate213inter7));
  inv1  gate2263(.a(G672), .O(gate213inter8));
  nand2 gate2264(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2265(.a(s_245), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2266(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2267(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2268(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate785(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate786(.a(gate215inter0), .b(s_34), .O(gate215inter1));
  and2  gate787(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate788(.a(s_34), .O(gate215inter3));
  inv1  gate789(.a(s_35), .O(gate215inter4));
  nand2 gate790(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate791(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate792(.a(G607), .O(gate215inter7));
  inv1  gate793(.a(G675), .O(gate215inter8));
  nand2 gate794(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate795(.a(s_35), .b(gate215inter3), .O(gate215inter10));
  nor2  gate796(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate797(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate798(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate3277(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate3278(.a(gate219inter0), .b(s_390), .O(gate219inter1));
  and2  gate3279(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate3280(.a(s_390), .O(gate219inter3));
  inv1  gate3281(.a(s_391), .O(gate219inter4));
  nand2 gate3282(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate3283(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate3284(.a(G632), .O(gate219inter7));
  inv1  gate3285(.a(G681), .O(gate219inter8));
  nand2 gate3286(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate3287(.a(s_391), .b(gate219inter3), .O(gate219inter10));
  nor2  gate3288(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate3289(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate3290(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate2395(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate2396(.a(gate222inter0), .b(s_264), .O(gate222inter1));
  and2  gate2397(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate2398(.a(s_264), .O(gate222inter3));
  inv1  gate2399(.a(s_265), .O(gate222inter4));
  nand2 gate2400(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate2401(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate2402(.a(G632), .O(gate222inter7));
  inv1  gate2403(.a(G684), .O(gate222inter8));
  nand2 gate2404(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate2405(.a(s_265), .b(gate222inter3), .O(gate222inter10));
  nor2  gate2406(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate2407(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate2408(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate2801(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate2802(.a(gate226inter0), .b(s_322), .O(gate226inter1));
  and2  gate2803(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate2804(.a(s_322), .O(gate226inter3));
  inv1  gate2805(.a(s_323), .O(gate226inter4));
  nand2 gate2806(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate2807(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate2808(.a(G692), .O(gate226inter7));
  inv1  gate2809(.a(G693), .O(gate226inter8));
  nand2 gate2810(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate2811(.a(s_323), .b(gate226inter3), .O(gate226inter10));
  nor2  gate2812(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate2813(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate2814(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1597(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1598(.a(gate227inter0), .b(s_150), .O(gate227inter1));
  and2  gate1599(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1600(.a(s_150), .O(gate227inter3));
  inv1  gate1601(.a(s_151), .O(gate227inter4));
  nand2 gate1602(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1603(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1604(.a(G694), .O(gate227inter7));
  inv1  gate1605(.a(G695), .O(gate227inter8));
  nand2 gate1606(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1607(.a(s_151), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1608(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1609(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1610(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate995(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate996(.a(gate230inter0), .b(s_64), .O(gate230inter1));
  and2  gate997(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate998(.a(s_64), .O(gate230inter3));
  inv1  gate999(.a(s_65), .O(gate230inter4));
  nand2 gate1000(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1001(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1002(.a(G700), .O(gate230inter7));
  inv1  gate1003(.a(G701), .O(gate230inter8));
  nand2 gate1004(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1005(.a(s_65), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1006(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1007(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1008(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2927(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2928(.a(gate232inter0), .b(s_340), .O(gate232inter1));
  and2  gate2929(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2930(.a(s_340), .O(gate232inter3));
  inv1  gate2931(.a(s_341), .O(gate232inter4));
  nand2 gate2932(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2933(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2934(.a(G704), .O(gate232inter7));
  inv1  gate2935(.a(G705), .O(gate232inter8));
  nand2 gate2936(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2937(.a(s_341), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2938(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2939(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2940(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate897(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate898(.a(gate233inter0), .b(s_50), .O(gate233inter1));
  and2  gate899(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate900(.a(s_50), .O(gate233inter3));
  inv1  gate901(.a(s_51), .O(gate233inter4));
  nand2 gate902(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate903(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate904(.a(G242), .O(gate233inter7));
  inv1  gate905(.a(G718), .O(gate233inter8));
  nand2 gate906(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate907(.a(s_51), .b(gate233inter3), .O(gate233inter10));
  nor2  gate908(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate909(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate910(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1051(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1052(.a(gate234inter0), .b(s_72), .O(gate234inter1));
  and2  gate1053(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1054(.a(s_72), .O(gate234inter3));
  inv1  gate1055(.a(s_73), .O(gate234inter4));
  nand2 gate1056(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1057(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1058(.a(G245), .O(gate234inter7));
  inv1  gate1059(.a(G721), .O(gate234inter8));
  nand2 gate1060(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1061(.a(s_73), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1062(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1063(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1064(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1135(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1136(.a(gate236inter0), .b(s_84), .O(gate236inter1));
  and2  gate1137(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1138(.a(s_84), .O(gate236inter3));
  inv1  gate1139(.a(s_85), .O(gate236inter4));
  nand2 gate1140(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1141(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1142(.a(G251), .O(gate236inter7));
  inv1  gate1143(.a(G727), .O(gate236inter8));
  nand2 gate1144(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1145(.a(s_85), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1146(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1147(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1148(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1611(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1612(.a(gate238inter0), .b(s_152), .O(gate238inter1));
  and2  gate1613(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1614(.a(s_152), .O(gate238inter3));
  inv1  gate1615(.a(s_153), .O(gate238inter4));
  nand2 gate1616(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1617(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1618(.a(G257), .O(gate238inter7));
  inv1  gate1619(.a(G709), .O(gate238inter8));
  nand2 gate1620(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1621(.a(s_153), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1622(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1623(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1624(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate2171(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2172(.a(gate239inter0), .b(s_232), .O(gate239inter1));
  and2  gate2173(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2174(.a(s_232), .O(gate239inter3));
  inv1  gate2175(.a(s_233), .O(gate239inter4));
  nand2 gate2176(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2177(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2178(.a(G260), .O(gate239inter7));
  inv1  gate2179(.a(G712), .O(gate239inter8));
  nand2 gate2180(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2181(.a(s_233), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2182(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2183(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2184(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2885(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2886(.a(gate241inter0), .b(s_334), .O(gate241inter1));
  and2  gate2887(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2888(.a(s_334), .O(gate241inter3));
  inv1  gate2889(.a(s_335), .O(gate241inter4));
  nand2 gate2890(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2891(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2892(.a(G242), .O(gate241inter7));
  inv1  gate2893(.a(G730), .O(gate241inter8));
  nand2 gate2894(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2895(.a(s_335), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2896(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2897(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2898(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1765(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1766(.a(gate243inter0), .b(s_174), .O(gate243inter1));
  and2  gate1767(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1768(.a(s_174), .O(gate243inter3));
  inv1  gate1769(.a(s_175), .O(gate243inter4));
  nand2 gate1770(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1771(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1772(.a(G245), .O(gate243inter7));
  inv1  gate1773(.a(G733), .O(gate243inter8));
  nand2 gate1774(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1775(.a(s_175), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1776(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1777(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1778(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate3165(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate3166(.a(gate245inter0), .b(s_374), .O(gate245inter1));
  and2  gate3167(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate3168(.a(s_374), .O(gate245inter3));
  inv1  gate3169(.a(s_375), .O(gate245inter4));
  nand2 gate3170(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate3171(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate3172(.a(G248), .O(gate245inter7));
  inv1  gate3173(.a(G736), .O(gate245inter8));
  nand2 gate3174(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate3175(.a(s_375), .b(gate245inter3), .O(gate245inter10));
  nor2  gate3176(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate3177(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate3178(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2899(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2900(.a(gate247inter0), .b(s_336), .O(gate247inter1));
  and2  gate2901(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2902(.a(s_336), .O(gate247inter3));
  inv1  gate2903(.a(s_337), .O(gate247inter4));
  nand2 gate2904(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2905(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2906(.a(G251), .O(gate247inter7));
  inv1  gate2907(.a(G739), .O(gate247inter8));
  nand2 gate2908(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2909(.a(s_337), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2910(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2911(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2912(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1345(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1346(.a(gate251inter0), .b(s_114), .O(gate251inter1));
  and2  gate1347(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1348(.a(s_114), .O(gate251inter3));
  inv1  gate1349(.a(s_115), .O(gate251inter4));
  nand2 gate1350(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1351(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1352(.a(G257), .O(gate251inter7));
  inv1  gate1353(.a(G745), .O(gate251inter8));
  nand2 gate1354(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1355(.a(s_115), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1356(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1357(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1358(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1793(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1794(.a(gate252inter0), .b(s_178), .O(gate252inter1));
  and2  gate1795(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1796(.a(s_178), .O(gate252inter3));
  inv1  gate1797(.a(s_179), .O(gate252inter4));
  nand2 gate1798(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1799(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1800(.a(G709), .O(gate252inter7));
  inv1  gate1801(.a(G745), .O(gate252inter8));
  nand2 gate1802(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1803(.a(s_179), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1804(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1805(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1806(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2493(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2494(.a(gate254inter0), .b(s_278), .O(gate254inter1));
  and2  gate2495(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2496(.a(s_278), .O(gate254inter3));
  inv1  gate2497(.a(s_279), .O(gate254inter4));
  nand2 gate2498(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2499(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2500(.a(G712), .O(gate254inter7));
  inv1  gate2501(.a(G748), .O(gate254inter8));
  nand2 gate2502(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2503(.a(s_279), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2504(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2505(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2506(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate3095(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate3096(.a(gate258inter0), .b(s_364), .O(gate258inter1));
  and2  gate3097(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate3098(.a(s_364), .O(gate258inter3));
  inv1  gate3099(.a(s_365), .O(gate258inter4));
  nand2 gate3100(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate3101(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate3102(.a(G756), .O(gate258inter7));
  inv1  gate3103(.a(G757), .O(gate258inter8));
  nand2 gate3104(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate3105(.a(s_365), .b(gate258inter3), .O(gate258inter10));
  nor2  gate3106(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate3107(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate3108(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1555(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1556(.a(gate259inter0), .b(s_144), .O(gate259inter1));
  and2  gate1557(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1558(.a(s_144), .O(gate259inter3));
  inv1  gate1559(.a(s_145), .O(gate259inter4));
  nand2 gate1560(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1561(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1562(.a(G758), .O(gate259inter7));
  inv1  gate1563(.a(G759), .O(gate259inter8));
  nand2 gate1564(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1565(.a(s_145), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1566(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1567(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1568(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate2129(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2130(.a(gate260inter0), .b(s_226), .O(gate260inter1));
  and2  gate2131(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2132(.a(s_226), .O(gate260inter3));
  inv1  gate2133(.a(s_227), .O(gate260inter4));
  nand2 gate2134(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2135(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2136(.a(G760), .O(gate260inter7));
  inv1  gate2137(.a(G761), .O(gate260inter8));
  nand2 gate2138(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2139(.a(s_227), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2140(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2141(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2142(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1219(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1220(.a(gate262inter0), .b(s_96), .O(gate262inter1));
  and2  gate1221(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1222(.a(s_96), .O(gate262inter3));
  inv1  gate1223(.a(s_97), .O(gate262inter4));
  nand2 gate1224(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1225(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1226(.a(G764), .O(gate262inter7));
  inv1  gate1227(.a(G765), .O(gate262inter8));
  nand2 gate1228(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1229(.a(s_97), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1230(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1231(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1232(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1415(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1416(.a(gate263inter0), .b(s_124), .O(gate263inter1));
  and2  gate1417(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1418(.a(s_124), .O(gate263inter3));
  inv1  gate1419(.a(s_125), .O(gate263inter4));
  nand2 gate1420(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1421(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1422(.a(G766), .O(gate263inter7));
  inv1  gate1423(.a(G767), .O(gate263inter8));
  nand2 gate1424(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1425(.a(s_125), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1426(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1427(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1428(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1639(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1640(.a(gate264inter0), .b(s_156), .O(gate264inter1));
  and2  gate1641(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1642(.a(s_156), .O(gate264inter3));
  inv1  gate1643(.a(s_157), .O(gate264inter4));
  nand2 gate1644(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1645(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1646(.a(G768), .O(gate264inter7));
  inv1  gate1647(.a(G769), .O(gate264inter8));
  nand2 gate1648(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1649(.a(s_157), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1650(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1651(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1652(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate911(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate912(.a(gate269inter0), .b(s_52), .O(gate269inter1));
  and2  gate913(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate914(.a(s_52), .O(gate269inter3));
  inv1  gate915(.a(s_53), .O(gate269inter4));
  nand2 gate916(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate917(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate918(.a(G654), .O(gate269inter7));
  inv1  gate919(.a(G782), .O(gate269inter8));
  nand2 gate920(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate921(.a(s_53), .b(gate269inter3), .O(gate269inter10));
  nor2  gate922(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate923(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate924(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2339(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2340(.a(gate272inter0), .b(s_256), .O(gate272inter1));
  and2  gate2341(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2342(.a(s_256), .O(gate272inter3));
  inv1  gate2343(.a(s_257), .O(gate272inter4));
  nand2 gate2344(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2345(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2346(.a(G663), .O(gate272inter7));
  inv1  gate2347(.a(G791), .O(gate272inter8));
  nand2 gate2348(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2349(.a(s_257), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2350(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2351(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2352(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate3081(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate3082(.a(gate274inter0), .b(s_362), .O(gate274inter1));
  and2  gate3083(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate3084(.a(s_362), .O(gate274inter3));
  inv1  gate3085(.a(s_363), .O(gate274inter4));
  nand2 gate3086(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate3087(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate3088(.a(G770), .O(gate274inter7));
  inv1  gate3089(.a(G794), .O(gate274inter8));
  nand2 gate3090(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate3091(.a(s_363), .b(gate274inter3), .O(gate274inter10));
  nor2  gate3092(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate3093(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate3094(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1387(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1388(.a(gate275inter0), .b(s_120), .O(gate275inter1));
  and2  gate1389(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1390(.a(s_120), .O(gate275inter3));
  inv1  gate1391(.a(s_121), .O(gate275inter4));
  nand2 gate1392(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1393(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1394(.a(G645), .O(gate275inter7));
  inv1  gate1395(.a(G797), .O(gate275inter8));
  nand2 gate1396(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1397(.a(s_121), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1398(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1399(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1400(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1919(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1920(.a(gate282inter0), .b(s_196), .O(gate282inter1));
  and2  gate1921(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1922(.a(s_196), .O(gate282inter3));
  inv1  gate1923(.a(s_197), .O(gate282inter4));
  nand2 gate1924(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1925(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1926(.a(G782), .O(gate282inter7));
  inv1  gate1927(.a(G806), .O(gate282inter8));
  nand2 gate1928(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1929(.a(s_197), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1930(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1931(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1932(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2703(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2704(.a(gate285inter0), .b(s_308), .O(gate285inter1));
  and2  gate2705(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2706(.a(s_308), .O(gate285inter3));
  inv1  gate2707(.a(s_309), .O(gate285inter4));
  nand2 gate2708(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2709(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2710(.a(G660), .O(gate285inter7));
  inv1  gate2711(.a(G812), .O(gate285inter8));
  nand2 gate2712(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2713(.a(s_309), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2714(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2715(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2716(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1107(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1108(.a(gate286inter0), .b(s_80), .O(gate286inter1));
  and2  gate1109(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1110(.a(s_80), .O(gate286inter3));
  inv1  gate1111(.a(s_81), .O(gate286inter4));
  nand2 gate1112(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1113(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1114(.a(G788), .O(gate286inter7));
  inv1  gate1115(.a(G812), .O(gate286inter8));
  nand2 gate1116(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1117(.a(s_81), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1118(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1119(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1120(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate827(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate828(.a(gate287inter0), .b(s_40), .O(gate287inter1));
  and2  gate829(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate830(.a(s_40), .O(gate287inter3));
  inv1  gate831(.a(s_41), .O(gate287inter4));
  nand2 gate832(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate833(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate834(.a(G663), .O(gate287inter7));
  inv1  gate835(.a(G815), .O(gate287inter8));
  nand2 gate836(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate837(.a(s_41), .b(gate287inter3), .O(gate287inter10));
  nor2  gate838(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate839(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate840(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate925(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate926(.a(gate288inter0), .b(s_54), .O(gate288inter1));
  and2  gate927(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate928(.a(s_54), .O(gate288inter3));
  inv1  gate929(.a(s_55), .O(gate288inter4));
  nand2 gate930(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate931(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate932(.a(G791), .O(gate288inter7));
  inv1  gate933(.a(G815), .O(gate288inter8));
  nand2 gate934(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate935(.a(s_55), .b(gate288inter3), .O(gate288inter10));
  nor2  gate936(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate937(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate938(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate757(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate758(.a(gate289inter0), .b(s_30), .O(gate289inter1));
  and2  gate759(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate760(.a(s_30), .O(gate289inter3));
  inv1  gate761(.a(s_31), .O(gate289inter4));
  nand2 gate762(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate763(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate764(.a(G818), .O(gate289inter7));
  inv1  gate765(.a(G819), .O(gate289inter8));
  nand2 gate766(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate767(.a(s_31), .b(gate289inter3), .O(gate289inter10));
  nor2  gate768(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate769(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate770(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1191(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1192(.a(gate291inter0), .b(s_92), .O(gate291inter1));
  and2  gate1193(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1194(.a(s_92), .O(gate291inter3));
  inv1  gate1195(.a(s_93), .O(gate291inter4));
  nand2 gate1196(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1197(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1198(.a(G822), .O(gate291inter7));
  inv1  gate1199(.a(G823), .O(gate291inter8));
  nand2 gate1200(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1201(.a(s_93), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1202(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1203(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1204(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate2241(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2242(.a(gate292inter0), .b(s_242), .O(gate292inter1));
  and2  gate2243(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2244(.a(s_242), .O(gate292inter3));
  inv1  gate2245(.a(s_243), .O(gate292inter4));
  nand2 gate2246(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2247(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2248(.a(G824), .O(gate292inter7));
  inv1  gate2249(.a(G825), .O(gate292inter8));
  nand2 gate2250(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2251(.a(s_243), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2252(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2253(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2254(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2997(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2998(.a(gate295inter0), .b(s_350), .O(gate295inter1));
  and2  gate2999(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate3000(.a(s_350), .O(gate295inter3));
  inv1  gate3001(.a(s_351), .O(gate295inter4));
  nand2 gate3002(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate3003(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate3004(.a(G830), .O(gate295inter7));
  inv1  gate3005(.a(G831), .O(gate295inter8));
  nand2 gate3006(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate3007(.a(s_351), .b(gate295inter3), .O(gate295inter10));
  nor2  gate3008(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate3009(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate3010(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1905(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1906(.a(gate296inter0), .b(s_194), .O(gate296inter1));
  and2  gate1907(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1908(.a(s_194), .O(gate296inter3));
  inv1  gate1909(.a(s_195), .O(gate296inter4));
  nand2 gate1910(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1911(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1912(.a(G826), .O(gate296inter7));
  inv1  gate1913(.a(G827), .O(gate296inter8));
  nand2 gate1914(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1915(.a(s_195), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1916(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1917(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1918(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2661(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2662(.a(gate387inter0), .b(s_302), .O(gate387inter1));
  and2  gate2663(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2664(.a(s_302), .O(gate387inter3));
  inv1  gate2665(.a(s_303), .O(gate387inter4));
  nand2 gate2666(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2667(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2668(.a(G1), .O(gate387inter7));
  inv1  gate2669(.a(G1036), .O(gate387inter8));
  nand2 gate2670(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2671(.a(s_303), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2672(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2673(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2674(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1513(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1514(.a(gate389inter0), .b(s_138), .O(gate389inter1));
  and2  gate1515(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1516(.a(s_138), .O(gate389inter3));
  inv1  gate1517(.a(s_139), .O(gate389inter4));
  nand2 gate1518(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1519(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1520(.a(G3), .O(gate389inter7));
  inv1  gate1521(.a(G1042), .O(gate389inter8));
  nand2 gate1522(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1523(.a(s_139), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1524(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1525(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1526(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate2003(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2004(.a(gate390inter0), .b(s_208), .O(gate390inter1));
  and2  gate2005(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2006(.a(s_208), .O(gate390inter3));
  inv1  gate2007(.a(s_209), .O(gate390inter4));
  nand2 gate2008(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2009(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2010(.a(G4), .O(gate390inter7));
  inv1  gate2011(.a(G1045), .O(gate390inter8));
  nand2 gate2012(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2013(.a(s_209), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2014(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2015(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2016(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2325(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2326(.a(gate392inter0), .b(s_254), .O(gate392inter1));
  and2  gate2327(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2328(.a(s_254), .O(gate392inter3));
  inv1  gate2329(.a(s_255), .O(gate392inter4));
  nand2 gate2330(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2331(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2332(.a(G6), .O(gate392inter7));
  inv1  gate2333(.a(G1051), .O(gate392inter8));
  nand2 gate2334(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2335(.a(s_255), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2336(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2337(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2338(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2101(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2102(.a(gate394inter0), .b(s_222), .O(gate394inter1));
  and2  gate2103(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2104(.a(s_222), .O(gate394inter3));
  inv1  gate2105(.a(s_223), .O(gate394inter4));
  nand2 gate2106(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2107(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2108(.a(G8), .O(gate394inter7));
  inv1  gate2109(.a(G1057), .O(gate394inter8));
  nand2 gate2110(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2111(.a(s_223), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2112(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2113(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2114(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate967(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate968(.a(gate395inter0), .b(s_60), .O(gate395inter1));
  and2  gate969(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate970(.a(s_60), .O(gate395inter3));
  inv1  gate971(.a(s_61), .O(gate395inter4));
  nand2 gate972(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate973(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate974(.a(G9), .O(gate395inter7));
  inv1  gate975(.a(G1060), .O(gate395inter8));
  nand2 gate976(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate977(.a(s_61), .b(gate395inter3), .O(gate395inter10));
  nor2  gate978(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate979(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate980(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1989(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1990(.a(gate396inter0), .b(s_206), .O(gate396inter1));
  and2  gate1991(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1992(.a(s_206), .O(gate396inter3));
  inv1  gate1993(.a(s_207), .O(gate396inter4));
  nand2 gate1994(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1995(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1996(.a(G10), .O(gate396inter7));
  inv1  gate1997(.a(G1063), .O(gate396inter8));
  nand2 gate1998(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1999(.a(s_207), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2000(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2001(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2002(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate659(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate660(.a(gate397inter0), .b(s_16), .O(gate397inter1));
  and2  gate661(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate662(.a(s_16), .O(gate397inter3));
  inv1  gate663(.a(s_17), .O(gate397inter4));
  nand2 gate664(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate665(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate666(.a(G11), .O(gate397inter7));
  inv1  gate667(.a(G1066), .O(gate397inter8));
  nand2 gate668(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate669(.a(s_17), .b(gate397inter3), .O(gate397inter10));
  nor2  gate670(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate671(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate672(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1233(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1234(.a(gate399inter0), .b(s_98), .O(gate399inter1));
  and2  gate1235(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1236(.a(s_98), .O(gate399inter3));
  inv1  gate1237(.a(s_99), .O(gate399inter4));
  nand2 gate1238(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1239(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1240(.a(G13), .O(gate399inter7));
  inv1  gate1241(.a(G1072), .O(gate399inter8));
  nand2 gate1242(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1243(.a(s_99), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1244(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1245(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1246(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1947(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1948(.a(gate401inter0), .b(s_200), .O(gate401inter1));
  and2  gate1949(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1950(.a(s_200), .O(gate401inter3));
  inv1  gate1951(.a(s_201), .O(gate401inter4));
  nand2 gate1952(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1953(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1954(.a(G15), .O(gate401inter7));
  inv1  gate1955(.a(G1078), .O(gate401inter8));
  nand2 gate1956(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1957(.a(s_201), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1958(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1959(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1960(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate3193(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate3194(.a(gate408inter0), .b(s_378), .O(gate408inter1));
  and2  gate3195(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate3196(.a(s_378), .O(gate408inter3));
  inv1  gate3197(.a(s_379), .O(gate408inter4));
  nand2 gate3198(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate3199(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate3200(.a(G22), .O(gate408inter7));
  inv1  gate3201(.a(G1099), .O(gate408inter8));
  nand2 gate3202(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate3203(.a(s_379), .b(gate408inter3), .O(gate408inter10));
  nor2  gate3204(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate3205(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate3206(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2185(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2186(.a(gate410inter0), .b(s_234), .O(gate410inter1));
  and2  gate2187(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2188(.a(s_234), .O(gate410inter3));
  inv1  gate2189(.a(s_235), .O(gate410inter4));
  nand2 gate2190(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2191(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2192(.a(G24), .O(gate410inter7));
  inv1  gate2193(.a(G1105), .O(gate410inter8));
  nand2 gate2194(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2195(.a(s_235), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2196(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2197(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2198(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1849(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1850(.a(gate413inter0), .b(s_186), .O(gate413inter1));
  and2  gate1851(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1852(.a(s_186), .O(gate413inter3));
  inv1  gate1853(.a(s_187), .O(gate413inter4));
  nand2 gate1854(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1855(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1856(.a(G27), .O(gate413inter7));
  inv1  gate1857(.a(G1114), .O(gate413inter8));
  nand2 gate1858(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1859(.a(s_187), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1860(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1861(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1862(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2073(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2074(.a(gate414inter0), .b(s_218), .O(gate414inter1));
  and2  gate2075(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2076(.a(s_218), .O(gate414inter3));
  inv1  gate2077(.a(s_219), .O(gate414inter4));
  nand2 gate2078(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2079(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2080(.a(G28), .O(gate414inter7));
  inv1  gate2081(.a(G1117), .O(gate414inter8));
  nand2 gate2082(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2083(.a(s_219), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2084(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2085(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2086(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2451(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2452(.a(gate416inter0), .b(s_272), .O(gate416inter1));
  and2  gate2453(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2454(.a(s_272), .O(gate416inter3));
  inv1  gate2455(.a(s_273), .O(gate416inter4));
  nand2 gate2456(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2457(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2458(.a(G30), .O(gate416inter7));
  inv1  gate2459(.a(G1123), .O(gate416inter8));
  nand2 gate2460(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2461(.a(s_273), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2462(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2463(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2464(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2381(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2382(.a(gate419inter0), .b(s_262), .O(gate419inter1));
  and2  gate2383(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2384(.a(s_262), .O(gate419inter3));
  inv1  gate2385(.a(s_263), .O(gate419inter4));
  nand2 gate2386(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2387(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2388(.a(G1), .O(gate419inter7));
  inv1  gate2389(.a(G1132), .O(gate419inter8));
  nand2 gate2390(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2391(.a(s_263), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2392(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2393(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2394(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2871(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2872(.a(gate420inter0), .b(s_332), .O(gate420inter1));
  and2  gate2873(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2874(.a(s_332), .O(gate420inter3));
  inv1  gate2875(.a(s_333), .O(gate420inter4));
  nand2 gate2876(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2877(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2878(.a(G1036), .O(gate420inter7));
  inv1  gate2879(.a(G1132), .O(gate420inter8));
  nand2 gate2880(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2881(.a(s_333), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2882(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2883(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2884(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2647(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2648(.a(gate421inter0), .b(s_300), .O(gate421inter1));
  and2  gate2649(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2650(.a(s_300), .O(gate421inter3));
  inv1  gate2651(.a(s_301), .O(gate421inter4));
  nand2 gate2652(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2653(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2654(.a(G2), .O(gate421inter7));
  inv1  gate2655(.a(G1135), .O(gate421inter8));
  nand2 gate2656(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2657(.a(s_301), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2658(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2659(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2660(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2773(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2774(.a(gate422inter0), .b(s_318), .O(gate422inter1));
  and2  gate2775(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2776(.a(s_318), .O(gate422inter3));
  inv1  gate2777(.a(s_319), .O(gate422inter4));
  nand2 gate2778(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2779(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2780(.a(G1039), .O(gate422inter7));
  inv1  gate2781(.a(G1135), .O(gate422inter8));
  nand2 gate2782(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2783(.a(s_319), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2784(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2785(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2786(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate981(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate982(.a(gate424inter0), .b(s_62), .O(gate424inter1));
  and2  gate983(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate984(.a(s_62), .O(gate424inter3));
  inv1  gate985(.a(s_63), .O(gate424inter4));
  nand2 gate986(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate987(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate988(.a(G1042), .O(gate424inter7));
  inv1  gate989(.a(G1138), .O(gate424inter8));
  nand2 gate990(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate991(.a(s_63), .b(gate424inter3), .O(gate424inter10));
  nor2  gate992(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate993(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate994(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1401(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1402(.a(gate428inter0), .b(s_122), .O(gate428inter1));
  and2  gate1403(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1404(.a(s_122), .O(gate428inter3));
  inv1  gate1405(.a(s_123), .O(gate428inter4));
  nand2 gate1406(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1407(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1408(.a(G1048), .O(gate428inter7));
  inv1  gate1409(.a(G1144), .O(gate428inter8));
  nand2 gate1410(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1411(.a(s_123), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1412(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1413(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1414(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1709(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1710(.a(gate429inter0), .b(s_166), .O(gate429inter1));
  and2  gate1711(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1712(.a(s_166), .O(gate429inter3));
  inv1  gate1713(.a(s_167), .O(gate429inter4));
  nand2 gate1714(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1715(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1716(.a(G6), .O(gate429inter7));
  inv1  gate1717(.a(G1147), .O(gate429inter8));
  nand2 gate1718(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1719(.a(s_167), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1720(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1721(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1722(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate687(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate688(.a(gate431inter0), .b(s_20), .O(gate431inter1));
  and2  gate689(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate690(.a(s_20), .O(gate431inter3));
  inv1  gate691(.a(s_21), .O(gate431inter4));
  nand2 gate692(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate693(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate694(.a(G7), .O(gate431inter7));
  inv1  gate695(.a(G1150), .O(gate431inter8));
  nand2 gate696(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate697(.a(s_21), .b(gate431inter3), .O(gate431inter10));
  nor2  gate698(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate699(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate700(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1149(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1150(.a(gate432inter0), .b(s_86), .O(gate432inter1));
  and2  gate1151(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1152(.a(s_86), .O(gate432inter3));
  inv1  gate1153(.a(s_87), .O(gate432inter4));
  nand2 gate1154(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1155(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1156(.a(G1054), .O(gate432inter7));
  inv1  gate1157(.a(G1150), .O(gate432inter8));
  nand2 gate1158(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1159(.a(s_87), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1160(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1161(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1162(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2717(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2718(.a(gate434inter0), .b(s_310), .O(gate434inter1));
  and2  gate2719(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2720(.a(s_310), .O(gate434inter3));
  inv1  gate2721(.a(s_311), .O(gate434inter4));
  nand2 gate2722(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2723(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2724(.a(G1057), .O(gate434inter7));
  inv1  gate2725(.a(G1153), .O(gate434inter8));
  nand2 gate2726(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2727(.a(s_311), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2728(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2729(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2730(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1065(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1066(.a(gate440inter0), .b(s_74), .O(gate440inter1));
  and2  gate1067(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1068(.a(s_74), .O(gate440inter3));
  inv1  gate1069(.a(s_75), .O(gate440inter4));
  nand2 gate1070(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1071(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1072(.a(G1066), .O(gate440inter7));
  inv1  gate1073(.a(G1162), .O(gate440inter8));
  nand2 gate1074(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1075(.a(s_75), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1076(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1077(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1078(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate3109(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate3110(.a(gate441inter0), .b(s_366), .O(gate441inter1));
  and2  gate3111(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate3112(.a(s_366), .O(gate441inter3));
  inv1  gate3113(.a(s_367), .O(gate441inter4));
  nand2 gate3114(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate3115(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate3116(.a(G12), .O(gate441inter7));
  inv1  gate3117(.a(G1165), .O(gate441inter8));
  nand2 gate3118(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate3119(.a(s_367), .b(gate441inter3), .O(gate441inter10));
  nor2  gate3120(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate3121(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate3122(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate701(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate702(.a(gate442inter0), .b(s_22), .O(gate442inter1));
  and2  gate703(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate704(.a(s_22), .O(gate442inter3));
  inv1  gate705(.a(s_23), .O(gate442inter4));
  nand2 gate706(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate707(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate708(.a(G1069), .O(gate442inter7));
  inv1  gate709(.a(G1165), .O(gate442inter8));
  nand2 gate710(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate711(.a(s_23), .b(gate442inter3), .O(gate442inter10));
  nor2  gate712(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate713(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate714(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate2045(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2046(.a(gate443inter0), .b(s_214), .O(gate443inter1));
  and2  gate2047(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2048(.a(s_214), .O(gate443inter3));
  inv1  gate2049(.a(s_215), .O(gate443inter4));
  nand2 gate2050(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2051(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2052(.a(G13), .O(gate443inter7));
  inv1  gate2053(.a(G1168), .O(gate443inter8));
  nand2 gate2054(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2055(.a(s_215), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2056(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2057(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2058(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2829(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2830(.a(gate446inter0), .b(s_326), .O(gate446inter1));
  and2  gate2831(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2832(.a(s_326), .O(gate446inter3));
  inv1  gate2833(.a(s_327), .O(gate446inter4));
  nand2 gate2834(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2835(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2836(.a(G1075), .O(gate446inter7));
  inv1  gate2837(.a(G1171), .O(gate446inter8));
  nand2 gate2838(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2839(.a(s_327), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2840(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2841(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2842(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate3025(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate3026(.a(gate447inter0), .b(s_354), .O(gate447inter1));
  and2  gate3027(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate3028(.a(s_354), .O(gate447inter3));
  inv1  gate3029(.a(s_355), .O(gate447inter4));
  nand2 gate3030(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate3031(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate3032(.a(G15), .O(gate447inter7));
  inv1  gate3033(.a(G1174), .O(gate447inter8));
  nand2 gate3034(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate3035(.a(s_355), .b(gate447inter3), .O(gate447inter10));
  nor2  gate3036(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate3037(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate3038(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1961(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1962(.a(gate452inter0), .b(s_202), .O(gate452inter1));
  and2  gate1963(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1964(.a(s_202), .O(gate452inter3));
  inv1  gate1965(.a(s_203), .O(gate452inter4));
  nand2 gate1966(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1967(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1968(.a(G1084), .O(gate452inter7));
  inv1  gate1969(.a(G1180), .O(gate452inter8));
  nand2 gate1970(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1971(.a(s_203), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1972(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1973(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1974(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2955(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2956(.a(gate455inter0), .b(s_344), .O(gate455inter1));
  and2  gate2957(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2958(.a(s_344), .O(gate455inter3));
  inv1  gate2959(.a(s_345), .O(gate455inter4));
  nand2 gate2960(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2961(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2962(.a(G19), .O(gate455inter7));
  inv1  gate2963(.a(G1186), .O(gate455inter8));
  nand2 gate2964(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2965(.a(s_345), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2966(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2967(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2968(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate771(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate772(.a(gate457inter0), .b(s_32), .O(gate457inter1));
  and2  gate773(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate774(.a(s_32), .O(gate457inter3));
  inv1  gate775(.a(s_33), .O(gate457inter4));
  nand2 gate776(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate777(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate778(.a(G20), .O(gate457inter7));
  inv1  gate779(.a(G1189), .O(gate457inter8));
  nand2 gate780(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate781(.a(s_33), .b(gate457inter3), .O(gate457inter10));
  nor2  gate782(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate783(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate784(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate883(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate884(.a(gate459inter0), .b(s_48), .O(gate459inter1));
  and2  gate885(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate886(.a(s_48), .O(gate459inter3));
  inv1  gate887(.a(s_49), .O(gate459inter4));
  nand2 gate888(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate889(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate890(.a(G21), .O(gate459inter7));
  inv1  gate891(.a(G1192), .O(gate459inter8));
  nand2 gate892(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate893(.a(s_49), .b(gate459inter3), .O(gate459inter10));
  nor2  gate894(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate895(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate896(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate855(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate856(.a(gate460inter0), .b(s_44), .O(gate460inter1));
  and2  gate857(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate858(.a(s_44), .O(gate460inter3));
  inv1  gate859(.a(s_45), .O(gate460inter4));
  nand2 gate860(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate861(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate862(.a(G1096), .O(gate460inter7));
  inv1  gate863(.a(G1192), .O(gate460inter8));
  nand2 gate864(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate865(.a(s_45), .b(gate460inter3), .O(gate460inter10));
  nor2  gate866(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate867(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate868(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2857(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2858(.a(gate461inter0), .b(s_330), .O(gate461inter1));
  and2  gate2859(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2860(.a(s_330), .O(gate461inter3));
  inv1  gate2861(.a(s_331), .O(gate461inter4));
  nand2 gate2862(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2863(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2864(.a(G22), .O(gate461inter7));
  inv1  gate2865(.a(G1195), .O(gate461inter8));
  nand2 gate2866(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2867(.a(s_331), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2868(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2869(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2870(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate673(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate674(.a(gate463inter0), .b(s_18), .O(gate463inter1));
  and2  gate675(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate676(.a(s_18), .O(gate463inter3));
  inv1  gate677(.a(s_19), .O(gate463inter4));
  nand2 gate678(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate679(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate680(.a(G23), .O(gate463inter7));
  inv1  gate681(.a(G1198), .O(gate463inter8));
  nand2 gate682(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate683(.a(s_19), .b(gate463inter3), .O(gate463inter10));
  nor2  gate684(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate685(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate686(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2605(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2606(.a(gate465inter0), .b(s_294), .O(gate465inter1));
  and2  gate2607(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2608(.a(s_294), .O(gate465inter3));
  inv1  gate2609(.a(s_295), .O(gate465inter4));
  nand2 gate2610(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2611(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2612(.a(G24), .O(gate465inter7));
  inv1  gate2613(.a(G1201), .O(gate465inter8));
  nand2 gate2614(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2615(.a(s_295), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2616(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2617(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2618(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2549(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2550(.a(gate466inter0), .b(s_286), .O(gate466inter1));
  and2  gate2551(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2552(.a(s_286), .O(gate466inter3));
  inv1  gate2553(.a(s_287), .O(gate466inter4));
  nand2 gate2554(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2555(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2556(.a(G1105), .O(gate466inter7));
  inv1  gate2557(.a(G1201), .O(gate466inter8));
  nand2 gate2558(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2559(.a(s_287), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2560(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2561(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2562(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1373(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1374(.a(gate467inter0), .b(s_118), .O(gate467inter1));
  and2  gate1375(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1376(.a(s_118), .O(gate467inter3));
  inv1  gate1377(.a(s_119), .O(gate467inter4));
  nand2 gate1378(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1379(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1380(.a(G25), .O(gate467inter7));
  inv1  gate1381(.a(G1204), .O(gate467inter8));
  nand2 gate1382(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1383(.a(s_119), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1384(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1385(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1386(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate2115(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2116(.a(gate468inter0), .b(s_224), .O(gate468inter1));
  and2  gate2117(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2118(.a(s_224), .O(gate468inter3));
  inv1  gate2119(.a(s_225), .O(gate468inter4));
  nand2 gate2120(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2121(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2122(.a(G1108), .O(gate468inter7));
  inv1  gate2123(.a(G1204), .O(gate468inter8));
  nand2 gate2124(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2125(.a(s_225), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2126(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2127(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2128(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1485(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1486(.a(gate470inter0), .b(s_134), .O(gate470inter1));
  and2  gate1487(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1488(.a(s_134), .O(gate470inter3));
  inv1  gate1489(.a(s_135), .O(gate470inter4));
  nand2 gate1490(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1491(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1492(.a(G1111), .O(gate470inter7));
  inv1  gate1493(.a(G1207), .O(gate470inter8));
  nand2 gate1494(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1495(.a(s_135), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1496(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1497(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1498(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2577(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2578(.a(gate471inter0), .b(s_290), .O(gate471inter1));
  and2  gate2579(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2580(.a(s_290), .O(gate471inter3));
  inv1  gate2581(.a(s_291), .O(gate471inter4));
  nand2 gate2582(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2583(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2584(.a(G27), .O(gate471inter7));
  inv1  gate2585(.a(G1210), .O(gate471inter8));
  nand2 gate2586(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2587(.a(s_291), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2588(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2589(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2590(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate3137(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate3138(.a(gate477inter0), .b(s_370), .O(gate477inter1));
  and2  gate3139(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate3140(.a(s_370), .O(gate477inter3));
  inv1  gate3141(.a(s_371), .O(gate477inter4));
  nand2 gate3142(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate3143(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate3144(.a(G30), .O(gate477inter7));
  inv1  gate3145(.a(G1219), .O(gate477inter8));
  nand2 gate3146(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate3147(.a(s_371), .b(gate477inter3), .O(gate477inter10));
  nor2  gate3148(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate3149(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate3150(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate813(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate814(.a(gate478inter0), .b(s_38), .O(gate478inter1));
  and2  gate815(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate816(.a(s_38), .O(gate478inter3));
  inv1  gate817(.a(s_39), .O(gate478inter4));
  nand2 gate818(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate819(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate820(.a(G1123), .O(gate478inter7));
  inv1  gate821(.a(G1219), .O(gate478inter8));
  nand2 gate822(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate823(.a(s_39), .b(gate478inter3), .O(gate478inter10));
  nor2  gate824(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate825(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate826(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2465(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2466(.a(gate480inter0), .b(s_274), .O(gate480inter1));
  and2  gate2467(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2468(.a(s_274), .O(gate480inter3));
  inv1  gate2469(.a(s_275), .O(gate480inter4));
  nand2 gate2470(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2471(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2472(.a(G1126), .O(gate480inter7));
  inv1  gate2473(.a(G1222), .O(gate480inter8));
  nand2 gate2474(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2475(.a(s_275), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2476(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2477(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2478(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1163(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1164(.a(gate482inter0), .b(s_88), .O(gate482inter1));
  and2  gate1165(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1166(.a(s_88), .O(gate482inter3));
  inv1  gate1167(.a(s_89), .O(gate482inter4));
  nand2 gate1168(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1169(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1170(.a(G1129), .O(gate482inter7));
  inv1  gate1171(.a(G1225), .O(gate482inter8));
  nand2 gate1172(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1173(.a(s_89), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1174(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1175(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1176(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2983(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2984(.a(gate486inter0), .b(s_348), .O(gate486inter1));
  and2  gate2985(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2986(.a(s_348), .O(gate486inter3));
  inv1  gate2987(.a(s_349), .O(gate486inter4));
  nand2 gate2988(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2989(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2990(.a(G1234), .O(gate486inter7));
  inv1  gate2991(.a(G1235), .O(gate486inter8));
  nand2 gate2992(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2993(.a(s_349), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2994(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2995(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2996(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2535(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2536(.a(gate487inter0), .b(s_284), .O(gate487inter1));
  and2  gate2537(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2538(.a(s_284), .O(gate487inter3));
  inv1  gate2539(.a(s_285), .O(gate487inter4));
  nand2 gate2540(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2541(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2542(.a(G1236), .O(gate487inter7));
  inv1  gate2543(.a(G1237), .O(gate487inter8));
  nand2 gate2544(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2545(.a(s_285), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2546(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2547(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2548(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2031(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2032(.a(gate490inter0), .b(s_212), .O(gate490inter1));
  and2  gate2033(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2034(.a(s_212), .O(gate490inter3));
  inv1  gate2035(.a(s_213), .O(gate490inter4));
  nand2 gate2036(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2037(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2038(.a(G1242), .O(gate490inter7));
  inv1  gate2039(.a(G1243), .O(gate490inter8));
  nand2 gate2040(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2041(.a(s_213), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2042(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2043(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2044(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1681(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1682(.a(gate492inter0), .b(s_162), .O(gate492inter1));
  and2  gate1683(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1684(.a(s_162), .O(gate492inter3));
  inv1  gate1685(.a(s_163), .O(gate492inter4));
  nand2 gate1686(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1687(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1688(.a(G1246), .O(gate492inter7));
  inv1  gate1689(.a(G1247), .O(gate492inter8));
  nand2 gate1690(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1691(.a(s_163), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1692(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1693(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1694(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1093(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1094(.a(gate493inter0), .b(s_78), .O(gate493inter1));
  and2  gate1095(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1096(.a(s_78), .O(gate493inter3));
  inv1  gate1097(.a(s_79), .O(gate493inter4));
  nand2 gate1098(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1099(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1100(.a(G1248), .O(gate493inter7));
  inv1  gate1101(.a(G1249), .O(gate493inter8));
  nand2 gate1102(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1103(.a(s_79), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1104(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1105(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1106(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1891(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1892(.a(gate494inter0), .b(s_192), .O(gate494inter1));
  and2  gate1893(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1894(.a(s_192), .O(gate494inter3));
  inv1  gate1895(.a(s_193), .O(gate494inter4));
  nand2 gate1896(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1897(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1898(.a(G1250), .O(gate494inter7));
  inv1  gate1899(.a(G1251), .O(gate494inter8));
  nand2 gate1900(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1901(.a(s_193), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1902(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1903(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1904(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2297(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2298(.a(gate495inter0), .b(s_250), .O(gate495inter1));
  and2  gate2299(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2300(.a(s_250), .O(gate495inter3));
  inv1  gate2301(.a(s_251), .O(gate495inter4));
  nand2 gate2302(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2303(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2304(.a(G1252), .O(gate495inter7));
  inv1  gate2305(.a(G1253), .O(gate495inter8));
  nand2 gate2306(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2307(.a(s_251), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2308(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2309(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2310(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate869(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate870(.a(gate500inter0), .b(s_46), .O(gate500inter1));
  and2  gate871(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate872(.a(s_46), .O(gate500inter3));
  inv1  gate873(.a(s_47), .O(gate500inter4));
  nand2 gate874(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate875(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate876(.a(G1262), .O(gate500inter7));
  inv1  gate877(.a(G1263), .O(gate500inter8));
  nand2 gate878(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate879(.a(s_47), .b(gate500inter3), .O(gate500inter10));
  nor2  gate880(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate881(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate882(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1863(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1864(.a(gate501inter0), .b(s_188), .O(gate501inter1));
  and2  gate1865(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1866(.a(s_188), .O(gate501inter3));
  inv1  gate1867(.a(s_189), .O(gate501inter4));
  nand2 gate1868(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1869(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1870(.a(G1264), .O(gate501inter7));
  inv1  gate1871(.a(G1265), .O(gate501inter8));
  nand2 gate1872(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1873(.a(s_189), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1874(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1875(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1876(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2479(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2480(.a(gate502inter0), .b(s_276), .O(gate502inter1));
  and2  gate2481(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2482(.a(s_276), .O(gate502inter3));
  inv1  gate2483(.a(s_277), .O(gate502inter4));
  nand2 gate2484(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2485(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2486(.a(G1266), .O(gate502inter7));
  inv1  gate2487(.a(G1267), .O(gate502inter8));
  nand2 gate2488(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2489(.a(s_277), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2490(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2491(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2492(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1653(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1654(.a(gate503inter0), .b(s_158), .O(gate503inter1));
  and2  gate1655(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1656(.a(s_158), .O(gate503inter3));
  inv1  gate1657(.a(s_159), .O(gate503inter4));
  nand2 gate1658(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1659(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1660(.a(G1268), .O(gate503inter7));
  inv1  gate1661(.a(G1269), .O(gate503inter8));
  nand2 gate1662(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1663(.a(s_159), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1664(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1665(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1666(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate617(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate618(.a(gate504inter0), .b(s_10), .O(gate504inter1));
  and2  gate619(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate620(.a(s_10), .O(gate504inter3));
  inv1  gate621(.a(s_11), .O(gate504inter4));
  nand2 gate622(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate623(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate624(.a(G1270), .O(gate504inter7));
  inv1  gate625(.a(G1271), .O(gate504inter8));
  nand2 gate626(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate627(.a(s_11), .b(gate504inter3), .O(gate504inter10));
  nor2  gate628(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate629(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate630(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1037(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1038(.a(gate505inter0), .b(s_70), .O(gate505inter1));
  and2  gate1039(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1040(.a(s_70), .O(gate505inter3));
  inv1  gate1041(.a(s_71), .O(gate505inter4));
  nand2 gate1042(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1043(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1044(.a(G1272), .O(gate505inter7));
  inv1  gate1045(.a(G1273), .O(gate505inter8));
  nand2 gate1046(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1047(.a(s_71), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1048(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1049(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1050(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate547(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate548(.a(gate506inter0), .b(s_0), .O(gate506inter1));
  and2  gate549(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate550(.a(s_0), .O(gate506inter3));
  inv1  gate551(.a(s_1), .O(gate506inter4));
  nand2 gate552(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate553(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate554(.a(G1274), .O(gate506inter7));
  inv1  gate555(.a(G1275), .O(gate506inter8));
  nand2 gate556(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate557(.a(s_1), .b(gate506inter3), .O(gate506inter10));
  nor2  gate558(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate559(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate560(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2633(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2634(.a(gate510inter0), .b(s_298), .O(gate510inter1));
  and2  gate2635(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2636(.a(s_298), .O(gate510inter3));
  inv1  gate2637(.a(s_299), .O(gate510inter4));
  nand2 gate2638(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2639(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2640(.a(G1282), .O(gate510inter7));
  inv1  gate2641(.a(G1283), .O(gate510inter8));
  nand2 gate2642(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2643(.a(s_299), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2644(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2645(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2646(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate3263(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate3264(.a(gate511inter0), .b(s_388), .O(gate511inter1));
  and2  gate3265(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate3266(.a(s_388), .O(gate511inter3));
  inv1  gate3267(.a(s_389), .O(gate511inter4));
  nand2 gate3268(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate3269(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate3270(.a(G1284), .O(gate511inter7));
  inv1  gate3271(.a(G1285), .O(gate511inter8));
  nand2 gate3272(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate3273(.a(s_389), .b(gate511inter3), .O(gate511inter10));
  nor2  gate3274(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate3275(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate3276(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1569(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1570(.a(gate513inter0), .b(s_146), .O(gate513inter1));
  and2  gate1571(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1572(.a(s_146), .O(gate513inter3));
  inv1  gate1573(.a(s_147), .O(gate513inter4));
  nand2 gate1574(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1575(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1576(.a(G1288), .O(gate513inter7));
  inv1  gate1577(.a(G1289), .O(gate513inter8));
  nand2 gate1578(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1579(.a(s_147), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1580(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1581(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1582(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule