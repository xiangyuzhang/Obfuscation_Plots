module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1289(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1290(.a(gate10inter0), .b(s_106), .O(gate10inter1));
  and2  gate1291(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1292(.a(s_106), .O(gate10inter3));
  inv1  gate1293(.a(s_107), .O(gate10inter4));
  nand2 gate1294(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1295(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1296(.a(G3), .O(gate10inter7));
  inv1  gate1297(.a(G4), .O(gate10inter8));
  nand2 gate1298(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1299(.a(s_107), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1300(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1301(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1302(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2395(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2396(.a(gate12inter0), .b(s_264), .O(gate12inter1));
  and2  gate2397(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2398(.a(s_264), .O(gate12inter3));
  inv1  gate2399(.a(s_265), .O(gate12inter4));
  nand2 gate2400(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2401(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2402(.a(G7), .O(gate12inter7));
  inv1  gate2403(.a(G8), .O(gate12inter8));
  nand2 gate2404(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2405(.a(s_265), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2406(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2407(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2408(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1135(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1136(.a(gate15inter0), .b(s_84), .O(gate15inter1));
  and2  gate1137(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1138(.a(s_84), .O(gate15inter3));
  inv1  gate1139(.a(s_85), .O(gate15inter4));
  nand2 gate1140(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1141(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1142(.a(G13), .O(gate15inter7));
  inv1  gate1143(.a(G14), .O(gate15inter8));
  nand2 gate1144(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1145(.a(s_85), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1146(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1147(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1148(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate631(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate632(.a(gate19inter0), .b(s_12), .O(gate19inter1));
  and2  gate633(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate634(.a(s_12), .O(gate19inter3));
  inv1  gate635(.a(s_13), .O(gate19inter4));
  nand2 gate636(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate637(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate638(.a(G21), .O(gate19inter7));
  inv1  gate639(.a(G22), .O(gate19inter8));
  nand2 gate640(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate641(.a(s_13), .b(gate19inter3), .O(gate19inter10));
  nor2  gate642(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate643(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate644(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate547(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate548(.a(gate21inter0), .b(s_0), .O(gate21inter1));
  and2  gate549(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate550(.a(s_0), .O(gate21inter3));
  inv1  gate551(.a(s_1), .O(gate21inter4));
  nand2 gate552(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate553(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate554(.a(G25), .O(gate21inter7));
  inv1  gate555(.a(G26), .O(gate21inter8));
  nand2 gate556(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate557(.a(s_1), .b(gate21inter3), .O(gate21inter10));
  nor2  gate558(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate559(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate560(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate757(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate758(.a(gate24inter0), .b(s_30), .O(gate24inter1));
  and2  gate759(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate760(.a(s_30), .O(gate24inter3));
  inv1  gate761(.a(s_31), .O(gate24inter4));
  nand2 gate762(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate763(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate764(.a(G31), .O(gate24inter7));
  inv1  gate765(.a(G32), .O(gate24inter8));
  nand2 gate766(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate767(.a(s_31), .b(gate24inter3), .O(gate24inter10));
  nor2  gate768(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate769(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate770(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate2773(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2774(.a(gate25inter0), .b(s_318), .O(gate25inter1));
  and2  gate2775(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2776(.a(s_318), .O(gate25inter3));
  inv1  gate2777(.a(s_319), .O(gate25inter4));
  nand2 gate2778(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2779(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2780(.a(G1), .O(gate25inter7));
  inv1  gate2781(.a(G5), .O(gate25inter8));
  nand2 gate2782(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2783(.a(s_319), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2784(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2785(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2786(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate561(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate562(.a(gate26inter0), .b(s_2), .O(gate26inter1));
  and2  gate563(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate564(.a(s_2), .O(gate26inter3));
  inv1  gate565(.a(s_3), .O(gate26inter4));
  nand2 gate566(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate567(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate568(.a(G9), .O(gate26inter7));
  inv1  gate569(.a(G13), .O(gate26inter8));
  nand2 gate570(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate571(.a(s_3), .b(gate26inter3), .O(gate26inter10));
  nor2  gate572(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate573(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate574(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate2759(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2760(.a(gate27inter0), .b(s_316), .O(gate27inter1));
  and2  gate2761(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2762(.a(s_316), .O(gate27inter3));
  inv1  gate2763(.a(s_317), .O(gate27inter4));
  nand2 gate2764(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2765(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2766(.a(G2), .O(gate27inter7));
  inv1  gate2767(.a(G6), .O(gate27inter8));
  nand2 gate2768(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2769(.a(s_317), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2770(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2771(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2772(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2605(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2606(.a(gate31inter0), .b(s_294), .O(gate31inter1));
  and2  gate2607(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2608(.a(s_294), .O(gate31inter3));
  inv1  gate2609(.a(s_295), .O(gate31inter4));
  nand2 gate2610(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2611(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2612(.a(G4), .O(gate31inter7));
  inv1  gate2613(.a(G8), .O(gate31inter8));
  nand2 gate2614(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2615(.a(s_295), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2616(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2617(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2618(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate855(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate856(.a(gate32inter0), .b(s_44), .O(gate32inter1));
  and2  gate857(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate858(.a(s_44), .O(gate32inter3));
  inv1  gate859(.a(s_45), .O(gate32inter4));
  nand2 gate860(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate861(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate862(.a(G12), .O(gate32inter7));
  inv1  gate863(.a(G16), .O(gate32inter8));
  nand2 gate864(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate865(.a(s_45), .b(gate32inter3), .O(gate32inter10));
  nor2  gate866(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate867(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate868(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1793(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1794(.a(gate34inter0), .b(s_178), .O(gate34inter1));
  and2  gate1795(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1796(.a(s_178), .O(gate34inter3));
  inv1  gate1797(.a(s_179), .O(gate34inter4));
  nand2 gate1798(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1799(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1800(.a(G25), .O(gate34inter7));
  inv1  gate1801(.a(G29), .O(gate34inter8));
  nand2 gate1802(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1803(.a(s_179), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1804(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1805(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1806(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1317(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1318(.a(gate37inter0), .b(s_110), .O(gate37inter1));
  and2  gate1319(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1320(.a(s_110), .O(gate37inter3));
  inv1  gate1321(.a(s_111), .O(gate37inter4));
  nand2 gate1322(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1323(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1324(.a(G19), .O(gate37inter7));
  inv1  gate1325(.a(G23), .O(gate37inter8));
  nand2 gate1326(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1327(.a(s_111), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1328(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1329(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1330(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate925(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate926(.a(gate42inter0), .b(s_54), .O(gate42inter1));
  and2  gate927(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate928(.a(s_54), .O(gate42inter3));
  inv1  gate929(.a(s_55), .O(gate42inter4));
  nand2 gate930(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate931(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate932(.a(G2), .O(gate42inter7));
  inv1  gate933(.a(G266), .O(gate42inter8));
  nand2 gate934(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate935(.a(s_55), .b(gate42inter3), .O(gate42inter10));
  nor2  gate936(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate937(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate938(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1163(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1164(.a(gate44inter0), .b(s_88), .O(gate44inter1));
  and2  gate1165(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1166(.a(s_88), .O(gate44inter3));
  inv1  gate1167(.a(s_89), .O(gate44inter4));
  nand2 gate1168(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1169(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1170(.a(G4), .O(gate44inter7));
  inv1  gate1171(.a(G269), .O(gate44inter8));
  nand2 gate1172(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1173(.a(s_89), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1174(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1175(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1176(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2703(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2704(.a(gate50inter0), .b(s_308), .O(gate50inter1));
  and2  gate2705(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2706(.a(s_308), .O(gate50inter3));
  inv1  gate2707(.a(s_309), .O(gate50inter4));
  nand2 gate2708(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2709(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2710(.a(G10), .O(gate50inter7));
  inv1  gate2711(.a(G278), .O(gate50inter8));
  nand2 gate2712(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2713(.a(s_309), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2714(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2715(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2716(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1121(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1122(.a(gate55inter0), .b(s_82), .O(gate55inter1));
  and2  gate1123(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1124(.a(s_82), .O(gate55inter3));
  inv1  gate1125(.a(s_83), .O(gate55inter4));
  nand2 gate1126(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1127(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1128(.a(G15), .O(gate55inter7));
  inv1  gate1129(.a(G287), .O(gate55inter8));
  nand2 gate1130(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1131(.a(s_83), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1132(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1133(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1134(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1247(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1248(.a(gate57inter0), .b(s_100), .O(gate57inter1));
  and2  gate1249(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1250(.a(s_100), .O(gate57inter3));
  inv1  gate1251(.a(s_101), .O(gate57inter4));
  nand2 gate1252(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1253(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1254(.a(G17), .O(gate57inter7));
  inv1  gate1255(.a(G290), .O(gate57inter8));
  nand2 gate1256(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1257(.a(s_101), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1258(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1259(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1260(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1947(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1948(.a(gate61inter0), .b(s_200), .O(gate61inter1));
  and2  gate1949(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1950(.a(s_200), .O(gate61inter3));
  inv1  gate1951(.a(s_201), .O(gate61inter4));
  nand2 gate1952(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1953(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1954(.a(G21), .O(gate61inter7));
  inv1  gate1955(.a(G296), .O(gate61inter8));
  nand2 gate1956(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1957(.a(s_201), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1958(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1959(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1960(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1457(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1458(.a(gate62inter0), .b(s_130), .O(gate62inter1));
  and2  gate1459(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1460(.a(s_130), .O(gate62inter3));
  inv1  gate1461(.a(s_131), .O(gate62inter4));
  nand2 gate1462(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1463(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1464(.a(G22), .O(gate62inter7));
  inv1  gate1465(.a(G296), .O(gate62inter8));
  nand2 gate1466(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1467(.a(s_131), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1468(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1469(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1470(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1639(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1640(.a(gate63inter0), .b(s_156), .O(gate63inter1));
  and2  gate1641(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1642(.a(s_156), .O(gate63inter3));
  inv1  gate1643(.a(s_157), .O(gate63inter4));
  nand2 gate1644(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1645(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1646(.a(G23), .O(gate63inter7));
  inv1  gate1647(.a(G299), .O(gate63inter8));
  nand2 gate1648(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1649(.a(s_157), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1650(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1651(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1652(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2549(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2550(.a(gate64inter0), .b(s_286), .O(gate64inter1));
  and2  gate2551(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2552(.a(s_286), .O(gate64inter3));
  inv1  gate2553(.a(s_287), .O(gate64inter4));
  nand2 gate2554(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2555(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2556(.a(G24), .O(gate64inter7));
  inv1  gate2557(.a(G299), .O(gate64inter8));
  nand2 gate2558(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2559(.a(s_287), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2560(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2561(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2562(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate2437(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2438(.a(gate65inter0), .b(s_270), .O(gate65inter1));
  and2  gate2439(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2440(.a(s_270), .O(gate65inter3));
  inv1  gate2441(.a(s_271), .O(gate65inter4));
  nand2 gate2442(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2443(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2444(.a(G25), .O(gate65inter7));
  inv1  gate2445(.a(G302), .O(gate65inter8));
  nand2 gate2446(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2447(.a(s_271), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2448(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2449(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2450(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1387(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1388(.a(gate75inter0), .b(s_120), .O(gate75inter1));
  and2  gate1389(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1390(.a(s_120), .O(gate75inter3));
  inv1  gate1391(.a(s_121), .O(gate75inter4));
  nand2 gate1392(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1393(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1394(.a(G9), .O(gate75inter7));
  inv1  gate1395(.a(G317), .O(gate75inter8));
  nand2 gate1396(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1397(.a(s_121), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1398(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1399(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1400(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1877(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1878(.a(gate79inter0), .b(s_190), .O(gate79inter1));
  and2  gate1879(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1880(.a(s_190), .O(gate79inter3));
  inv1  gate1881(.a(s_191), .O(gate79inter4));
  nand2 gate1882(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1883(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1884(.a(G10), .O(gate79inter7));
  inv1  gate1885(.a(G323), .O(gate79inter8));
  nand2 gate1886(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1887(.a(s_191), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1888(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1889(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1890(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1513(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1514(.a(gate83inter0), .b(s_138), .O(gate83inter1));
  and2  gate1515(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1516(.a(s_138), .O(gate83inter3));
  inv1  gate1517(.a(s_139), .O(gate83inter4));
  nand2 gate1518(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1519(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1520(.a(G11), .O(gate83inter7));
  inv1  gate1521(.a(G329), .O(gate83inter8));
  nand2 gate1522(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1523(.a(s_139), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1524(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1525(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1526(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate2563(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2564(.a(gate84inter0), .b(s_288), .O(gate84inter1));
  and2  gate2565(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2566(.a(s_288), .O(gate84inter3));
  inv1  gate2567(.a(s_289), .O(gate84inter4));
  nand2 gate2568(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2569(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2570(.a(G15), .O(gate84inter7));
  inv1  gate2571(.a(G329), .O(gate84inter8));
  nand2 gate2572(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2573(.a(s_289), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2574(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2575(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2576(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2213(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2214(.a(gate92inter0), .b(s_238), .O(gate92inter1));
  and2  gate2215(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2216(.a(s_238), .O(gate92inter3));
  inv1  gate2217(.a(s_239), .O(gate92inter4));
  nand2 gate2218(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2219(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2220(.a(G29), .O(gate92inter7));
  inv1  gate2221(.a(G341), .O(gate92inter8));
  nand2 gate2222(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2223(.a(s_239), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2224(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2225(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2226(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate575(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate576(.a(gate97inter0), .b(s_4), .O(gate97inter1));
  and2  gate577(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate578(.a(s_4), .O(gate97inter3));
  inv1  gate579(.a(s_5), .O(gate97inter4));
  nand2 gate580(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate581(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate582(.a(G19), .O(gate97inter7));
  inv1  gate583(.a(G350), .O(gate97inter8));
  nand2 gate584(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate585(.a(s_5), .b(gate97inter3), .O(gate97inter10));
  nor2  gate586(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate587(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate588(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1737(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1738(.a(gate98inter0), .b(s_170), .O(gate98inter1));
  and2  gate1739(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1740(.a(s_170), .O(gate98inter3));
  inv1  gate1741(.a(s_171), .O(gate98inter4));
  nand2 gate1742(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1743(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1744(.a(G23), .O(gate98inter7));
  inv1  gate1745(.a(G350), .O(gate98inter8));
  nand2 gate1746(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1747(.a(s_171), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1748(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1749(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1750(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate967(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate968(.a(gate99inter0), .b(s_60), .O(gate99inter1));
  and2  gate969(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate970(.a(s_60), .O(gate99inter3));
  inv1  gate971(.a(s_61), .O(gate99inter4));
  nand2 gate972(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate973(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate974(.a(G27), .O(gate99inter7));
  inv1  gate975(.a(G353), .O(gate99inter8));
  nand2 gate976(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate977(.a(s_61), .b(gate99inter3), .O(gate99inter10));
  nor2  gate978(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate979(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate980(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate2325(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2326(.a(gate100inter0), .b(s_254), .O(gate100inter1));
  and2  gate2327(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2328(.a(s_254), .O(gate100inter3));
  inv1  gate2329(.a(s_255), .O(gate100inter4));
  nand2 gate2330(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2331(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2332(.a(G31), .O(gate100inter7));
  inv1  gate2333(.a(G353), .O(gate100inter8));
  nand2 gate2334(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2335(.a(s_255), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2336(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2337(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2338(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1023(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1024(.a(gate102inter0), .b(s_68), .O(gate102inter1));
  and2  gate1025(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1026(.a(s_68), .O(gate102inter3));
  inv1  gate1027(.a(s_69), .O(gate102inter4));
  nand2 gate1028(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1029(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1030(.a(G24), .O(gate102inter7));
  inv1  gate1031(.a(G356), .O(gate102inter8));
  nand2 gate1032(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1033(.a(s_69), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1034(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1035(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1036(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2227(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2228(.a(gate106inter0), .b(s_240), .O(gate106inter1));
  and2  gate2229(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2230(.a(s_240), .O(gate106inter3));
  inv1  gate2231(.a(s_241), .O(gate106inter4));
  nand2 gate2232(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2233(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2234(.a(G364), .O(gate106inter7));
  inv1  gate2235(.a(G365), .O(gate106inter8));
  nand2 gate2236(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2237(.a(s_241), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2238(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2239(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2240(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1961(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1962(.a(gate111inter0), .b(s_202), .O(gate111inter1));
  and2  gate1963(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1964(.a(s_202), .O(gate111inter3));
  inv1  gate1965(.a(s_203), .O(gate111inter4));
  nand2 gate1966(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1967(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1968(.a(G374), .O(gate111inter7));
  inv1  gate1969(.a(G375), .O(gate111inter8));
  nand2 gate1970(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1971(.a(s_203), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1972(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1973(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1974(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1471(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1472(.a(gate112inter0), .b(s_132), .O(gate112inter1));
  and2  gate1473(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1474(.a(s_132), .O(gate112inter3));
  inv1  gate1475(.a(s_133), .O(gate112inter4));
  nand2 gate1476(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1477(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1478(.a(G376), .O(gate112inter7));
  inv1  gate1479(.a(G377), .O(gate112inter8));
  nand2 gate1480(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1481(.a(s_133), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1482(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1483(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1484(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2619(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2620(.a(gate118inter0), .b(s_296), .O(gate118inter1));
  and2  gate2621(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2622(.a(s_296), .O(gate118inter3));
  inv1  gate2623(.a(s_297), .O(gate118inter4));
  nand2 gate2624(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2625(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2626(.a(G388), .O(gate118inter7));
  inv1  gate2627(.a(G389), .O(gate118inter8));
  nand2 gate2628(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2629(.a(s_297), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2630(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2631(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2632(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate2157(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2158(.a(gate119inter0), .b(s_230), .O(gate119inter1));
  and2  gate2159(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2160(.a(s_230), .O(gate119inter3));
  inv1  gate2161(.a(s_231), .O(gate119inter4));
  nand2 gate2162(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2163(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2164(.a(G390), .O(gate119inter7));
  inv1  gate2165(.a(G391), .O(gate119inter8));
  nand2 gate2166(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2167(.a(s_231), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2168(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2169(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2170(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1849(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1850(.a(gate123inter0), .b(s_186), .O(gate123inter1));
  and2  gate1851(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1852(.a(s_186), .O(gate123inter3));
  inv1  gate1853(.a(s_187), .O(gate123inter4));
  nand2 gate1854(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1855(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1856(.a(G398), .O(gate123inter7));
  inv1  gate1857(.a(G399), .O(gate123inter8));
  nand2 gate1858(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1859(.a(s_187), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1860(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1861(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1862(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1975(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1976(.a(gate124inter0), .b(s_204), .O(gate124inter1));
  and2  gate1977(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1978(.a(s_204), .O(gate124inter3));
  inv1  gate1979(.a(s_205), .O(gate124inter4));
  nand2 gate1980(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1981(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1982(.a(G400), .O(gate124inter7));
  inv1  gate1983(.a(G401), .O(gate124inter8));
  nand2 gate1984(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1985(.a(s_205), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1986(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1987(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1988(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate869(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate870(.a(gate131inter0), .b(s_46), .O(gate131inter1));
  and2  gate871(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate872(.a(s_46), .O(gate131inter3));
  inv1  gate873(.a(s_47), .O(gate131inter4));
  nand2 gate874(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate875(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate876(.a(G414), .O(gate131inter7));
  inv1  gate877(.a(G415), .O(gate131inter8));
  nand2 gate878(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate879(.a(s_47), .b(gate131inter3), .O(gate131inter10));
  nor2  gate880(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate881(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate882(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1765(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1766(.a(gate132inter0), .b(s_174), .O(gate132inter1));
  and2  gate1767(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1768(.a(s_174), .O(gate132inter3));
  inv1  gate1769(.a(s_175), .O(gate132inter4));
  nand2 gate1770(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1771(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1772(.a(G416), .O(gate132inter7));
  inv1  gate1773(.a(G417), .O(gate132inter8));
  nand2 gate1774(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1775(.a(s_175), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1776(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1777(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1778(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate659(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate660(.a(gate133inter0), .b(s_16), .O(gate133inter1));
  and2  gate661(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate662(.a(s_16), .O(gate133inter3));
  inv1  gate663(.a(s_17), .O(gate133inter4));
  nand2 gate664(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate665(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate666(.a(G418), .O(gate133inter7));
  inv1  gate667(.a(G419), .O(gate133inter8));
  nand2 gate668(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate669(.a(s_17), .b(gate133inter3), .O(gate133inter10));
  nor2  gate670(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate671(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate672(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2731(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2732(.a(gate138inter0), .b(s_312), .O(gate138inter1));
  and2  gate2733(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2734(.a(s_312), .O(gate138inter3));
  inv1  gate2735(.a(s_313), .O(gate138inter4));
  nand2 gate2736(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2737(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2738(.a(G432), .O(gate138inter7));
  inv1  gate2739(.a(G435), .O(gate138inter8));
  nand2 gate2740(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2741(.a(s_313), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2742(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2743(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2744(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate939(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate940(.a(gate147inter0), .b(s_56), .O(gate147inter1));
  and2  gate941(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate942(.a(s_56), .O(gate147inter3));
  inv1  gate943(.a(s_57), .O(gate147inter4));
  nand2 gate944(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate945(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate946(.a(G486), .O(gate147inter7));
  inv1  gate947(.a(G489), .O(gate147inter8));
  nand2 gate948(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate949(.a(s_57), .b(gate147inter3), .O(gate147inter10));
  nor2  gate950(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate951(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate952(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1807(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1808(.a(gate150inter0), .b(s_180), .O(gate150inter1));
  and2  gate1809(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1810(.a(s_180), .O(gate150inter3));
  inv1  gate1811(.a(s_181), .O(gate150inter4));
  nand2 gate1812(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1813(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1814(.a(G504), .O(gate150inter7));
  inv1  gate1815(.a(G507), .O(gate150inter8));
  nand2 gate1816(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1817(.a(s_181), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1818(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1819(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1820(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1401(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1402(.a(gate151inter0), .b(s_122), .O(gate151inter1));
  and2  gate1403(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1404(.a(s_122), .O(gate151inter3));
  inv1  gate1405(.a(s_123), .O(gate151inter4));
  nand2 gate1406(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1407(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1408(.a(G510), .O(gate151inter7));
  inv1  gate1409(.a(G513), .O(gate151inter8));
  nand2 gate1410(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1411(.a(s_123), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1412(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1413(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1414(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1373(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1374(.a(gate152inter0), .b(s_118), .O(gate152inter1));
  and2  gate1375(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1376(.a(s_118), .O(gate152inter3));
  inv1  gate1377(.a(s_119), .O(gate152inter4));
  nand2 gate1378(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1379(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1380(.a(G516), .O(gate152inter7));
  inv1  gate1381(.a(G519), .O(gate152inter8));
  nand2 gate1382(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1383(.a(s_119), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1384(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1385(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1386(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate603(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate604(.a(gate154inter0), .b(s_8), .O(gate154inter1));
  and2  gate605(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate606(.a(s_8), .O(gate154inter3));
  inv1  gate607(.a(s_9), .O(gate154inter4));
  nand2 gate608(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate609(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate610(.a(G429), .O(gate154inter7));
  inv1  gate611(.a(G522), .O(gate154inter8));
  nand2 gate612(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate613(.a(s_9), .b(gate154inter3), .O(gate154inter10));
  nor2  gate614(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate615(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate616(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate673(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate674(.a(gate155inter0), .b(s_18), .O(gate155inter1));
  and2  gate675(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate676(.a(s_18), .O(gate155inter3));
  inv1  gate677(.a(s_19), .O(gate155inter4));
  nand2 gate678(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate679(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate680(.a(G432), .O(gate155inter7));
  inv1  gate681(.a(G525), .O(gate155inter8));
  nand2 gate682(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate683(.a(s_19), .b(gate155inter3), .O(gate155inter10));
  nor2  gate684(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate685(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate686(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2129(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2130(.a(gate157inter0), .b(s_226), .O(gate157inter1));
  and2  gate2131(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2132(.a(s_226), .O(gate157inter3));
  inv1  gate2133(.a(s_227), .O(gate157inter4));
  nand2 gate2134(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2135(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2136(.a(G438), .O(gate157inter7));
  inv1  gate2137(.a(G528), .O(gate157inter8));
  nand2 gate2138(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2139(.a(s_227), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2140(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2141(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2142(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate2073(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2074(.a(gate168inter0), .b(s_218), .O(gate168inter1));
  and2  gate2075(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2076(.a(s_218), .O(gate168inter3));
  inv1  gate2077(.a(s_219), .O(gate168inter4));
  nand2 gate2078(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2079(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2080(.a(G471), .O(gate168inter7));
  inv1  gate2081(.a(G543), .O(gate168inter8));
  nand2 gate2082(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2083(.a(s_219), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2084(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2085(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2086(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate995(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate996(.a(gate170inter0), .b(s_64), .O(gate170inter1));
  and2  gate997(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate998(.a(s_64), .O(gate170inter3));
  inv1  gate999(.a(s_65), .O(gate170inter4));
  nand2 gate1000(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1001(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1002(.a(G477), .O(gate170inter7));
  inv1  gate1003(.a(G546), .O(gate170inter8));
  nand2 gate1004(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1005(.a(s_65), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1006(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1007(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1008(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1527(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1528(.a(gate174inter0), .b(s_140), .O(gate174inter1));
  and2  gate1529(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1530(.a(s_140), .O(gate174inter3));
  inv1  gate1531(.a(s_141), .O(gate174inter4));
  nand2 gate1532(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1533(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1534(.a(G489), .O(gate174inter7));
  inv1  gate1535(.a(G552), .O(gate174inter8));
  nand2 gate1536(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1537(.a(s_141), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1538(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1539(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1540(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate715(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate716(.a(gate178inter0), .b(s_24), .O(gate178inter1));
  and2  gate717(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate718(.a(s_24), .O(gate178inter3));
  inv1  gate719(.a(s_25), .O(gate178inter4));
  nand2 gate720(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate721(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate722(.a(G501), .O(gate178inter7));
  inv1  gate723(.a(G558), .O(gate178inter8));
  nand2 gate724(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate725(.a(s_25), .b(gate178inter3), .O(gate178inter10));
  nor2  gate726(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate727(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate728(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate645(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate646(.a(gate179inter0), .b(s_14), .O(gate179inter1));
  and2  gate647(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate648(.a(s_14), .O(gate179inter3));
  inv1  gate649(.a(s_15), .O(gate179inter4));
  nand2 gate650(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate651(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate652(.a(G504), .O(gate179inter7));
  inv1  gate653(.a(G561), .O(gate179inter8));
  nand2 gate654(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate655(.a(s_15), .b(gate179inter3), .O(gate179inter10));
  nor2  gate656(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate657(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate658(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2297(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2298(.a(gate183inter0), .b(s_250), .O(gate183inter1));
  and2  gate2299(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2300(.a(s_250), .O(gate183inter3));
  inv1  gate2301(.a(s_251), .O(gate183inter4));
  nand2 gate2302(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2303(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2304(.a(G516), .O(gate183inter7));
  inv1  gate2305(.a(G567), .O(gate183inter8));
  nand2 gate2306(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2307(.a(s_251), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2308(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2309(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2310(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2465(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2466(.a(gate191inter0), .b(s_274), .O(gate191inter1));
  and2  gate2467(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2468(.a(s_274), .O(gate191inter3));
  inv1  gate2469(.a(s_275), .O(gate191inter4));
  nand2 gate2470(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2471(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2472(.a(G582), .O(gate191inter7));
  inv1  gate2473(.a(G583), .O(gate191inter8));
  nand2 gate2474(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2475(.a(s_275), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2476(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2477(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2478(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2311(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2312(.a(gate192inter0), .b(s_252), .O(gate192inter1));
  and2  gate2313(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2314(.a(s_252), .O(gate192inter3));
  inv1  gate2315(.a(s_253), .O(gate192inter4));
  nand2 gate2316(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2317(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2318(.a(G584), .O(gate192inter7));
  inv1  gate2319(.a(G585), .O(gate192inter8));
  nand2 gate2320(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2321(.a(s_253), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2322(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2323(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2324(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2087(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2088(.a(gate195inter0), .b(s_220), .O(gate195inter1));
  and2  gate2089(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2090(.a(s_220), .O(gate195inter3));
  inv1  gate2091(.a(s_221), .O(gate195inter4));
  nand2 gate2092(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2093(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2094(.a(G590), .O(gate195inter7));
  inv1  gate2095(.a(G591), .O(gate195inter8));
  nand2 gate2096(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2097(.a(s_221), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2098(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2099(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2100(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2059(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2060(.a(gate198inter0), .b(s_216), .O(gate198inter1));
  and2  gate2061(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2062(.a(s_216), .O(gate198inter3));
  inv1  gate2063(.a(s_217), .O(gate198inter4));
  nand2 gate2064(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2065(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2066(.a(G596), .O(gate198inter7));
  inv1  gate2067(.a(G597), .O(gate198inter8));
  nand2 gate2068(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2069(.a(s_217), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2070(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2071(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2072(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1429(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1430(.a(gate200inter0), .b(s_126), .O(gate200inter1));
  and2  gate1431(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1432(.a(s_126), .O(gate200inter3));
  inv1  gate1433(.a(s_127), .O(gate200inter4));
  nand2 gate1434(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1435(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1436(.a(G600), .O(gate200inter7));
  inv1  gate1437(.a(G601), .O(gate200inter8));
  nand2 gate1438(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1439(.a(s_127), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1440(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1441(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1442(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1695(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1696(.a(gate201inter0), .b(s_164), .O(gate201inter1));
  and2  gate1697(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1698(.a(s_164), .O(gate201inter3));
  inv1  gate1699(.a(s_165), .O(gate201inter4));
  nand2 gate1700(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1701(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1702(.a(G602), .O(gate201inter7));
  inv1  gate1703(.a(G607), .O(gate201inter8));
  nand2 gate1704(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1705(.a(s_165), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1706(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1707(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1708(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1667(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1668(.a(gate204inter0), .b(s_160), .O(gate204inter1));
  and2  gate1669(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1670(.a(s_160), .O(gate204inter3));
  inv1  gate1671(.a(s_161), .O(gate204inter4));
  nand2 gate1672(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1673(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1674(.a(G607), .O(gate204inter7));
  inv1  gate1675(.a(G617), .O(gate204inter8));
  nand2 gate1676(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1677(.a(s_161), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1678(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1679(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1680(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1079(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1080(.a(gate205inter0), .b(s_76), .O(gate205inter1));
  and2  gate1081(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1082(.a(s_76), .O(gate205inter3));
  inv1  gate1083(.a(s_77), .O(gate205inter4));
  nand2 gate1084(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1085(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1086(.a(G622), .O(gate205inter7));
  inv1  gate1087(.a(G627), .O(gate205inter8));
  nand2 gate1088(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1089(.a(s_77), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1090(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1091(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1092(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2507(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2508(.a(gate206inter0), .b(s_280), .O(gate206inter1));
  and2  gate2509(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2510(.a(s_280), .O(gate206inter3));
  inv1  gate2511(.a(s_281), .O(gate206inter4));
  nand2 gate2512(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2513(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2514(.a(G632), .O(gate206inter7));
  inv1  gate2515(.a(G637), .O(gate206inter8));
  nand2 gate2516(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2517(.a(s_281), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2518(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2519(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2520(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1919(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1920(.a(gate207inter0), .b(s_196), .O(gate207inter1));
  and2  gate1921(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1922(.a(s_196), .O(gate207inter3));
  inv1  gate1923(.a(s_197), .O(gate207inter4));
  nand2 gate1924(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1925(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1926(.a(G622), .O(gate207inter7));
  inv1  gate1927(.a(G632), .O(gate207inter8));
  nand2 gate1928(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1929(.a(s_197), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1930(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1931(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1932(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1345(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1346(.a(gate208inter0), .b(s_114), .O(gate208inter1));
  and2  gate1347(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1348(.a(s_114), .O(gate208inter3));
  inv1  gate1349(.a(s_115), .O(gate208inter4));
  nand2 gate1350(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1351(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1352(.a(G627), .O(gate208inter7));
  inv1  gate1353(.a(G637), .O(gate208inter8));
  nand2 gate1354(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1355(.a(s_115), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1356(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1357(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1358(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2283(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2284(.a(gate211inter0), .b(s_248), .O(gate211inter1));
  and2  gate2285(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2286(.a(s_248), .O(gate211inter3));
  inv1  gate2287(.a(s_249), .O(gate211inter4));
  nand2 gate2288(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2289(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2290(.a(G612), .O(gate211inter7));
  inv1  gate2291(.a(G669), .O(gate211inter8));
  nand2 gate2292(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2293(.a(s_249), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2294(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2295(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2296(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate2675(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2676(.a(gate212inter0), .b(s_304), .O(gate212inter1));
  and2  gate2677(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2678(.a(s_304), .O(gate212inter3));
  inv1  gate2679(.a(s_305), .O(gate212inter4));
  nand2 gate2680(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2681(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2682(.a(G617), .O(gate212inter7));
  inv1  gate2683(.a(G669), .O(gate212inter8));
  nand2 gate2684(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2685(.a(s_305), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2686(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2687(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2688(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1751(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1752(.a(gate214inter0), .b(s_172), .O(gate214inter1));
  and2  gate1753(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1754(.a(s_172), .O(gate214inter3));
  inv1  gate1755(.a(s_173), .O(gate214inter4));
  nand2 gate1756(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1757(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1758(.a(G612), .O(gate214inter7));
  inv1  gate1759(.a(G672), .O(gate214inter8));
  nand2 gate1760(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1761(.a(s_173), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1762(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1763(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1764(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1779(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1780(.a(gate215inter0), .b(s_176), .O(gate215inter1));
  and2  gate1781(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1782(.a(s_176), .O(gate215inter3));
  inv1  gate1783(.a(s_177), .O(gate215inter4));
  nand2 gate1784(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1785(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1786(.a(G607), .O(gate215inter7));
  inv1  gate1787(.a(G675), .O(gate215inter8));
  nand2 gate1788(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1789(.a(s_177), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1790(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1791(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1792(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1233(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1234(.a(gate216inter0), .b(s_98), .O(gate216inter1));
  and2  gate1235(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1236(.a(s_98), .O(gate216inter3));
  inv1  gate1237(.a(s_99), .O(gate216inter4));
  nand2 gate1238(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1239(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1240(.a(G617), .O(gate216inter7));
  inv1  gate1241(.a(G675), .O(gate216inter8));
  nand2 gate1242(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1243(.a(s_99), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1244(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1245(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1246(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1933(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1934(.a(gate221inter0), .b(s_198), .O(gate221inter1));
  and2  gate1935(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1936(.a(s_198), .O(gate221inter3));
  inv1  gate1937(.a(s_199), .O(gate221inter4));
  nand2 gate1938(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1939(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1940(.a(G622), .O(gate221inter7));
  inv1  gate1941(.a(G684), .O(gate221inter8));
  nand2 gate1942(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1943(.a(s_199), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1944(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1945(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1946(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate771(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate772(.a(gate223inter0), .b(s_32), .O(gate223inter1));
  and2  gate773(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate774(.a(s_32), .O(gate223inter3));
  inv1  gate775(.a(s_33), .O(gate223inter4));
  nand2 gate776(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate777(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate778(.a(G627), .O(gate223inter7));
  inv1  gate779(.a(G687), .O(gate223inter8));
  nand2 gate780(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate781(.a(s_33), .b(gate223inter3), .O(gate223inter10));
  nor2  gate782(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate783(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate784(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate2031(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2032(.a(gate224inter0), .b(s_212), .O(gate224inter1));
  and2  gate2033(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2034(.a(s_212), .O(gate224inter3));
  inv1  gate2035(.a(s_213), .O(gate224inter4));
  nand2 gate2036(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2037(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2038(.a(G637), .O(gate224inter7));
  inv1  gate2039(.a(G687), .O(gate224inter8));
  nand2 gate2040(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2041(.a(s_213), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2042(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2043(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2044(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1569(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1570(.a(gate225inter0), .b(s_146), .O(gate225inter1));
  and2  gate1571(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1572(.a(s_146), .O(gate225inter3));
  inv1  gate1573(.a(s_147), .O(gate225inter4));
  nand2 gate1574(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1575(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1576(.a(G690), .O(gate225inter7));
  inv1  gate1577(.a(G691), .O(gate225inter8));
  nand2 gate1578(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1579(.a(s_147), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1580(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1581(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1582(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1653(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1654(.a(gate230inter0), .b(s_158), .O(gate230inter1));
  and2  gate1655(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1656(.a(s_158), .O(gate230inter3));
  inv1  gate1657(.a(s_159), .O(gate230inter4));
  nand2 gate1658(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1659(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1660(.a(G700), .O(gate230inter7));
  inv1  gate1661(.a(G701), .O(gate230inter8));
  nand2 gate1662(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1663(.a(s_159), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1664(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1665(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1666(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1863(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1864(.a(gate231inter0), .b(s_188), .O(gate231inter1));
  and2  gate1865(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1866(.a(s_188), .O(gate231inter3));
  inv1  gate1867(.a(s_189), .O(gate231inter4));
  nand2 gate1868(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1869(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1870(.a(G702), .O(gate231inter7));
  inv1  gate1871(.a(G703), .O(gate231inter8));
  nand2 gate1872(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1873(.a(s_189), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1874(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1875(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1876(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2535(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2536(.a(gate232inter0), .b(s_284), .O(gate232inter1));
  and2  gate2537(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2538(.a(s_284), .O(gate232inter3));
  inv1  gate2539(.a(s_285), .O(gate232inter4));
  nand2 gate2540(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2541(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2542(.a(G704), .O(gate232inter7));
  inv1  gate2543(.a(G705), .O(gate232inter8));
  nand2 gate2544(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2545(.a(s_285), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2546(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2547(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2548(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1597(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1598(.a(gate234inter0), .b(s_150), .O(gate234inter1));
  and2  gate1599(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1600(.a(s_150), .O(gate234inter3));
  inv1  gate1601(.a(s_151), .O(gate234inter4));
  nand2 gate1602(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1603(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1604(.a(G245), .O(gate234inter7));
  inv1  gate1605(.a(G721), .O(gate234inter8));
  nand2 gate1606(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1607(.a(s_151), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1608(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1609(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1610(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1149(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1150(.a(gate236inter0), .b(s_86), .O(gate236inter1));
  and2  gate1151(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1152(.a(s_86), .O(gate236inter3));
  inv1  gate1153(.a(s_87), .O(gate236inter4));
  nand2 gate1154(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1155(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1156(.a(G251), .O(gate236inter7));
  inv1  gate1157(.a(G727), .O(gate236inter8));
  nand2 gate1158(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1159(.a(s_87), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1160(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1161(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1162(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate2255(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2256(.a(gate237inter0), .b(s_244), .O(gate237inter1));
  and2  gate2257(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2258(.a(s_244), .O(gate237inter3));
  inv1  gate2259(.a(s_245), .O(gate237inter4));
  nand2 gate2260(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2261(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2262(.a(G254), .O(gate237inter7));
  inv1  gate2263(.a(G706), .O(gate237inter8));
  nand2 gate2264(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2265(.a(s_245), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2266(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2267(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2268(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate785(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate786(.a(gate239inter0), .b(s_34), .O(gate239inter1));
  and2  gate787(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate788(.a(s_34), .O(gate239inter3));
  inv1  gate789(.a(s_35), .O(gate239inter4));
  nand2 gate790(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate791(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate792(.a(G260), .O(gate239inter7));
  inv1  gate793(.a(G712), .O(gate239inter8));
  nand2 gate794(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate795(.a(s_35), .b(gate239inter3), .O(gate239inter10));
  nor2  gate796(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate797(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate798(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate2339(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2340(.a(gate240inter0), .b(s_256), .O(gate240inter1));
  and2  gate2341(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2342(.a(s_256), .O(gate240inter3));
  inv1  gate2343(.a(s_257), .O(gate240inter4));
  nand2 gate2344(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2345(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2346(.a(G263), .O(gate240inter7));
  inv1  gate2347(.a(G715), .O(gate240inter8));
  nand2 gate2348(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2349(.a(s_257), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2350(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2351(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2352(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1555(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1556(.a(gate244inter0), .b(s_144), .O(gate244inter1));
  and2  gate1557(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1558(.a(s_144), .O(gate244inter3));
  inv1  gate1559(.a(s_145), .O(gate244inter4));
  nand2 gate1560(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1561(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1562(.a(G721), .O(gate244inter7));
  inv1  gate1563(.a(G733), .O(gate244inter8));
  nand2 gate1564(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1565(.a(s_145), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1566(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1567(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1568(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1443(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1444(.a(gate247inter0), .b(s_128), .O(gate247inter1));
  and2  gate1445(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1446(.a(s_128), .O(gate247inter3));
  inv1  gate1447(.a(s_129), .O(gate247inter4));
  nand2 gate1448(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1449(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1450(.a(G251), .O(gate247inter7));
  inv1  gate1451(.a(G739), .O(gate247inter8));
  nand2 gate1452(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1453(.a(s_129), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1454(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1455(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1456(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2017(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2018(.a(gate248inter0), .b(s_210), .O(gate248inter1));
  and2  gate2019(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2020(.a(s_210), .O(gate248inter3));
  inv1  gate2021(.a(s_211), .O(gate248inter4));
  nand2 gate2022(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2023(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2024(.a(G727), .O(gate248inter7));
  inv1  gate2025(.a(G739), .O(gate248inter8));
  nand2 gate2026(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2027(.a(s_211), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2028(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2029(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2030(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1681(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1682(.a(gate250inter0), .b(s_162), .O(gate250inter1));
  and2  gate1683(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1684(.a(s_162), .O(gate250inter3));
  inv1  gate1685(.a(s_163), .O(gate250inter4));
  nand2 gate1686(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1687(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1688(.a(G706), .O(gate250inter7));
  inv1  gate1689(.a(G742), .O(gate250inter8));
  nand2 gate1690(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1691(.a(s_163), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1692(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1693(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1694(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2717(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2718(.a(gate252inter0), .b(s_310), .O(gate252inter1));
  and2  gate2719(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2720(.a(s_310), .O(gate252inter3));
  inv1  gate2721(.a(s_311), .O(gate252inter4));
  nand2 gate2722(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2723(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2724(.a(G709), .O(gate252inter7));
  inv1  gate2725(.a(G745), .O(gate252inter8));
  nand2 gate2726(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2727(.a(s_311), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2728(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2729(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2730(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2591(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2592(.a(gate255inter0), .b(s_292), .O(gate255inter1));
  and2  gate2593(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2594(.a(s_292), .O(gate255inter3));
  inv1  gate2595(.a(s_293), .O(gate255inter4));
  nand2 gate2596(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2597(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2598(.a(G263), .O(gate255inter7));
  inv1  gate2599(.a(G751), .O(gate255inter8));
  nand2 gate2600(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2601(.a(s_293), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2602(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2603(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2604(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2353(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2354(.a(gate257inter0), .b(s_258), .O(gate257inter1));
  and2  gate2355(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2356(.a(s_258), .O(gate257inter3));
  inv1  gate2357(.a(s_259), .O(gate257inter4));
  nand2 gate2358(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2359(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2360(.a(G754), .O(gate257inter7));
  inv1  gate2361(.a(G755), .O(gate257inter8));
  nand2 gate2362(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2363(.a(s_259), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2364(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2365(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2366(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1709(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1710(.a(gate258inter0), .b(s_166), .O(gate258inter1));
  and2  gate1711(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1712(.a(s_166), .O(gate258inter3));
  inv1  gate1713(.a(s_167), .O(gate258inter4));
  nand2 gate1714(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1715(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1716(.a(G756), .O(gate258inter7));
  inv1  gate1717(.a(G757), .O(gate258inter8));
  nand2 gate1718(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1719(.a(s_167), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1720(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1721(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1722(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1177(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1178(.a(gate261inter0), .b(s_90), .O(gate261inter1));
  and2  gate1179(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1180(.a(s_90), .O(gate261inter3));
  inv1  gate1181(.a(s_91), .O(gate261inter4));
  nand2 gate1182(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1183(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1184(.a(G762), .O(gate261inter7));
  inv1  gate1185(.a(G763), .O(gate261inter8));
  nand2 gate1186(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1187(.a(s_91), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1188(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1189(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1190(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2409(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2410(.a(gate265inter0), .b(s_266), .O(gate265inter1));
  and2  gate2411(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2412(.a(s_266), .O(gate265inter3));
  inv1  gate2413(.a(s_267), .O(gate265inter4));
  nand2 gate2414(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2415(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2416(.a(G642), .O(gate265inter7));
  inv1  gate2417(.a(G770), .O(gate265inter8));
  nand2 gate2418(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2419(.a(s_267), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2420(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2421(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2422(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1485(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1486(.a(gate268inter0), .b(s_134), .O(gate268inter1));
  and2  gate1487(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1488(.a(s_134), .O(gate268inter3));
  inv1  gate1489(.a(s_135), .O(gate268inter4));
  nand2 gate1490(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1491(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1492(.a(G651), .O(gate268inter7));
  inv1  gate1493(.a(G779), .O(gate268inter8));
  nand2 gate1494(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1495(.a(s_135), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1496(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1497(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1498(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2787(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2788(.a(gate274inter0), .b(s_320), .O(gate274inter1));
  and2  gate2789(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2790(.a(s_320), .O(gate274inter3));
  inv1  gate2791(.a(s_321), .O(gate274inter4));
  nand2 gate2792(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2793(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2794(.a(G770), .O(gate274inter7));
  inv1  gate2795(.a(G794), .O(gate274inter8));
  nand2 gate2796(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2797(.a(s_321), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2798(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2799(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2800(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1499(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1500(.a(gate277inter0), .b(s_136), .O(gate277inter1));
  and2  gate1501(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1502(.a(s_136), .O(gate277inter3));
  inv1  gate1503(.a(s_137), .O(gate277inter4));
  nand2 gate1504(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1505(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1506(.a(G648), .O(gate277inter7));
  inv1  gate1507(.a(G800), .O(gate277inter8));
  nand2 gate1508(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1509(.a(s_137), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1510(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1511(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1512(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate2171(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2172(.a(gate278inter0), .b(s_232), .O(gate278inter1));
  and2  gate2173(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2174(.a(s_232), .O(gate278inter3));
  inv1  gate2175(.a(s_233), .O(gate278inter4));
  nand2 gate2176(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2177(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2178(.a(G776), .O(gate278inter7));
  inv1  gate2179(.a(G800), .O(gate278inter8));
  nand2 gate2180(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2181(.a(s_233), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2182(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2183(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2184(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2521(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2522(.a(gate282inter0), .b(s_282), .O(gate282inter1));
  and2  gate2523(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2524(.a(s_282), .O(gate282inter3));
  inv1  gate2525(.a(s_283), .O(gate282inter4));
  nand2 gate2526(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2527(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2528(.a(G782), .O(gate282inter7));
  inv1  gate2529(.a(G806), .O(gate282inter8));
  nand2 gate2530(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2531(.a(s_283), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2532(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2533(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2534(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2185(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2186(.a(gate283inter0), .b(s_234), .O(gate283inter1));
  and2  gate2187(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2188(.a(s_234), .O(gate283inter3));
  inv1  gate2189(.a(s_235), .O(gate283inter4));
  nand2 gate2190(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2191(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2192(.a(G657), .O(gate283inter7));
  inv1  gate2193(.a(G809), .O(gate283inter8));
  nand2 gate2194(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2195(.a(s_235), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2196(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2197(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2198(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1821(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1822(.a(gate284inter0), .b(s_182), .O(gate284inter1));
  and2  gate1823(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1824(.a(s_182), .O(gate284inter3));
  inv1  gate1825(.a(s_183), .O(gate284inter4));
  nand2 gate1826(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1827(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1828(.a(G785), .O(gate284inter7));
  inv1  gate1829(.a(G809), .O(gate284inter8));
  nand2 gate1830(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1831(.a(s_183), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1832(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1833(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1834(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2647(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2648(.a(gate285inter0), .b(s_300), .O(gate285inter1));
  and2  gate2649(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2650(.a(s_300), .O(gate285inter3));
  inv1  gate2651(.a(s_301), .O(gate285inter4));
  nand2 gate2652(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2653(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2654(.a(G660), .O(gate285inter7));
  inv1  gate2655(.a(G812), .O(gate285inter8));
  nand2 gate2656(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2657(.a(s_301), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2658(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2659(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2660(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2745(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2746(.a(gate287inter0), .b(s_314), .O(gate287inter1));
  and2  gate2747(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2748(.a(s_314), .O(gate287inter3));
  inv1  gate2749(.a(s_315), .O(gate287inter4));
  nand2 gate2750(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2751(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2752(.a(G663), .O(gate287inter7));
  inv1  gate2753(.a(G815), .O(gate287inter8));
  nand2 gate2754(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2755(.a(s_315), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2756(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2757(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2758(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1261(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1262(.a(gate288inter0), .b(s_102), .O(gate288inter1));
  and2  gate1263(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1264(.a(s_102), .O(gate288inter3));
  inv1  gate1265(.a(s_103), .O(gate288inter4));
  nand2 gate1266(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1267(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1268(.a(G791), .O(gate288inter7));
  inv1  gate1269(.a(G815), .O(gate288inter8));
  nand2 gate1270(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1271(.a(s_103), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1272(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1273(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1274(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate841(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate842(.a(gate292inter0), .b(s_42), .O(gate292inter1));
  and2  gate843(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate844(.a(s_42), .O(gate292inter3));
  inv1  gate845(.a(s_43), .O(gate292inter4));
  nand2 gate846(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate847(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate848(.a(G824), .O(gate292inter7));
  inv1  gate849(.a(G825), .O(gate292inter8));
  nand2 gate850(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate851(.a(s_43), .b(gate292inter3), .O(gate292inter10));
  nor2  gate852(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate853(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate854(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2101(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2102(.a(gate296inter0), .b(s_222), .O(gate296inter1));
  and2  gate2103(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2104(.a(s_222), .O(gate296inter3));
  inv1  gate2105(.a(s_223), .O(gate296inter4));
  nand2 gate2106(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2107(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2108(.a(G826), .O(gate296inter7));
  inv1  gate2109(.a(G827), .O(gate296inter8));
  nand2 gate2110(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2111(.a(s_223), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2112(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2113(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2114(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate813(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate814(.a(gate391inter0), .b(s_38), .O(gate391inter1));
  and2  gate815(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate816(.a(s_38), .O(gate391inter3));
  inv1  gate817(.a(s_39), .O(gate391inter4));
  nand2 gate818(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate819(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate820(.a(G5), .O(gate391inter7));
  inv1  gate821(.a(G1048), .O(gate391inter8));
  nand2 gate822(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate823(.a(s_39), .b(gate391inter3), .O(gate391inter10));
  nor2  gate824(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate825(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate826(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1107(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1108(.a(gate394inter0), .b(s_80), .O(gate394inter1));
  and2  gate1109(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1110(.a(s_80), .O(gate394inter3));
  inv1  gate1111(.a(s_81), .O(gate394inter4));
  nand2 gate1112(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1113(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1114(.a(G8), .O(gate394inter7));
  inv1  gate1115(.a(G1057), .O(gate394inter8));
  nand2 gate1116(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1117(.a(s_81), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1118(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1119(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1120(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2269(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2270(.a(gate396inter0), .b(s_246), .O(gate396inter1));
  and2  gate2271(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2272(.a(s_246), .O(gate396inter3));
  inv1  gate2273(.a(s_247), .O(gate396inter4));
  nand2 gate2274(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2275(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2276(.a(G10), .O(gate396inter7));
  inv1  gate2277(.a(G1063), .O(gate396inter8));
  nand2 gate2278(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2279(.a(s_247), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2280(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2281(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2282(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2199(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2200(.a(gate400inter0), .b(s_236), .O(gate400inter1));
  and2  gate2201(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2202(.a(s_236), .O(gate400inter3));
  inv1  gate2203(.a(s_237), .O(gate400inter4));
  nand2 gate2204(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2205(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2206(.a(G14), .O(gate400inter7));
  inv1  gate2207(.a(G1075), .O(gate400inter8));
  nand2 gate2208(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2209(.a(s_237), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2210(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2211(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2212(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1989(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1990(.a(gate402inter0), .b(s_206), .O(gate402inter1));
  and2  gate1991(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1992(.a(s_206), .O(gate402inter3));
  inv1  gate1993(.a(s_207), .O(gate402inter4));
  nand2 gate1994(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1995(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1996(.a(G16), .O(gate402inter7));
  inv1  gate1997(.a(G1081), .O(gate402inter8));
  nand2 gate1998(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1999(.a(s_207), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2000(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2001(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2002(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1331(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1332(.a(gate408inter0), .b(s_112), .O(gate408inter1));
  and2  gate1333(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1334(.a(s_112), .O(gate408inter3));
  inv1  gate1335(.a(s_113), .O(gate408inter4));
  nand2 gate1336(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1337(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1338(.a(G22), .O(gate408inter7));
  inv1  gate1339(.a(G1099), .O(gate408inter8));
  nand2 gate1340(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1341(.a(s_113), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1342(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1343(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1344(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1275(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1276(.a(gate409inter0), .b(s_104), .O(gate409inter1));
  and2  gate1277(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1278(.a(s_104), .O(gate409inter3));
  inv1  gate1279(.a(s_105), .O(gate409inter4));
  nand2 gate1280(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1281(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1282(.a(G23), .O(gate409inter7));
  inv1  gate1283(.a(G1102), .O(gate409inter8));
  nand2 gate1284(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1285(.a(s_105), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1286(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1287(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1288(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1065(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1066(.a(gate410inter0), .b(s_74), .O(gate410inter1));
  and2  gate1067(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1068(.a(s_74), .O(gate410inter3));
  inv1  gate1069(.a(s_75), .O(gate410inter4));
  nand2 gate1070(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1071(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1072(.a(G24), .O(gate410inter7));
  inv1  gate1073(.a(G1105), .O(gate410inter8));
  nand2 gate1074(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1075(.a(s_75), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1076(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1077(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1078(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2241(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2242(.a(gate412inter0), .b(s_242), .O(gate412inter1));
  and2  gate2243(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2244(.a(s_242), .O(gate412inter3));
  inv1  gate2245(.a(s_243), .O(gate412inter4));
  nand2 gate2246(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2247(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2248(.a(G26), .O(gate412inter7));
  inv1  gate2249(.a(G1111), .O(gate412inter8));
  nand2 gate2250(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2251(.a(s_243), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2252(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2253(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2254(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1303(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1304(.a(gate414inter0), .b(s_108), .O(gate414inter1));
  and2  gate1305(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1306(.a(s_108), .O(gate414inter3));
  inv1  gate1307(.a(s_109), .O(gate414inter4));
  nand2 gate1308(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1309(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1310(.a(G28), .O(gate414inter7));
  inv1  gate1311(.a(G1117), .O(gate414inter8));
  nand2 gate1312(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1313(.a(s_109), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1314(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1315(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1316(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate981(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate982(.a(gate415inter0), .b(s_62), .O(gate415inter1));
  and2  gate983(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate984(.a(s_62), .O(gate415inter3));
  inv1  gate985(.a(s_63), .O(gate415inter4));
  nand2 gate986(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate987(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate988(.a(G29), .O(gate415inter7));
  inv1  gate989(.a(G1120), .O(gate415inter8));
  nand2 gate990(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate991(.a(s_63), .b(gate415inter3), .O(gate415inter10));
  nor2  gate992(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate993(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate994(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate2451(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2452(.a(gate416inter0), .b(s_272), .O(gate416inter1));
  and2  gate2453(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2454(.a(s_272), .O(gate416inter3));
  inv1  gate2455(.a(s_273), .O(gate416inter4));
  nand2 gate2456(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2457(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2458(.a(G30), .O(gate416inter7));
  inv1  gate2459(.a(G1123), .O(gate416inter8));
  nand2 gate2460(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2461(.a(s_273), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2462(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2463(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2464(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1359(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1360(.a(gate417inter0), .b(s_116), .O(gate417inter1));
  and2  gate1361(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1362(.a(s_116), .O(gate417inter3));
  inv1  gate1363(.a(s_117), .O(gate417inter4));
  nand2 gate1364(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1365(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1366(.a(G31), .O(gate417inter7));
  inv1  gate1367(.a(G1126), .O(gate417inter8));
  nand2 gate1368(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1369(.a(s_117), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1370(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1371(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1372(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1191(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1192(.a(gate420inter0), .b(s_92), .O(gate420inter1));
  and2  gate1193(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1194(.a(s_92), .O(gate420inter3));
  inv1  gate1195(.a(s_93), .O(gate420inter4));
  nand2 gate1196(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1197(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1198(.a(G1036), .O(gate420inter7));
  inv1  gate1199(.a(G1132), .O(gate420inter8));
  nand2 gate1200(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1201(.a(s_93), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1202(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1203(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1204(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2381(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2382(.a(gate422inter0), .b(s_262), .O(gate422inter1));
  and2  gate2383(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2384(.a(s_262), .O(gate422inter3));
  inv1  gate2385(.a(s_263), .O(gate422inter4));
  nand2 gate2386(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2387(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2388(.a(G1039), .O(gate422inter7));
  inv1  gate2389(.a(G1135), .O(gate422inter8));
  nand2 gate2390(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2391(.a(s_263), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2392(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2393(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2394(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1051(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1052(.a(gate424inter0), .b(s_72), .O(gate424inter1));
  and2  gate1053(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1054(.a(s_72), .O(gate424inter3));
  inv1  gate1055(.a(s_73), .O(gate424inter4));
  nand2 gate1056(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1057(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1058(.a(G1042), .O(gate424inter7));
  inv1  gate1059(.a(G1138), .O(gate424inter8));
  nand2 gate1060(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1061(.a(s_73), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1062(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1063(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1064(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate617(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate618(.a(gate426inter0), .b(s_10), .O(gate426inter1));
  and2  gate619(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate620(.a(s_10), .O(gate426inter3));
  inv1  gate621(.a(s_11), .O(gate426inter4));
  nand2 gate622(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate623(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate624(.a(G1045), .O(gate426inter7));
  inv1  gate625(.a(G1141), .O(gate426inter8));
  nand2 gate626(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate627(.a(s_11), .b(gate426inter3), .O(gate426inter10));
  nor2  gate628(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate629(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate630(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1891(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1892(.a(gate430inter0), .b(s_192), .O(gate430inter1));
  and2  gate1893(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1894(.a(s_192), .O(gate430inter3));
  inv1  gate1895(.a(s_193), .O(gate430inter4));
  nand2 gate1896(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1897(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1898(.a(G1051), .O(gate430inter7));
  inv1  gate1899(.a(G1147), .O(gate430inter8));
  nand2 gate1900(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1901(.a(s_193), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1902(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1903(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1904(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate729(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate730(.a(gate439inter0), .b(s_26), .O(gate439inter1));
  and2  gate731(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate732(.a(s_26), .O(gate439inter3));
  inv1  gate733(.a(s_27), .O(gate439inter4));
  nand2 gate734(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate735(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate736(.a(G11), .O(gate439inter7));
  inv1  gate737(.a(G1162), .O(gate439inter8));
  nand2 gate738(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate739(.a(s_27), .b(gate439inter3), .O(gate439inter10));
  nor2  gate740(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate741(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate742(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1009(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1010(.a(gate441inter0), .b(s_66), .O(gate441inter1));
  and2  gate1011(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1012(.a(s_66), .O(gate441inter3));
  inv1  gate1013(.a(s_67), .O(gate441inter4));
  nand2 gate1014(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1015(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1016(.a(G12), .O(gate441inter7));
  inv1  gate1017(.a(G1165), .O(gate441inter8));
  nand2 gate1018(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1019(.a(s_67), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1020(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1021(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1022(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1723(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1724(.a(gate442inter0), .b(s_168), .O(gate442inter1));
  and2  gate1725(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1726(.a(s_168), .O(gate442inter3));
  inv1  gate1727(.a(s_169), .O(gate442inter4));
  nand2 gate1728(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1729(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1730(.a(G1069), .O(gate442inter7));
  inv1  gate1731(.a(G1165), .O(gate442inter8));
  nand2 gate1732(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1733(.a(s_169), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1734(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1735(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1736(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate911(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate912(.a(gate443inter0), .b(s_52), .O(gate443inter1));
  and2  gate913(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate914(.a(s_52), .O(gate443inter3));
  inv1  gate915(.a(s_53), .O(gate443inter4));
  nand2 gate916(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate917(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate918(.a(G13), .O(gate443inter7));
  inv1  gate919(.a(G1168), .O(gate443inter8));
  nand2 gate920(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate921(.a(s_53), .b(gate443inter3), .O(gate443inter10));
  nor2  gate922(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate923(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate924(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate2115(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2116(.a(gate446inter0), .b(s_224), .O(gate446inter1));
  and2  gate2117(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2118(.a(s_224), .O(gate446inter3));
  inv1  gate2119(.a(s_225), .O(gate446inter4));
  nand2 gate2120(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2121(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2122(.a(G1075), .O(gate446inter7));
  inv1  gate2123(.a(G1171), .O(gate446inter8));
  nand2 gate2124(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2125(.a(s_225), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2126(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2127(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2128(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1611(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1612(.a(gate448inter0), .b(s_152), .O(gate448inter1));
  and2  gate1613(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1614(.a(s_152), .O(gate448inter3));
  inv1  gate1615(.a(s_153), .O(gate448inter4));
  nand2 gate1616(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1617(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1618(.a(G1078), .O(gate448inter7));
  inv1  gate1619(.a(G1174), .O(gate448inter8));
  nand2 gate1620(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1621(.a(s_153), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1622(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1623(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1624(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1625(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1626(.a(gate451inter0), .b(s_154), .O(gate451inter1));
  and2  gate1627(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1628(.a(s_154), .O(gate451inter3));
  inv1  gate1629(.a(s_155), .O(gate451inter4));
  nand2 gate1630(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1631(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1632(.a(G17), .O(gate451inter7));
  inv1  gate1633(.a(G1180), .O(gate451inter8));
  nand2 gate1634(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1635(.a(s_155), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1636(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1637(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1638(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1205(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1206(.a(gate452inter0), .b(s_94), .O(gate452inter1));
  and2  gate1207(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1208(.a(s_94), .O(gate452inter3));
  inv1  gate1209(.a(s_95), .O(gate452inter4));
  nand2 gate1210(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1211(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1212(.a(G1084), .O(gate452inter7));
  inv1  gate1213(.a(G1180), .O(gate452inter8));
  nand2 gate1214(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1215(.a(s_95), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1216(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1217(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1218(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2577(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2578(.a(gate455inter0), .b(s_290), .O(gate455inter1));
  and2  gate2579(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2580(.a(s_290), .O(gate455inter3));
  inv1  gate2581(.a(s_291), .O(gate455inter4));
  nand2 gate2582(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2583(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2584(.a(G19), .O(gate455inter7));
  inv1  gate2585(.a(G1186), .O(gate455inter8));
  nand2 gate2586(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2587(.a(s_291), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2588(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2589(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2590(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2367(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2368(.a(gate459inter0), .b(s_260), .O(gate459inter1));
  and2  gate2369(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2370(.a(s_260), .O(gate459inter3));
  inv1  gate2371(.a(s_261), .O(gate459inter4));
  nand2 gate2372(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2373(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2374(.a(G21), .O(gate459inter7));
  inv1  gate2375(.a(G1192), .O(gate459inter8));
  nand2 gate2376(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2377(.a(s_261), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2378(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2379(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2380(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1583(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1584(.a(gate460inter0), .b(s_148), .O(gate460inter1));
  and2  gate1585(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1586(.a(s_148), .O(gate460inter3));
  inv1  gate1587(.a(s_149), .O(gate460inter4));
  nand2 gate1588(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1589(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1590(.a(G1096), .O(gate460inter7));
  inv1  gate1591(.a(G1192), .O(gate460inter8));
  nand2 gate1592(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1593(.a(s_149), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1594(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1595(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1596(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2493(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2494(.a(gate465inter0), .b(s_278), .O(gate465inter1));
  and2  gate2495(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2496(.a(s_278), .O(gate465inter3));
  inv1  gate2497(.a(s_279), .O(gate465inter4));
  nand2 gate2498(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2499(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2500(.a(G24), .O(gate465inter7));
  inv1  gate2501(.a(G1201), .O(gate465inter8));
  nand2 gate2502(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2503(.a(s_279), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2504(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2505(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2506(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2423(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2424(.a(gate466inter0), .b(s_268), .O(gate466inter1));
  and2  gate2425(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2426(.a(s_268), .O(gate466inter3));
  inv1  gate2427(.a(s_269), .O(gate466inter4));
  nand2 gate2428(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2429(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2430(.a(G1105), .O(gate466inter7));
  inv1  gate2431(.a(G1201), .O(gate466inter8));
  nand2 gate2432(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2433(.a(s_269), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2434(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2435(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2436(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate883(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate884(.a(gate468inter0), .b(s_48), .O(gate468inter1));
  and2  gate885(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate886(.a(s_48), .O(gate468inter3));
  inv1  gate887(.a(s_49), .O(gate468inter4));
  nand2 gate888(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate889(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate890(.a(G1108), .O(gate468inter7));
  inv1  gate891(.a(G1204), .O(gate468inter8));
  nand2 gate892(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate893(.a(s_49), .b(gate468inter3), .O(gate468inter10));
  nor2  gate894(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate895(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate896(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1219(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1220(.a(gate471inter0), .b(s_96), .O(gate471inter1));
  and2  gate1221(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1222(.a(s_96), .O(gate471inter3));
  inv1  gate1223(.a(s_97), .O(gate471inter4));
  nand2 gate1224(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1225(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1226(.a(G27), .O(gate471inter7));
  inv1  gate1227(.a(G1210), .O(gate471inter8));
  nand2 gate1228(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1229(.a(s_97), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1230(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1231(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1232(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate953(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate954(.a(gate472inter0), .b(s_58), .O(gate472inter1));
  and2  gate955(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate956(.a(s_58), .O(gate472inter3));
  inv1  gate957(.a(s_59), .O(gate472inter4));
  nand2 gate958(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate959(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate960(.a(G1114), .O(gate472inter7));
  inv1  gate961(.a(G1210), .O(gate472inter8));
  nand2 gate962(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate963(.a(s_59), .b(gate472inter3), .O(gate472inter10));
  nor2  gate964(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate965(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate966(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1037(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1038(.a(gate475inter0), .b(s_70), .O(gate475inter1));
  and2  gate1039(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1040(.a(s_70), .O(gate475inter3));
  inv1  gate1041(.a(s_71), .O(gate475inter4));
  nand2 gate1042(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1043(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1044(.a(G29), .O(gate475inter7));
  inv1  gate1045(.a(G1216), .O(gate475inter8));
  nand2 gate1046(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1047(.a(s_71), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1048(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1049(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1050(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate827(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate828(.a(gate476inter0), .b(s_40), .O(gate476inter1));
  and2  gate829(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate830(.a(s_40), .O(gate476inter3));
  inv1  gate831(.a(s_41), .O(gate476inter4));
  nand2 gate832(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate833(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate834(.a(G1120), .O(gate476inter7));
  inv1  gate835(.a(G1216), .O(gate476inter8));
  nand2 gate836(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate837(.a(s_41), .b(gate476inter3), .O(gate476inter10));
  nor2  gate838(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate839(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate840(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1905(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1906(.a(gate477inter0), .b(s_194), .O(gate477inter1));
  and2  gate1907(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1908(.a(s_194), .O(gate477inter3));
  inv1  gate1909(.a(s_195), .O(gate477inter4));
  nand2 gate1910(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1911(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1912(.a(G30), .O(gate477inter7));
  inv1  gate1913(.a(G1219), .O(gate477inter8));
  nand2 gate1914(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1915(.a(s_195), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1916(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1917(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1918(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate687(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate688(.a(gate480inter0), .b(s_20), .O(gate480inter1));
  and2  gate689(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate690(.a(s_20), .O(gate480inter3));
  inv1  gate691(.a(s_21), .O(gate480inter4));
  nand2 gate692(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate693(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate694(.a(G1126), .O(gate480inter7));
  inv1  gate695(.a(G1222), .O(gate480inter8));
  nand2 gate696(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate697(.a(s_21), .b(gate480inter3), .O(gate480inter10));
  nor2  gate698(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate699(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate700(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1093(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1094(.a(gate486inter0), .b(s_78), .O(gate486inter1));
  and2  gate1095(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1096(.a(s_78), .O(gate486inter3));
  inv1  gate1097(.a(s_79), .O(gate486inter4));
  nand2 gate1098(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1099(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1100(.a(G1234), .O(gate486inter7));
  inv1  gate1101(.a(G1235), .O(gate486inter8));
  nand2 gate1102(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1103(.a(s_79), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1104(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1105(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1106(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2633(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2634(.a(gate487inter0), .b(s_298), .O(gate487inter1));
  and2  gate2635(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2636(.a(s_298), .O(gate487inter3));
  inv1  gate2637(.a(s_299), .O(gate487inter4));
  nand2 gate2638(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2639(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2640(.a(G1236), .O(gate487inter7));
  inv1  gate2641(.a(G1237), .O(gate487inter8));
  nand2 gate2642(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2643(.a(s_299), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2644(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2645(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2646(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate743(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate744(.a(gate488inter0), .b(s_28), .O(gate488inter1));
  and2  gate745(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate746(.a(s_28), .O(gate488inter3));
  inv1  gate747(.a(s_29), .O(gate488inter4));
  nand2 gate748(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate749(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate750(.a(G1238), .O(gate488inter7));
  inv1  gate751(.a(G1239), .O(gate488inter8));
  nand2 gate752(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate753(.a(s_29), .b(gate488inter3), .O(gate488inter10));
  nor2  gate754(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate755(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate756(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2689(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2690(.a(gate490inter0), .b(s_306), .O(gate490inter1));
  and2  gate2691(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2692(.a(s_306), .O(gate490inter3));
  inv1  gate2693(.a(s_307), .O(gate490inter4));
  nand2 gate2694(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2695(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2696(.a(G1242), .O(gate490inter7));
  inv1  gate2697(.a(G1243), .O(gate490inter8));
  nand2 gate2698(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2699(.a(s_307), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2700(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2701(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2702(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2143(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2144(.a(gate492inter0), .b(s_228), .O(gate492inter1));
  and2  gate2145(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2146(.a(s_228), .O(gate492inter3));
  inv1  gate2147(.a(s_229), .O(gate492inter4));
  nand2 gate2148(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2149(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2150(.a(G1246), .O(gate492inter7));
  inv1  gate2151(.a(G1247), .O(gate492inter8));
  nand2 gate2152(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2153(.a(s_229), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2154(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2155(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2156(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate701(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate702(.a(gate493inter0), .b(s_22), .O(gate493inter1));
  and2  gate703(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate704(.a(s_22), .O(gate493inter3));
  inv1  gate705(.a(s_23), .O(gate493inter4));
  nand2 gate706(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate707(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate708(.a(G1248), .O(gate493inter7));
  inv1  gate709(.a(G1249), .O(gate493inter8));
  nand2 gate710(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate711(.a(s_23), .b(gate493inter3), .O(gate493inter10));
  nor2  gate712(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate713(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate714(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate589(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate590(.a(gate496inter0), .b(s_6), .O(gate496inter1));
  and2  gate591(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate592(.a(s_6), .O(gate496inter3));
  inv1  gate593(.a(s_7), .O(gate496inter4));
  nand2 gate594(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate595(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate596(.a(G1254), .O(gate496inter7));
  inv1  gate597(.a(G1255), .O(gate496inter8));
  nand2 gate598(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate599(.a(s_7), .b(gate496inter3), .O(gate496inter10));
  nor2  gate600(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate601(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate602(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate2479(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2480(.a(gate497inter0), .b(s_276), .O(gate497inter1));
  and2  gate2481(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2482(.a(s_276), .O(gate497inter3));
  inv1  gate2483(.a(s_277), .O(gate497inter4));
  nand2 gate2484(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2485(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2486(.a(G1256), .O(gate497inter7));
  inv1  gate2487(.a(G1257), .O(gate497inter8));
  nand2 gate2488(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2489(.a(s_277), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2490(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2491(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2492(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate799(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate800(.a(gate498inter0), .b(s_36), .O(gate498inter1));
  and2  gate801(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate802(.a(s_36), .O(gate498inter3));
  inv1  gate803(.a(s_37), .O(gate498inter4));
  nand2 gate804(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate805(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate806(.a(G1258), .O(gate498inter7));
  inv1  gate807(.a(G1259), .O(gate498inter8));
  nand2 gate808(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate809(.a(s_37), .b(gate498inter3), .O(gate498inter10));
  nor2  gate810(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate811(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate812(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1835(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1836(.a(gate499inter0), .b(s_184), .O(gate499inter1));
  and2  gate1837(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1838(.a(s_184), .O(gate499inter3));
  inv1  gate1839(.a(s_185), .O(gate499inter4));
  nand2 gate1840(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1841(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1842(.a(G1260), .O(gate499inter7));
  inv1  gate1843(.a(G1261), .O(gate499inter8));
  nand2 gate1844(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1845(.a(s_185), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1846(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1847(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1848(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2045(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2046(.a(gate500inter0), .b(s_214), .O(gate500inter1));
  and2  gate2047(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2048(.a(s_214), .O(gate500inter3));
  inv1  gate2049(.a(s_215), .O(gate500inter4));
  nand2 gate2050(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2051(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2052(.a(G1262), .O(gate500inter7));
  inv1  gate2053(.a(G1263), .O(gate500inter8));
  nand2 gate2054(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2055(.a(s_215), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2056(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2057(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2058(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate897(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate898(.a(gate501inter0), .b(s_50), .O(gate501inter1));
  and2  gate899(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate900(.a(s_50), .O(gate501inter3));
  inv1  gate901(.a(s_51), .O(gate501inter4));
  nand2 gate902(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate903(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate904(.a(G1264), .O(gate501inter7));
  inv1  gate905(.a(G1265), .O(gate501inter8));
  nand2 gate906(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate907(.a(s_51), .b(gate501inter3), .O(gate501inter10));
  nor2  gate908(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate909(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate910(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2003(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2004(.a(gate503inter0), .b(s_208), .O(gate503inter1));
  and2  gate2005(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2006(.a(s_208), .O(gate503inter3));
  inv1  gate2007(.a(s_209), .O(gate503inter4));
  nand2 gate2008(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2009(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2010(.a(G1268), .O(gate503inter7));
  inv1  gate2011(.a(G1269), .O(gate503inter8));
  nand2 gate2012(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2013(.a(s_209), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2014(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2015(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2016(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1541(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1542(.a(gate507inter0), .b(s_142), .O(gate507inter1));
  and2  gate1543(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1544(.a(s_142), .O(gate507inter3));
  inv1  gate1545(.a(s_143), .O(gate507inter4));
  nand2 gate1546(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1547(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1548(.a(G1276), .O(gate507inter7));
  inv1  gate1549(.a(G1277), .O(gate507inter8));
  nand2 gate1550(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1551(.a(s_143), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1552(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1553(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1554(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2661(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2662(.a(gate511inter0), .b(s_302), .O(gate511inter1));
  and2  gate2663(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2664(.a(s_302), .O(gate511inter3));
  inv1  gate2665(.a(s_303), .O(gate511inter4));
  nand2 gate2666(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2667(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2668(.a(G1284), .O(gate511inter7));
  inv1  gate2669(.a(G1285), .O(gate511inter8));
  nand2 gate2670(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2671(.a(s_303), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2672(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2673(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2674(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1415(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1416(.a(gate513inter0), .b(s_124), .O(gate513inter1));
  and2  gate1417(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1418(.a(s_124), .O(gate513inter3));
  inv1  gate1419(.a(s_125), .O(gate513inter4));
  nand2 gate1420(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1421(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1422(.a(G1288), .O(gate513inter7));
  inv1  gate1423(.a(G1289), .O(gate513inter8));
  nand2 gate1424(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1425(.a(s_125), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1426(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1427(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1428(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule