module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate631(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate632(.a(gate14inter0), .b(s_12), .O(gate14inter1));
  and2  gate633(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate634(.a(s_12), .O(gate14inter3));
  inv1  gate635(.a(s_13), .O(gate14inter4));
  nand2 gate636(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate637(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate638(.a(G11), .O(gate14inter7));
  inv1  gate639(.a(G12), .O(gate14inter8));
  nand2 gate640(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate641(.a(s_13), .b(gate14inter3), .O(gate14inter10));
  nor2  gate642(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate643(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate644(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate911(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate912(.a(gate19inter0), .b(s_52), .O(gate19inter1));
  and2  gate913(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate914(.a(s_52), .O(gate19inter3));
  inv1  gate915(.a(s_53), .O(gate19inter4));
  nand2 gate916(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate917(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate918(.a(G21), .O(gate19inter7));
  inv1  gate919(.a(G22), .O(gate19inter8));
  nand2 gate920(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate921(.a(s_53), .b(gate19inter3), .O(gate19inter10));
  nor2  gate922(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate923(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate924(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1737(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1738(.a(gate20inter0), .b(s_170), .O(gate20inter1));
  and2  gate1739(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1740(.a(s_170), .O(gate20inter3));
  inv1  gate1741(.a(s_171), .O(gate20inter4));
  nand2 gate1742(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1743(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1744(.a(G23), .O(gate20inter7));
  inv1  gate1745(.a(G24), .O(gate20inter8));
  nand2 gate1746(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1747(.a(s_171), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1748(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1749(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1750(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1401(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1402(.a(gate22inter0), .b(s_122), .O(gate22inter1));
  and2  gate1403(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1404(.a(s_122), .O(gate22inter3));
  inv1  gate1405(.a(s_123), .O(gate22inter4));
  nand2 gate1406(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1407(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1408(.a(G27), .O(gate22inter7));
  inv1  gate1409(.a(G28), .O(gate22inter8));
  nand2 gate1410(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1411(.a(s_123), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1412(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1413(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1414(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate995(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate996(.a(gate23inter0), .b(s_64), .O(gate23inter1));
  and2  gate997(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate998(.a(s_64), .O(gate23inter3));
  inv1  gate999(.a(s_65), .O(gate23inter4));
  nand2 gate1000(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1001(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1002(.a(G29), .O(gate23inter7));
  inv1  gate1003(.a(G30), .O(gate23inter8));
  nand2 gate1004(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1005(.a(s_65), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1006(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1007(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1008(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1359(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1360(.a(gate27inter0), .b(s_116), .O(gate27inter1));
  and2  gate1361(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1362(.a(s_116), .O(gate27inter3));
  inv1  gate1363(.a(s_117), .O(gate27inter4));
  nand2 gate1364(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1365(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1366(.a(G2), .O(gate27inter7));
  inv1  gate1367(.a(G6), .O(gate27inter8));
  nand2 gate1368(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1369(.a(s_117), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1370(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1371(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1372(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1065(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1066(.a(gate31inter0), .b(s_74), .O(gate31inter1));
  and2  gate1067(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1068(.a(s_74), .O(gate31inter3));
  inv1  gate1069(.a(s_75), .O(gate31inter4));
  nand2 gate1070(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1071(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1072(.a(G4), .O(gate31inter7));
  inv1  gate1073(.a(G8), .O(gate31inter8));
  nand2 gate1074(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1075(.a(s_75), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1076(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1077(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1078(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate673(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate674(.a(gate32inter0), .b(s_18), .O(gate32inter1));
  and2  gate675(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate676(.a(s_18), .O(gate32inter3));
  inv1  gate677(.a(s_19), .O(gate32inter4));
  nand2 gate678(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate679(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate680(.a(G12), .O(gate32inter7));
  inv1  gate681(.a(G16), .O(gate32inter8));
  nand2 gate682(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate683(.a(s_19), .b(gate32inter3), .O(gate32inter10));
  nor2  gate684(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate685(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate686(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate785(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate786(.a(gate33inter0), .b(s_34), .O(gate33inter1));
  and2  gate787(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate788(.a(s_34), .O(gate33inter3));
  inv1  gate789(.a(s_35), .O(gate33inter4));
  nand2 gate790(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate791(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate792(.a(G17), .O(gate33inter7));
  inv1  gate793(.a(G21), .O(gate33inter8));
  nand2 gate794(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate795(.a(s_35), .b(gate33inter3), .O(gate33inter10));
  nor2  gate796(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate797(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate798(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1457(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1458(.a(gate40inter0), .b(s_130), .O(gate40inter1));
  and2  gate1459(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1460(.a(s_130), .O(gate40inter3));
  inv1  gate1461(.a(s_131), .O(gate40inter4));
  nand2 gate1462(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1463(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1464(.a(G28), .O(gate40inter7));
  inv1  gate1465(.a(G32), .O(gate40inter8));
  nand2 gate1466(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1467(.a(s_131), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1468(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1469(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1470(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1723(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1724(.a(gate48inter0), .b(s_168), .O(gate48inter1));
  and2  gate1725(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1726(.a(s_168), .O(gate48inter3));
  inv1  gate1727(.a(s_169), .O(gate48inter4));
  nand2 gate1728(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1729(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1730(.a(G8), .O(gate48inter7));
  inv1  gate1731(.a(G275), .O(gate48inter8));
  nand2 gate1732(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1733(.a(s_169), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1734(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1735(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1736(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate575(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate576(.a(gate52inter0), .b(s_4), .O(gate52inter1));
  and2  gate577(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate578(.a(s_4), .O(gate52inter3));
  inv1  gate579(.a(s_5), .O(gate52inter4));
  nand2 gate580(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate581(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate582(.a(G12), .O(gate52inter7));
  inv1  gate583(.a(G281), .O(gate52inter8));
  nand2 gate584(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate585(.a(s_5), .b(gate52inter3), .O(gate52inter10));
  nor2  gate586(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate587(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate588(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate883(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate884(.a(gate71inter0), .b(s_48), .O(gate71inter1));
  and2  gate885(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate886(.a(s_48), .O(gate71inter3));
  inv1  gate887(.a(s_49), .O(gate71inter4));
  nand2 gate888(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate889(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate890(.a(G31), .O(gate71inter7));
  inv1  gate891(.a(G311), .O(gate71inter8));
  nand2 gate892(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate893(.a(s_49), .b(gate71inter3), .O(gate71inter10));
  nor2  gate894(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate895(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate896(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1681(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1682(.a(gate72inter0), .b(s_162), .O(gate72inter1));
  and2  gate1683(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1684(.a(s_162), .O(gate72inter3));
  inv1  gate1685(.a(s_163), .O(gate72inter4));
  nand2 gate1686(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1687(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1688(.a(G32), .O(gate72inter7));
  inv1  gate1689(.a(G311), .O(gate72inter8));
  nand2 gate1690(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1691(.a(s_163), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1692(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1693(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1694(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate827(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate828(.a(gate92inter0), .b(s_40), .O(gate92inter1));
  and2  gate829(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate830(.a(s_40), .O(gate92inter3));
  inv1  gate831(.a(s_41), .O(gate92inter4));
  nand2 gate832(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate833(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate834(.a(G29), .O(gate92inter7));
  inv1  gate835(.a(G341), .O(gate92inter8));
  nand2 gate836(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate837(.a(s_41), .b(gate92inter3), .O(gate92inter10));
  nor2  gate838(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate839(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate840(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1303(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1304(.a(gate100inter0), .b(s_108), .O(gate100inter1));
  and2  gate1305(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1306(.a(s_108), .O(gate100inter3));
  inv1  gate1307(.a(s_109), .O(gate100inter4));
  nand2 gate1308(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1309(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1310(.a(G31), .O(gate100inter7));
  inv1  gate1311(.a(G353), .O(gate100inter8));
  nand2 gate1312(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1313(.a(s_109), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1314(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1315(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1316(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1051(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1052(.a(gate115inter0), .b(s_72), .O(gate115inter1));
  and2  gate1053(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1054(.a(s_72), .O(gate115inter3));
  inv1  gate1055(.a(s_73), .O(gate115inter4));
  nand2 gate1056(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1057(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1058(.a(G382), .O(gate115inter7));
  inv1  gate1059(.a(G383), .O(gate115inter8));
  nand2 gate1060(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1061(.a(s_73), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1062(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1063(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1064(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate855(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate856(.a(gate117inter0), .b(s_44), .O(gate117inter1));
  and2  gate857(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate858(.a(s_44), .O(gate117inter3));
  inv1  gate859(.a(s_45), .O(gate117inter4));
  nand2 gate860(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate861(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate862(.a(G386), .O(gate117inter7));
  inv1  gate863(.a(G387), .O(gate117inter8));
  nand2 gate864(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate865(.a(s_45), .b(gate117inter3), .O(gate117inter10));
  nor2  gate866(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate867(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate868(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1583(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1584(.a(gate120inter0), .b(s_148), .O(gate120inter1));
  and2  gate1585(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1586(.a(s_148), .O(gate120inter3));
  inv1  gate1587(.a(s_149), .O(gate120inter4));
  nand2 gate1588(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1589(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1590(.a(G392), .O(gate120inter7));
  inv1  gate1591(.a(G393), .O(gate120inter8));
  nand2 gate1592(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1593(.a(s_149), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1594(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1595(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1596(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1093(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1094(.a(gate128inter0), .b(s_78), .O(gate128inter1));
  and2  gate1095(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1096(.a(s_78), .O(gate128inter3));
  inv1  gate1097(.a(s_79), .O(gate128inter4));
  nand2 gate1098(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1099(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1100(.a(G408), .O(gate128inter7));
  inv1  gate1101(.a(G409), .O(gate128inter8));
  nand2 gate1102(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1103(.a(s_79), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1104(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1105(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1106(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1695(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1696(.a(gate138inter0), .b(s_164), .O(gate138inter1));
  and2  gate1697(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1698(.a(s_164), .O(gate138inter3));
  inv1  gate1699(.a(s_165), .O(gate138inter4));
  nand2 gate1700(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1701(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1702(.a(G432), .O(gate138inter7));
  inv1  gate1703(.a(G435), .O(gate138inter8));
  nand2 gate1704(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1705(.a(s_165), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1706(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1707(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1708(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1233(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1234(.a(gate146inter0), .b(s_98), .O(gate146inter1));
  and2  gate1235(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1236(.a(s_98), .O(gate146inter3));
  inv1  gate1237(.a(s_99), .O(gate146inter4));
  nand2 gate1238(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1239(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1240(.a(G480), .O(gate146inter7));
  inv1  gate1241(.a(G483), .O(gate146inter8));
  nand2 gate1242(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1243(.a(s_99), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1244(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1245(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1246(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate617(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate618(.a(gate147inter0), .b(s_10), .O(gate147inter1));
  and2  gate619(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate620(.a(s_10), .O(gate147inter3));
  inv1  gate621(.a(s_11), .O(gate147inter4));
  nand2 gate622(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate623(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate624(.a(G486), .O(gate147inter7));
  inv1  gate625(.a(G489), .O(gate147inter8));
  nand2 gate626(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate627(.a(s_11), .b(gate147inter3), .O(gate147inter10));
  nor2  gate628(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate629(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate630(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1611(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1612(.a(gate151inter0), .b(s_152), .O(gate151inter1));
  and2  gate1613(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1614(.a(s_152), .O(gate151inter3));
  inv1  gate1615(.a(s_153), .O(gate151inter4));
  nand2 gate1616(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1617(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1618(.a(G510), .O(gate151inter7));
  inv1  gate1619(.a(G513), .O(gate151inter8));
  nand2 gate1620(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1621(.a(s_153), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1622(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1623(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1624(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate813(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate814(.a(gate154inter0), .b(s_38), .O(gate154inter1));
  and2  gate815(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate816(.a(s_38), .O(gate154inter3));
  inv1  gate817(.a(s_39), .O(gate154inter4));
  nand2 gate818(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate819(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate820(.a(G429), .O(gate154inter7));
  inv1  gate821(.a(G522), .O(gate154inter8));
  nand2 gate822(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate823(.a(s_39), .b(gate154inter3), .O(gate154inter10));
  nor2  gate824(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate825(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate826(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1107(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1108(.a(gate155inter0), .b(s_80), .O(gate155inter1));
  and2  gate1109(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1110(.a(s_80), .O(gate155inter3));
  inv1  gate1111(.a(s_81), .O(gate155inter4));
  nand2 gate1112(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1113(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1114(.a(G432), .O(gate155inter7));
  inv1  gate1115(.a(G525), .O(gate155inter8));
  nand2 gate1116(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1117(.a(s_81), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1118(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1119(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1120(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate547(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate548(.a(gate157inter0), .b(s_0), .O(gate157inter1));
  and2  gate549(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate550(.a(s_0), .O(gate157inter3));
  inv1  gate551(.a(s_1), .O(gate157inter4));
  nand2 gate552(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate553(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate554(.a(G438), .O(gate157inter7));
  inv1  gate555(.a(G528), .O(gate157inter8));
  nand2 gate556(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate557(.a(s_1), .b(gate157inter3), .O(gate157inter10));
  nor2  gate558(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate559(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate560(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate743(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate744(.a(gate168inter0), .b(s_28), .O(gate168inter1));
  and2  gate745(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate746(.a(s_28), .O(gate168inter3));
  inv1  gate747(.a(s_29), .O(gate168inter4));
  nand2 gate748(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate749(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate750(.a(G471), .O(gate168inter7));
  inv1  gate751(.a(G543), .O(gate168inter8));
  nand2 gate752(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate753(.a(s_29), .b(gate168inter3), .O(gate168inter10));
  nor2  gate754(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate755(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate756(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1079(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1080(.a(gate169inter0), .b(s_76), .O(gate169inter1));
  and2  gate1081(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1082(.a(s_76), .O(gate169inter3));
  inv1  gate1083(.a(s_77), .O(gate169inter4));
  nand2 gate1084(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1085(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1086(.a(G474), .O(gate169inter7));
  inv1  gate1087(.a(G546), .O(gate169inter8));
  nand2 gate1088(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1089(.a(s_77), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1090(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1091(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1092(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1177(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1178(.a(gate171inter0), .b(s_90), .O(gate171inter1));
  and2  gate1179(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1180(.a(s_90), .O(gate171inter3));
  inv1  gate1181(.a(s_91), .O(gate171inter4));
  nand2 gate1182(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1183(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1184(.a(G480), .O(gate171inter7));
  inv1  gate1185(.a(G549), .O(gate171inter8));
  nand2 gate1186(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1187(.a(s_91), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1188(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1189(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1190(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1667(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1668(.a(gate172inter0), .b(s_160), .O(gate172inter1));
  and2  gate1669(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1670(.a(s_160), .O(gate172inter3));
  inv1  gate1671(.a(s_161), .O(gate172inter4));
  nand2 gate1672(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1673(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1674(.a(G483), .O(gate172inter7));
  inv1  gate1675(.a(G549), .O(gate172inter8));
  nand2 gate1676(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1677(.a(s_161), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1678(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1679(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1680(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1527(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1528(.a(gate177inter0), .b(s_140), .O(gate177inter1));
  and2  gate1529(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1530(.a(s_140), .O(gate177inter3));
  inv1  gate1531(.a(s_141), .O(gate177inter4));
  nand2 gate1532(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1533(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1534(.a(G498), .O(gate177inter7));
  inv1  gate1535(.a(G558), .O(gate177inter8));
  nand2 gate1536(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1537(.a(s_141), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1538(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1539(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1540(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate715(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate716(.a(gate184inter0), .b(s_24), .O(gate184inter1));
  and2  gate717(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate718(.a(s_24), .O(gate184inter3));
  inv1  gate719(.a(s_25), .O(gate184inter4));
  nand2 gate720(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate721(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate722(.a(G519), .O(gate184inter7));
  inv1  gate723(.a(G567), .O(gate184inter8));
  nand2 gate724(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate725(.a(s_25), .b(gate184inter3), .O(gate184inter10));
  nor2  gate726(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate727(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate728(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1037(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1038(.a(gate185inter0), .b(s_70), .O(gate185inter1));
  and2  gate1039(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1040(.a(s_70), .O(gate185inter3));
  inv1  gate1041(.a(s_71), .O(gate185inter4));
  nand2 gate1042(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1043(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1044(.a(G570), .O(gate185inter7));
  inv1  gate1045(.a(G571), .O(gate185inter8));
  nand2 gate1046(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1047(.a(s_71), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1048(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1049(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1050(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1597(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1598(.a(gate189inter0), .b(s_150), .O(gate189inter1));
  and2  gate1599(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1600(.a(s_150), .O(gate189inter3));
  inv1  gate1601(.a(s_151), .O(gate189inter4));
  nand2 gate1602(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1603(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1604(.a(G578), .O(gate189inter7));
  inv1  gate1605(.a(G579), .O(gate189inter8));
  nand2 gate1606(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1607(.a(s_151), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1608(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1609(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1610(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1163(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1164(.a(gate193inter0), .b(s_88), .O(gate193inter1));
  and2  gate1165(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1166(.a(s_88), .O(gate193inter3));
  inv1  gate1167(.a(s_89), .O(gate193inter4));
  nand2 gate1168(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1169(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1170(.a(G586), .O(gate193inter7));
  inv1  gate1171(.a(G587), .O(gate193inter8));
  nand2 gate1172(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1173(.a(s_89), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1174(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1175(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1176(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1541(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1542(.a(gate194inter0), .b(s_142), .O(gate194inter1));
  and2  gate1543(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1544(.a(s_142), .O(gate194inter3));
  inv1  gate1545(.a(s_143), .O(gate194inter4));
  nand2 gate1546(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1547(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1548(.a(G588), .O(gate194inter7));
  inv1  gate1549(.a(G589), .O(gate194inter8));
  nand2 gate1550(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1551(.a(s_143), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1552(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1553(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1554(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1345(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1346(.a(gate196inter0), .b(s_114), .O(gate196inter1));
  and2  gate1347(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1348(.a(s_114), .O(gate196inter3));
  inv1  gate1349(.a(s_115), .O(gate196inter4));
  nand2 gate1350(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1351(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1352(.a(G592), .O(gate196inter7));
  inv1  gate1353(.a(G593), .O(gate196inter8));
  nand2 gate1354(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1355(.a(s_115), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1356(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1357(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1358(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate729(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate730(.a(gate197inter0), .b(s_26), .O(gate197inter1));
  and2  gate731(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate732(.a(s_26), .O(gate197inter3));
  inv1  gate733(.a(s_27), .O(gate197inter4));
  nand2 gate734(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate735(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate736(.a(G594), .O(gate197inter7));
  inv1  gate737(.a(G595), .O(gate197inter8));
  nand2 gate738(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate739(.a(s_27), .b(gate197inter3), .O(gate197inter10));
  nor2  gate740(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate741(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate742(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate687(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate688(.a(gate198inter0), .b(s_20), .O(gate198inter1));
  and2  gate689(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate690(.a(s_20), .O(gate198inter3));
  inv1  gate691(.a(s_21), .O(gate198inter4));
  nand2 gate692(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate693(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate694(.a(G596), .O(gate198inter7));
  inv1  gate695(.a(G597), .O(gate198inter8));
  nand2 gate696(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate697(.a(s_21), .b(gate198inter3), .O(gate198inter10));
  nor2  gate698(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate699(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate700(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1149(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1150(.a(gate201inter0), .b(s_86), .O(gate201inter1));
  and2  gate1151(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1152(.a(s_86), .O(gate201inter3));
  inv1  gate1153(.a(s_87), .O(gate201inter4));
  nand2 gate1154(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1155(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1156(.a(G602), .O(gate201inter7));
  inv1  gate1157(.a(G607), .O(gate201inter8));
  nand2 gate1158(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1159(.a(s_87), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1160(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1161(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1162(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1121(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1122(.a(gate202inter0), .b(s_82), .O(gate202inter1));
  and2  gate1123(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1124(.a(s_82), .O(gate202inter3));
  inv1  gate1125(.a(s_83), .O(gate202inter4));
  nand2 gate1126(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1127(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1128(.a(G612), .O(gate202inter7));
  inv1  gate1129(.a(G617), .O(gate202inter8));
  nand2 gate1130(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1131(.a(s_83), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1132(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1133(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1134(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1289(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1290(.a(gate210inter0), .b(s_106), .O(gate210inter1));
  and2  gate1291(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1292(.a(s_106), .O(gate210inter3));
  inv1  gate1293(.a(s_107), .O(gate210inter4));
  nand2 gate1294(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1295(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1296(.a(G607), .O(gate210inter7));
  inv1  gate1297(.a(G666), .O(gate210inter8));
  nand2 gate1298(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1299(.a(s_107), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1300(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1301(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1302(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate589(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate590(.a(gate212inter0), .b(s_6), .O(gate212inter1));
  and2  gate591(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate592(.a(s_6), .O(gate212inter3));
  inv1  gate593(.a(s_7), .O(gate212inter4));
  nand2 gate594(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate595(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate596(.a(G617), .O(gate212inter7));
  inv1  gate597(.a(G669), .O(gate212inter8));
  nand2 gate598(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate599(.a(s_7), .b(gate212inter3), .O(gate212inter10));
  nor2  gate600(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate601(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate602(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate659(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate660(.a(gate213inter0), .b(s_16), .O(gate213inter1));
  and2  gate661(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate662(.a(s_16), .O(gate213inter3));
  inv1  gate663(.a(s_17), .O(gate213inter4));
  nand2 gate664(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate665(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate666(.a(G602), .O(gate213inter7));
  inv1  gate667(.a(G672), .O(gate213inter8));
  nand2 gate668(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate669(.a(s_17), .b(gate213inter3), .O(gate213inter10));
  nor2  gate670(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate671(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate672(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate561(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate562(.a(gate223inter0), .b(s_2), .O(gate223inter1));
  and2  gate563(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate564(.a(s_2), .O(gate223inter3));
  inv1  gate565(.a(s_3), .O(gate223inter4));
  nand2 gate566(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate567(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate568(.a(G627), .O(gate223inter7));
  inv1  gate569(.a(G687), .O(gate223inter8));
  nand2 gate570(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate571(.a(s_3), .b(gate223inter3), .O(gate223inter10));
  nor2  gate572(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate573(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate574(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1555(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1556(.a(gate230inter0), .b(s_144), .O(gate230inter1));
  and2  gate1557(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1558(.a(s_144), .O(gate230inter3));
  inv1  gate1559(.a(s_145), .O(gate230inter4));
  nand2 gate1560(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1561(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1562(.a(G700), .O(gate230inter7));
  inv1  gate1563(.a(G701), .O(gate230inter8));
  nand2 gate1564(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1565(.a(s_145), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1566(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1567(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1568(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1331(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1332(.a(gate235inter0), .b(s_112), .O(gate235inter1));
  and2  gate1333(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1334(.a(s_112), .O(gate235inter3));
  inv1  gate1335(.a(s_113), .O(gate235inter4));
  nand2 gate1336(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1337(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1338(.a(G248), .O(gate235inter7));
  inv1  gate1339(.a(G724), .O(gate235inter8));
  nand2 gate1340(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1341(.a(s_113), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1342(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1343(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1344(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate869(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate870(.a(gate238inter0), .b(s_46), .O(gate238inter1));
  and2  gate871(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate872(.a(s_46), .O(gate238inter3));
  inv1  gate873(.a(s_47), .O(gate238inter4));
  nand2 gate874(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate875(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate876(.a(G257), .O(gate238inter7));
  inv1  gate877(.a(G709), .O(gate238inter8));
  nand2 gate878(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate879(.a(s_47), .b(gate238inter3), .O(gate238inter10));
  nor2  gate880(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate881(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate882(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1275(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1276(.a(gate240inter0), .b(s_104), .O(gate240inter1));
  and2  gate1277(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1278(.a(s_104), .O(gate240inter3));
  inv1  gate1279(.a(s_105), .O(gate240inter4));
  nand2 gate1280(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1281(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1282(.a(G263), .O(gate240inter7));
  inv1  gate1283(.a(G715), .O(gate240inter8));
  nand2 gate1284(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1285(.a(s_105), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1286(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1287(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1288(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate925(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate926(.a(gate244inter0), .b(s_54), .O(gate244inter1));
  and2  gate927(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate928(.a(s_54), .O(gate244inter3));
  inv1  gate929(.a(s_55), .O(gate244inter4));
  nand2 gate930(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate931(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate932(.a(G721), .O(gate244inter7));
  inv1  gate933(.a(G733), .O(gate244inter8));
  nand2 gate934(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate935(.a(s_55), .b(gate244inter3), .O(gate244inter10));
  nor2  gate936(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate937(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate938(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate1219(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1220(.a(gate245inter0), .b(s_96), .O(gate245inter1));
  and2  gate1221(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1222(.a(s_96), .O(gate245inter3));
  inv1  gate1223(.a(s_97), .O(gate245inter4));
  nand2 gate1224(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1225(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1226(.a(G248), .O(gate245inter7));
  inv1  gate1227(.a(G736), .O(gate245inter8));
  nand2 gate1228(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1229(.a(s_97), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1230(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1231(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1232(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1443(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1444(.a(gate262inter0), .b(s_128), .O(gate262inter1));
  and2  gate1445(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1446(.a(s_128), .O(gate262inter3));
  inv1  gate1447(.a(s_129), .O(gate262inter4));
  nand2 gate1448(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1449(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1450(.a(G764), .O(gate262inter7));
  inv1  gate1451(.a(G765), .O(gate262inter8));
  nand2 gate1452(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1453(.a(s_129), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1454(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1455(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1456(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1415(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1416(.a(gate270inter0), .b(s_124), .O(gate270inter1));
  and2  gate1417(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1418(.a(s_124), .O(gate270inter3));
  inv1  gate1419(.a(s_125), .O(gate270inter4));
  nand2 gate1420(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1421(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1422(.a(G657), .O(gate270inter7));
  inv1  gate1423(.a(G785), .O(gate270inter8));
  nand2 gate1424(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1425(.a(s_125), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1426(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1427(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1428(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate771(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate772(.a(gate275inter0), .b(s_32), .O(gate275inter1));
  and2  gate773(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate774(.a(s_32), .O(gate275inter3));
  inv1  gate775(.a(s_33), .O(gate275inter4));
  nand2 gate776(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate777(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate778(.a(G645), .O(gate275inter7));
  inv1  gate779(.a(G797), .O(gate275inter8));
  nand2 gate780(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate781(.a(s_33), .b(gate275inter3), .O(gate275inter10));
  nor2  gate782(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate783(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate784(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate841(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate842(.a(gate277inter0), .b(s_42), .O(gate277inter1));
  and2  gate843(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate844(.a(s_42), .O(gate277inter3));
  inv1  gate845(.a(s_43), .O(gate277inter4));
  nand2 gate846(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate847(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate848(.a(G648), .O(gate277inter7));
  inv1  gate849(.a(G800), .O(gate277inter8));
  nand2 gate850(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate851(.a(s_43), .b(gate277inter3), .O(gate277inter10));
  nor2  gate852(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate853(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate854(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1653(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1654(.a(gate280inter0), .b(s_158), .O(gate280inter1));
  and2  gate1655(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1656(.a(s_158), .O(gate280inter3));
  inv1  gate1657(.a(s_159), .O(gate280inter4));
  nand2 gate1658(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1659(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1660(.a(G779), .O(gate280inter7));
  inv1  gate1661(.a(G803), .O(gate280inter8));
  nand2 gate1662(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1663(.a(s_159), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1664(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1665(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1666(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1009(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1010(.a(gate294inter0), .b(s_66), .O(gate294inter1));
  and2  gate1011(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1012(.a(s_66), .O(gate294inter3));
  inv1  gate1013(.a(s_67), .O(gate294inter4));
  nand2 gate1014(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1015(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1016(.a(G832), .O(gate294inter7));
  inv1  gate1017(.a(G833), .O(gate294inter8));
  nand2 gate1018(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1019(.a(s_67), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1020(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1021(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1022(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1317(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1318(.a(gate295inter0), .b(s_110), .O(gate295inter1));
  and2  gate1319(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1320(.a(s_110), .O(gate295inter3));
  inv1  gate1321(.a(s_111), .O(gate295inter4));
  nand2 gate1322(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1323(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1324(.a(G830), .O(gate295inter7));
  inv1  gate1325(.a(G831), .O(gate295inter8));
  nand2 gate1326(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1327(.a(s_111), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1328(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1329(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1330(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1639(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1640(.a(gate296inter0), .b(s_156), .O(gate296inter1));
  and2  gate1641(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1642(.a(s_156), .O(gate296inter3));
  inv1  gate1643(.a(s_157), .O(gate296inter4));
  nand2 gate1644(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1645(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1646(.a(G826), .O(gate296inter7));
  inv1  gate1647(.a(G827), .O(gate296inter8));
  nand2 gate1648(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1649(.a(s_157), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1650(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1651(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1652(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1429(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1430(.a(gate388inter0), .b(s_126), .O(gate388inter1));
  and2  gate1431(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1432(.a(s_126), .O(gate388inter3));
  inv1  gate1433(.a(s_127), .O(gate388inter4));
  nand2 gate1434(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1435(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1436(.a(G2), .O(gate388inter7));
  inv1  gate1437(.a(G1039), .O(gate388inter8));
  nand2 gate1438(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1439(.a(s_127), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1440(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1441(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1442(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate701(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate702(.a(gate393inter0), .b(s_22), .O(gate393inter1));
  and2  gate703(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate704(.a(s_22), .O(gate393inter3));
  inv1  gate705(.a(s_23), .O(gate393inter4));
  nand2 gate706(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate707(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate708(.a(G7), .O(gate393inter7));
  inv1  gate709(.a(G1054), .O(gate393inter8));
  nand2 gate710(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate711(.a(s_23), .b(gate393inter3), .O(gate393inter10));
  nor2  gate712(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate713(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate714(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate1373(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1374(.a(gate394inter0), .b(s_118), .O(gate394inter1));
  and2  gate1375(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1376(.a(s_118), .O(gate394inter3));
  inv1  gate1377(.a(s_119), .O(gate394inter4));
  nand2 gate1378(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1379(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1380(.a(G8), .O(gate394inter7));
  inv1  gate1381(.a(G1057), .O(gate394inter8));
  nand2 gate1382(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1383(.a(s_119), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1384(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1385(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1386(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate603(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate604(.a(gate396inter0), .b(s_8), .O(gate396inter1));
  and2  gate605(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate606(.a(s_8), .O(gate396inter3));
  inv1  gate607(.a(s_9), .O(gate396inter4));
  nand2 gate608(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate609(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate610(.a(G10), .O(gate396inter7));
  inv1  gate611(.a(G1063), .O(gate396inter8));
  nand2 gate612(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate613(.a(s_9), .b(gate396inter3), .O(gate396inter10));
  nor2  gate614(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate615(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate616(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1625(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1626(.a(gate398inter0), .b(s_154), .O(gate398inter1));
  and2  gate1627(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1628(.a(s_154), .O(gate398inter3));
  inv1  gate1629(.a(s_155), .O(gate398inter4));
  nand2 gate1630(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1631(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1632(.a(G12), .O(gate398inter7));
  inv1  gate1633(.a(G1069), .O(gate398inter8));
  nand2 gate1634(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1635(.a(s_155), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1636(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1637(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1638(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1261(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1262(.a(gate402inter0), .b(s_102), .O(gate402inter1));
  and2  gate1263(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1264(.a(s_102), .O(gate402inter3));
  inv1  gate1265(.a(s_103), .O(gate402inter4));
  nand2 gate1266(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1267(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1268(.a(G16), .O(gate402inter7));
  inv1  gate1269(.a(G1081), .O(gate402inter8));
  nand2 gate1270(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1271(.a(s_103), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1272(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1273(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1274(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate981(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate982(.a(gate403inter0), .b(s_62), .O(gate403inter1));
  and2  gate983(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate984(.a(s_62), .O(gate403inter3));
  inv1  gate985(.a(s_63), .O(gate403inter4));
  nand2 gate986(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate987(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate988(.a(G17), .O(gate403inter7));
  inv1  gate989(.a(G1084), .O(gate403inter8));
  nand2 gate990(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate991(.a(s_63), .b(gate403inter3), .O(gate403inter10));
  nor2  gate992(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate993(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate994(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate967(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate968(.a(gate410inter0), .b(s_60), .O(gate410inter1));
  and2  gate969(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate970(.a(s_60), .O(gate410inter3));
  inv1  gate971(.a(s_61), .O(gate410inter4));
  nand2 gate972(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate973(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate974(.a(G24), .O(gate410inter7));
  inv1  gate975(.a(G1105), .O(gate410inter8));
  nand2 gate976(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate977(.a(s_61), .b(gate410inter3), .O(gate410inter10));
  nor2  gate978(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate979(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate980(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1569(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1570(.a(gate412inter0), .b(s_146), .O(gate412inter1));
  and2  gate1571(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1572(.a(s_146), .O(gate412inter3));
  inv1  gate1573(.a(s_147), .O(gate412inter4));
  nand2 gate1574(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1575(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1576(.a(G26), .O(gate412inter7));
  inv1  gate1577(.a(G1111), .O(gate412inter8));
  nand2 gate1578(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1579(.a(s_147), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1580(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1581(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1582(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate953(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate954(.a(gate414inter0), .b(s_58), .O(gate414inter1));
  and2  gate955(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate956(.a(s_58), .O(gate414inter3));
  inv1  gate957(.a(s_59), .O(gate414inter4));
  nand2 gate958(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate959(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate960(.a(G28), .O(gate414inter7));
  inv1  gate961(.a(G1117), .O(gate414inter8));
  nand2 gate962(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate963(.a(s_59), .b(gate414inter3), .O(gate414inter10));
  nor2  gate964(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate965(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate966(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1023(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1024(.a(gate418inter0), .b(s_68), .O(gate418inter1));
  and2  gate1025(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1026(.a(s_68), .O(gate418inter3));
  inv1  gate1027(.a(s_69), .O(gate418inter4));
  nand2 gate1028(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1029(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1030(.a(G32), .O(gate418inter7));
  inv1  gate1031(.a(G1129), .O(gate418inter8));
  nand2 gate1032(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1033(.a(s_69), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1034(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1035(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1036(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1387(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1388(.a(gate427inter0), .b(s_120), .O(gate427inter1));
  and2  gate1389(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1390(.a(s_120), .O(gate427inter3));
  inv1  gate1391(.a(s_121), .O(gate427inter4));
  nand2 gate1392(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1393(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1394(.a(G5), .O(gate427inter7));
  inv1  gate1395(.a(G1144), .O(gate427inter8));
  nand2 gate1396(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1397(.a(s_121), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1398(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1399(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1400(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1513(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1514(.a(gate435inter0), .b(s_138), .O(gate435inter1));
  and2  gate1515(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1516(.a(s_138), .O(gate435inter3));
  inv1  gate1517(.a(s_139), .O(gate435inter4));
  nand2 gate1518(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1519(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1520(.a(G9), .O(gate435inter7));
  inv1  gate1521(.a(G1156), .O(gate435inter8));
  nand2 gate1522(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1523(.a(s_139), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1524(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1525(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1526(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1247(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1248(.a(gate446inter0), .b(s_100), .O(gate446inter1));
  and2  gate1249(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1250(.a(s_100), .O(gate446inter3));
  inv1  gate1251(.a(s_101), .O(gate446inter4));
  nand2 gate1252(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1253(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1254(.a(G1075), .O(gate446inter7));
  inv1  gate1255(.a(G1171), .O(gate446inter8));
  nand2 gate1256(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1257(.a(s_101), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1258(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1259(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1260(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1471(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1472(.a(gate448inter0), .b(s_132), .O(gate448inter1));
  and2  gate1473(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1474(.a(s_132), .O(gate448inter3));
  inv1  gate1475(.a(s_133), .O(gate448inter4));
  nand2 gate1476(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1477(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1478(.a(G1078), .O(gate448inter7));
  inv1  gate1479(.a(G1174), .O(gate448inter8));
  nand2 gate1480(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1481(.a(s_133), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1482(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1483(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1484(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate645(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate646(.a(gate449inter0), .b(s_14), .O(gate449inter1));
  and2  gate647(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate648(.a(s_14), .O(gate449inter3));
  inv1  gate649(.a(s_15), .O(gate449inter4));
  nand2 gate650(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate651(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate652(.a(G16), .O(gate449inter7));
  inv1  gate653(.a(G1177), .O(gate449inter8));
  nand2 gate654(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate655(.a(s_15), .b(gate449inter3), .O(gate449inter10));
  nor2  gate656(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate657(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate658(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1485(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1486(.a(gate451inter0), .b(s_134), .O(gate451inter1));
  and2  gate1487(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1488(.a(s_134), .O(gate451inter3));
  inv1  gate1489(.a(s_135), .O(gate451inter4));
  nand2 gate1490(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1491(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1492(.a(G17), .O(gate451inter7));
  inv1  gate1493(.a(G1180), .O(gate451inter8));
  nand2 gate1494(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1495(.a(s_135), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1496(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1497(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1498(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate799(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate800(.a(gate477inter0), .b(s_36), .O(gate477inter1));
  and2  gate801(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate802(.a(s_36), .O(gate477inter3));
  inv1  gate803(.a(s_37), .O(gate477inter4));
  nand2 gate804(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate805(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate806(.a(G30), .O(gate477inter7));
  inv1  gate807(.a(G1219), .O(gate477inter8));
  nand2 gate808(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate809(.a(s_37), .b(gate477inter3), .O(gate477inter10));
  nor2  gate810(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate811(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate812(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1499(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1500(.a(gate481inter0), .b(s_136), .O(gate481inter1));
  and2  gate1501(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1502(.a(s_136), .O(gate481inter3));
  inv1  gate1503(.a(s_137), .O(gate481inter4));
  nand2 gate1504(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1505(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1506(.a(G32), .O(gate481inter7));
  inv1  gate1507(.a(G1225), .O(gate481inter8));
  nand2 gate1508(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1509(.a(s_137), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1510(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1511(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1512(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1205(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1206(.a(gate487inter0), .b(s_94), .O(gate487inter1));
  and2  gate1207(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1208(.a(s_94), .O(gate487inter3));
  inv1  gate1209(.a(s_95), .O(gate487inter4));
  nand2 gate1210(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1211(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1212(.a(G1236), .O(gate487inter7));
  inv1  gate1213(.a(G1237), .O(gate487inter8));
  nand2 gate1214(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1215(.a(s_95), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1216(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1217(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1218(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate939(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate940(.a(gate490inter0), .b(s_56), .O(gate490inter1));
  and2  gate941(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate942(.a(s_56), .O(gate490inter3));
  inv1  gate943(.a(s_57), .O(gate490inter4));
  nand2 gate944(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate945(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate946(.a(G1242), .O(gate490inter7));
  inv1  gate947(.a(G1243), .O(gate490inter8));
  nand2 gate948(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate949(.a(s_57), .b(gate490inter3), .O(gate490inter10));
  nor2  gate950(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate951(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate952(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate757(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate758(.a(gate496inter0), .b(s_30), .O(gate496inter1));
  and2  gate759(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate760(.a(s_30), .O(gate496inter3));
  inv1  gate761(.a(s_31), .O(gate496inter4));
  nand2 gate762(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate763(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate764(.a(G1254), .O(gate496inter7));
  inv1  gate765(.a(G1255), .O(gate496inter8));
  nand2 gate766(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate767(.a(s_31), .b(gate496inter3), .O(gate496inter10));
  nor2  gate768(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate769(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate770(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1135(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1136(.a(gate499inter0), .b(s_84), .O(gate499inter1));
  and2  gate1137(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1138(.a(s_84), .O(gate499inter3));
  inv1  gate1139(.a(s_85), .O(gate499inter4));
  nand2 gate1140(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1141(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1142(.a(G1260), .O(gate499inter7));
  inv1  gate1143(.a(G1261), .O(gate499inter8));
  nand2 gate1144(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1145(.a(s_85), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1146(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1147(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1148(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate897(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate898(.a(gate504inter0), .b(s_50), .O(gate504inter1));
  and2  gate899(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate900(.a(s_50), .O(gate504inter3));
  inv1  gate901(.a(s_51), .O(gate504inter4));
  nand2 gate902(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate903(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate904(.a(G1270), .O(gate504inter7));
  inv1  gate905(.a(G1271), .O(gate504inter8));
  nand2 gate906(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate907(.a(s_51), .b(gate504inter3), .O(gate504inter10));
  nor2  gate908(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate909(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate910(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1191(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1192(.a(gate509inter0), .b(s_92), .O(gate509inter1));
  and2  gate1193(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1194(.a(s_92), .O(gate509inter3));
  inv1  gate1195(.a(s_93), .O(gate509inter4));
  nand2 gate1196(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1197(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1198(.a(G1280), .O(gate509inter7));
  inv1  gate1199(.a(G1281), .O(gate509inter8));
  nand2 gate1200(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1201(.a(s_93), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1202(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1203(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1204(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1709(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1710(.a(gate511inter0), .b(s_166), .O(gate511inter1));
  and2  gate1711(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1712(.a(s_166), .O(gate511inter3));
  inv1  gate1713(.a(s_167), .O(gate511inter4));
  nand2 gate1714(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1715(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1716(.a(G1284), .O(gate511inter7));
  inv1  gate1717(.a(G1285), .O(gate511inter8));
  nand2 gate1718(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1719(.a(s_167), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1720(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1721(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1722(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule