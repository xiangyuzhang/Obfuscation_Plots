module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate7inter0, gate7inter1, gate7inter2, gate7inter3, gate7inter4, gate7inter5, gate7inter6, gate7inter7, gate7inter8, gate7inter9, gate7inter10, gate7inter11, gate7inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );

  xor2  gate301(.a(N53), .b(N49), .O(gate7inter0));
  nand2 gate302(.a(gate7inter0), .b(s_14), .O(gate7inter1));
  and2  gate303(.a(N53), .b(N49), .O(gate7inter2));
  inv1  gate304(.a(s_14), .O(gate7inter3));
  inv1  gate305(.a(s_15), .O(gate7inter4));
  nand2 gate306(.a(gate7inter4), .b(gate7inter3), .O(gate7inter5));
  nor2  gate307(.a(gate7inter5), .b(gate7inter2), .O(gate7inter6));
  inv1  gate308(.a(N49), .O(gate7inter7));
  inv1  gate309(.a(N53), .O(gate7inter8));
  nand2 gate310(.a(gate7inter8), .b(gate7inter7), .O(gate7inter9));
  nand2 gate311(.a(s_15), .b(gate7inter3), .O(gate7inter10));
  nor2  gate312(.a(gate7inter10), .b(gate7inter9), .O(gate7inter11));
  nor2  gate313(.a(gate7inter11), .b(gate7inter6), .O(gate7inter12));
  nand2 gate314(.a(gate7inter12), .b(gate7inter1), .O(N256));
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );

  xor2  gate371(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate372(.a(gate13inter0), .b(s_24), .O(gate13inter1));
  and2  gate373(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate374(.a(s_24), .O(gate13inter3));
  inv1  gate375(.a(s_25), .O(gate13inter4));
  nand2 gate376(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate377(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate378(.a(N97), .O(gate13inter7));
  inv1  gate379(.a(N101), .O(gate13inter8));
  nand2 gate380(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate381(.a(s_25), .b(gate13inter3), .O(gate13inter10));
  nor2  gate382(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate383(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate384(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate343(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate344(.a(gate42inter0), .b(s_20), .O(gate42inter1));
  and2  gate345(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate346(.a(s_20), .O(gate42inter3));
  inv1  gate347(.a(s_21), .O(gate42inter4));
  nand2 gate348(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate349(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate350(.a(N252), .O(gate42inter7));
  inv1  gate351(.a(N253), .O(gate42inter8));
  nand2 gate352(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate353(.a(s_21), .b(gate42inter3), .O(gate42inter10));
  nor2  gate354(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate355(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate356(.a(gate42inter12), .b(gate42inter1), .O(N293));

  xor2  gate329(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate330(.a(gate43inter0), .b(s_18), .O(gate43inter1));
  and2  gate331(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate332(.a(s_18), .O(gate43inter3));
  inv1  gate333(.a(s_19), .O(gate43inter4));
  nand2 gate334(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate335(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate336(.a(N254), .O(gate43inter7));
  inv1  gate337(.a(N255), .O(gate43inter8));
  nand2 gate338(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate339(.a(s_19), .b(gate43inter3), .O(gate43inter10));
  nor2  gate340(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate341(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate342(.a(gate43inter12), .b(gate43inter1), .O(N296));
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );

  xor2  gate399(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate400(.a(gate51inter0), .b(s_28), .O(gate51inter1));
  and2  gate401(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate402(.a(s_28), .O(gate51inter3));
  inv1  gate403(.a(s_29), .O(gate51inter4));
  nand2 gate404(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate405(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate406(.a(N278), .O(gate51inter7));
  inv1  gate407(.a(N279), .O(gate51inter8));
  nand2 gate408(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate409(.a(s_29), .b(gate51inter3), .O(gate51inter10));
  nor2  gate410(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate411(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate412(.a(gate51inter12), .b(gate51inter1), .O(N316));
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );

  xor2  gate413(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate414(.a(gate57inter0), .b(s_30), .O(gate57inter1));
  and2  gate415(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate416(.a(s_30), .O(gate57inter3));
  inv1  gate417(.a(s_31), .O(gate57inter4));
  nand2 gate418(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate419(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate420(.a(N290), .O(gate57inter7));
  inv1  gate421(.a(N293), .O(gate57inter8));
  nand2 gate422(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate423(.a(s_31), .b(gate57inter3), .O(gate57inter10));
  nor2  gate424(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate425(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate426(.a(gate57inter12), .b(gate57inter1), .O(N338));
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );

  xor2  gate385(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate386(.a(gate60inter0), .b(s_26), .O(gate60inter1));
  and2  gate387(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate388(.a(s_26), .O(gate60inter3));
  inv1  gate389(.a(s_27), .O(gate60inter4));
  nand2 gate390(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate391(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate392(.a(N293), .O(gate60inter7));
  inv1  gate393(.a(N299), .O(gate60inter8));
  nand2 gate394(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate395(.a(s_27), .b(gate60inter3), .O(gate60inter10));
  nor2  gate396(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate397(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate398(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate259(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate260(.a(gate62inter0), .b(s_8), .O(gate62inter1));
  and2  gate261(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate262(.a(s_8), .O(gate62inter3));
  inv1  gate263(.a(s_9), .O(gate62inter4));
  nand2 gate264(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate265(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate266(.a(N308), .O(gate62inter7));
  inv1  gate267(.a(N311), .O(gate62inter8));
  nand2 gate268(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate269(.a(s_9), .b(gate62inter3), .O(gate62inter10));
  nor2  gate270(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate271(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate272(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );

  xor2  gate231(.a(N695), .b(N13), .O(gate174inter0));
  nand2 gate232(.a(gate174inter0), .b(s_4), .O(gate174inter1));
  and2  gate233(.a(N695), .b(N13), .O(gate174inter2));
  inv1  gate234(.a(s_4), .O(gate174inter3));
  inv1  gate235(.a(s_5), .O(gate174inter4));
  nand2 gate236(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate237(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate238(.a(N13), .O(gate174inter7));
  inv1  gate239(.a(N695), .O(gate174inter8));
  nand2 gate240(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate241(.a(s_5), .b(gate174inter3), .O(gate174inter10));
  nor2  gate242(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate243(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate244(.a(gate174inter12), .b(gate174inter1), .O(N727));
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );

  xor2  gate315(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate316(.a(gate178inter0), .b(s_16), .O(gate178inter1));
  and2  gate317(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate318(.a(s_16), .O(gate178inter3));
  inv1  gate319(.a(s_17), .O(gate178inter4));
  nand2 gate320(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate321(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate322(.a(N29), .O(gate178inter7));
  inv1  gate323(.a(N699), .O(gate178inter8));
  nand2 gate324(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate325(.a(s_17), .b(gate178inter3), .O(gate178inter10));
  nor2  gate326(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate327(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate328(.a(gate178inter12), .b(gate178inter1), .O(N731));

  xor2  gate287(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate288(.a(gate179inter0), .b(s_12), .O(gate179inter1));
  and2  gate289(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate290(.a(s_12), .O(gate179inter3));
  inv1  gate291(.a(s_13), .O(gate179inter4));
  nand2 gate292(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate293(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate294(.a(N33), .O(gate179inter7));
  inv1  gate295(.a(N700), .O(gate179inter8));
  nand2 gate296(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate297(.a(s_13), .b(gate179inter3), .O(gate179inter10));
  nor2  gate298(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate299(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate300(.a(gate179inter12), .b(gate179inter1), .O(N732));

  xor2  gate217(.a(N701), .b(N37), .O(gate180inter0));
  nand2 gate218(.a(gate180inter0), .b(s_2), .O(gate180inter1));
  and2  gate219(.a(N701), .b(N37), .O(gate180inter2));
  inv1  gate220(.a(s_2), .O(gate180inter3));
  inv1  gate221(.a(s_3), .O(gate180inter4));
  nand2 gate222(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate223(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate224(.a(N37), .O(gate180inter7));
  inv1  gate225(.a(N701), .O(gate180inter8));
  nand2 gate226(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate227(.a(s_3), .b(gate180inter3), .O(gate180inter10));
  nor2  gate228(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate229(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate230(.a(gate180inter12), .b(gate180inter1), .O(N733));
xor2 gate181( .a(N41), .b(N702), .O(N734) );

  xor2  gate245(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate246(.a(gate182inter0), .b(s_6), .O(gate182inter1));
  and2  gate247(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate248(.a(s_6), .O(gate182inter3));
  inv1  gate249(.a(s_7), .O(gate182inter4));
  nand2 gate250(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate251(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate252(.a(N45), .O(gate182inter7));
  inv1  gate253(.a(N703), .O(gate182inter8));
  nand2 gate254(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate255(.a(s_7), .b(gate182inter3), .O(gate182inter10));
  nor2  gate256(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate257(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate258(.a(gate182inter12), .b(gate182inter1), .O(N735));
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );

  xor2  gate203(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate204(.a(gate194inter0), .b(s_0), .O(gate194inter1));
  and2  gate205(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate206(.a(s_0), .O(gate194inter3));
  inv1  gate207(.a(s_1), .O(gate194inter4));
  nand2 gate208(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate209(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate210(.a(N93), .O(gate194inter7));
  inv1  gate211(.a(N715), .O(gate194inter8));
  nand2 gate212(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate213(.a(s_1), .b(gate194inter3), .O(gate194inter10));
  nor2  gate214(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate215(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate216(.a(gate194inter12), .b(gate194inter1), .O(N747));
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );

  xor2  gate273(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate274(.a(gate198inter0), .b(s_10), .O(gate198inter1));
  and2  gate275(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate276(.a(s_10), .O(gate198inter3));
  inv1  gate277(.a(s_11), .O(gate198inter4));
  nand2 gate278(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate279(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate280(.a(N109), .O(gate198inter7));
  inv1  gate281(.a(N719), .O(gate198inter8));
  nand2 gate282(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate283(.a(s_11), .b(gate198inter3), .O(gate198inter10));
  nor2  gate284(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate285(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate286(.a(gate198inter12), .b(gate198inter1), .O(N751));

  xor2  gate357(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate358(.a(gate199inter0), .b(s_22), .O(gate199inter1));
  and2  gate359(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate360(.a(s_22), .O(gate199inter3));
  inv1  gate361(.a(s_23), .O(gate199inter4));
  nand2 gate362(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate363(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate364(.a(N113), .O(gate199inter7));
  inv1  gate365(.a(N720), .O(gate199inter8));
  nand2 gate366(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate367(.a(s_23), .b(gate199inter3), .O(gate199inter10));
  nor2  gate368(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate369(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate370(.a(gate199inter12), .b(gate199inter1), .O(N752));
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule