module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;
wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877, gate348inter0, gate348inter1, gate348inter2, gate348inter3, gate348inter4, gate348inter5, gate348inter6, gate348inter7, gate348inter8, gate348inter9, gate348inter10, gate348inter11, gate348inter12, gate344inter0, gate344inter1, gate344inter2, gate344inter3, gate344inter4, gate344inter5, gate344inter6, gate344inter7, gate344inter8, gate344inter9, gate344inter10, gate344inter11, gate344inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate311inter0, gate311inter1, gate311inter2, gate311inter3, gate311inter4, gate311inter5, gate311inter6, gate311inter7, gate311inter8, gate311inter9, gate311inter10, gate311inter11, gate311inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate315inter0, gate315inter1, gate315inter2, gate315inter3, gate315inter4, gate315inter5, gate315inter6, gate315inter7, gate315inter8, gate315inter9, gate315inter10, gate315inter11, gate315inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate327inter0, gate327inter1, gate327inter2, gate327inter3, gate327inter4, gate327inter5, gate327inter6, gate327inter7, gate327inter8, gate327inter9, gate327inter10, gate327inter11, gate327inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate307inter0, gate307inter1, gate307inter2, gate307inter3, gate307inter4, gate307inter5, gate307inter6, gate307inter7, gate307inter8, gate307inter9, gate307inter10, gate307inter11, gate307inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate302inter0, gate302inter1, gate302inter2, gate302inter3, gate302inter4, gate302inter5, gate302inter6, gate302inter7, gate302inter8, gate302inter9, gate302inter10, gate302inter11, gate302inter12, gate328inter0, gate328inter1, gate328inter2, gate328inter3, gate328inter4, gate328inter5, gate328inter6, gate328inter7, gate328inter8, gate328inter9, gate328inter10, gate328inter11, gate328inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate347inter0, gate347inter1, gate347inter2, gate347inter3, gate347inter4, gate347inter5, gate347inter6, gate347inter7, gate347inter8, gate347inter9, gate347inter10, gate347inter11, gate347inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12;


nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );
nand2 gate20( .a(N91), .b(N96), .O(N301) );
or2 gate21( .a(N91), .b(N96), .O(N302) );

  xor2  gate888(.a(N106), .b(N101), .O(gate22inter0));
  nand2 gate889(.a(gate22inter0), .b(s_72), .O(gate22inter1));
  and2  gate890(.a(N106), .b(N101), .O(gate22inter2));
  inv1  gate891(.a(s_72), .O(gate22inter3));
  inv1  gate892(.a(s_73), .O(gate22inter4));
  nand2 gate893(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate894(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate895(.a(N101), .O(gate22inter7));
  inv1  gate896(.a(N106), .O(gate22inter8));
  nand2 gate897(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate898(.a(s_73), .b(gate22inter3), .O(gate22inter10));
  nor2  gate899(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate900(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate901(.a(gate22inter12), .b(gate22inter1), .O(N303));
or2 gate23( .a(N101), .b(N106), .O(N304) );
nand2 gate24( .a(N111), .b(N116), .O(N305) );
or2 gate25( .a(N111), .b(N116), .O(N306) );
nand2 gate26( .a(N121), .b(N126), .O(N307) );
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );
nand2 gate33( .a(N59), .b(N156), .O(N319) );
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17), .b(N42), .O(N323) );

  xor2  gate426(.a(N165), .b(N159), .O(gate36inter0));
  nand2 gate427(.a(gate36inter0), .b(s_6), .O(gate36inter1));
  and2  gate428(.a(N165), .b(N159), .O(gate36inter2));
  inv1  gate429(.a(s_6), .O(gate36inter3));
  inv1  gate430(.a(s_7), .O(gate36inter4));
  nand2 gate431(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate432(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate433(.a(N159), .O(gate36inter7));
  inv1  gate434(.a(N165), .O(gate36inter8));
  nand2 gate435(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate436(.a(s_7), .b(gate36inter3), .O(gate36inter10));
  nor2  gate437(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate438(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate439(.a(gate36inter12), .b(gate36inter1), .O(N324));
or2 gate37( .a(N159), .b(N165), .O(N325) );
nand2 gate38( .a(N171), .b(N177), .O(N326) );
or2 gate39( .a(N171), .b(N177), .O(N327) );
nand2 gate40( .a(N183), .b(N189), .O(N328) );
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
and2 gate49( .a(N255), .b(N259), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );
nor2 gate60( .a(N280), .b(N284), .O(N348) );
or2 gate61( .a(N280), .b(N285), .O(N349) );
or2 gate62( .a(N280), .b(N286), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );
nand2 gate67( .a(N89), .b(N298), .O(N355) );
and2 gate68( .a(N90), .b(N298), .O(N356) );

  xor2  gate608(.a(N302), .b(N301), .O(gate69inter0));
  nand2 gate609(.a(gate69inter0), .b(s_32), .O(gate69inter1));
  and2  gate610(.a(N302), .b(N301), .O(gate69inter2));
  inv1  gate611(.a(s_32), .O(gate69inter3));
  inv1  gate612(.a(s_33), .O(gate69inter4));
  nand2 gate613(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate614(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate615(.a(N301), .O(gate69inter7));
  inv1  gate616(.a(N302), .O(gate69inter8));
  nand2 gate617(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate618(.a(s_33), .b(gate69inter3), .O(gate69inter10));
  nor2  gate619(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate620(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate621(.a(gate69inter12), .b(gate69inter1), .O(N357));
nand2 gate70( .a(N303), .b(N304), .O(N360) );

  xor2  gate412(.a(N306), .b(N305), .O(gate71inter0));
  nand2 gate413(.a(gate71inter0), .b(s_4), .O(gate71inter1));
  and2  gate414(.a(N306), .b(N305), .O(gate71inter2));
  inv1  gate415(.a(s_4), .O(gate71inter3));
  inv1  gate416(.a(s_5), .O(gate71inter4));
  nand2 gate417(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate418(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate419(.a(N305), .O(gate71inter7));
  inv1  gate420(.a(N306), .O(gate71inter8));
  nand2 gate421(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate422(.a(s_5), .b(gate71inter3), .O(gate71inter10));
  nor2  gate423(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate424(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate425(.a(gate71inter12), .b(gate71inter1), .O(N363));

  xor2  gate510(.a(N308), .b(N307), .O(gate72inter0));
  nand2 gate511(.a(gate72inter0), .b(s_18), .O(gate72inter1));
  and2  gate512(.a(N308), .b(N307), .O(gate72inter2));
  inv1  gate513(.a(s_18), .O(gate72inter3));
  inv1  gate514(.a(s_19), .O(gate72inter4));
  nand2 gate515(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate516(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate517(.a(N307), .O(gate72inter7));
  inv1  gate518(.a(N308), .O(gate72inter8));
  nand2 gate519(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate520(.a(s_19), .b(gate72inter3), .O(gate72inter10));
  nor2  gate521(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate522(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate523(.a(gate72inter12), .b(gate72inter1), .O(N366));
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );
nand2 gate76( .a(N326), .b(N327), .O(N379) );

  xor2  gate944(.a(N329), .b(N328), .O(gate77inter0));
  nand2 gate945(.a(gate77inter0), .b(s_80), .O(gate77inter1));
  and2  gate946(.a(N329), .b(N328), .O(gate77inter2));
  inv1  gate947(.a(s_80), .O(gate77inter3));
  inv1  gate948(.a(s_81), .O(gate77inter4));
  nand2 gate949(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate950(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate951(.a(N328), .O(gate77inter7));
  inv1  gate952(.a(N329), .O(gate77inter8));
  nand2 gate953(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate954(.a(s_81), .b(gate77inter3), .O(gate77inter10));
  nor2  gate955(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate956(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate957(.a(gate77inter12), .b(gate77inter1), .O(N382));
nand2 gate78( .a(N330), .b(N331), .O(N385) );
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );
nand2 gate96( .a(N347), .b(N352), .O(N410) );
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );
nor2 gate126( .a(N406), .b(N425), .O(N460) );

  xor2  gate818(.a(N426), .b(N409), .O(gate127inter0));
  nand2 gate819(.a(gate127inter0), .b(s_62), .O(gate127inter1));
  and2  gate820(.a(N426), .b(N409), .O(gate127inter2));
  inv1  gate821(.a(s_62), .O(gate127inter3));
  inv1  gate822(.a(s_63), .O(gate127inter4));
  nand2 gate823(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate824(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate825(.a(N409), .O(gate127inter7));
  inv1  gate826(.a(N426), .O(gate127inter8));
  nand2 gate827(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate828(.a(s_63), .b(gate127inter3), .O(gate127inter10));
  nor2  gate829(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate830(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate831(.a(gate127inter12), .b(gate127inter1), .O(N463));
nand2 gate128( .a(N442), .b(N410), .O(N466) );
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );
nand2 gate137( .a(N443), .b(N1), .O(N483) );
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );
nor2 gate142( .a(N413), .b(N444), .O(N492) );
nor2 gate143( .a(N416), .b(N445), .O(N495) );
nand2 gate144( .a(N130), .b(N460), .O(N498) );
or2 gate145( .a(N130), .b(N460), .O(N499) );
nand2 gate146( .a(N463), .b(N135), .O(N500) );
or2 gate147( .a(N463), .b(N135), .O(N501) );
and2 gate148( .a(N91), .b(N466), .O(N502) );

  xor2  gate524(.a(N476), .b(N475), .O(gate149inter0));
  nand2 gate525(.a(gate149inter0), .b(s_20), .O(gate149inter1));
  and2  gate526(.a(N476), .b(N475), .O(gate149inter2));
  inv1  gate527(.a(s_20), .O(gate149inter3));
  inv1  gate528(.a(s_21), .O(gate149inter4));
  nand2 gate529(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate530(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate531(.a(N475), .O(gate149inter7));
  inv1  gate532(.a(N476), .O(gate149inter8));
  nand2 gate533(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate534(.a(s_21), .b(gate149inter3), .O(gate149inter10));
  nor2  gate535(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate536(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate537(.a(gate149inter12), .b(gate149inter1), .O(N503));
and2 gate150( .a(N96), .b(N466), .O(N504) );
nor2 gate151( .a(N477), .b(N478), .O(N505) );
and2 gate152( .a(N101), .b(N466), .O(N506) );

  xor2  gate930(.a(N480), .b(N479), .O(gate153inter0));
  nand2 gate931(.a(gate153inter0), .b(s_78), .O(gate153inter1));
  and2  gate932(.a(N480), .b(N479), .O(gate153inter2));
  inv1  gate933(.a(s_78), .O(gate153inter3));
  inv1  gate934(.a(s_79), .O(gate153inter4));
  nand2 gate935(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate936(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate937(.a(N479), .O(gate153inter7));
  inv1  gate938(.a(N480), .O(gate153inter8));
  nand2 gate939(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate940(.a(s_79), .b(gate153inter3), .O(gate153inter10));
  nor2  gate941(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate942(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate943(.a(gate153inter12), .b(gate153inter1), .O(N507));
and2 gate154( .a(N106), .b(N466), .O(N508) );
nor2 gate155( .a(N481), .b(N482), .O(N509) );
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );

  xor2  gate496(.a(N492), .b(N130), .O(gate164inter0));
  nand2 gate497(.a(gate164inter0), .b(s_16), .O(gate164inter1));
  and2  gate498(.a(N492), .b(N130), .O(gate164inter2));
  inv1  gate499(.a(s_16), .O(gate164inter3));
  inv1  gate500(.a(s_17), .O(gate164inter4));
  nand2 gate501(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate502(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate503(.a(N130), .O(gate164inter7));
  inv1  gate504(.a(N492), .O(gate164inter8));
  nand2 gate505(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate506(.a(s_17), .b(gate164inter3), .O(gate164inter10));
  nor2  gate507(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate508(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate509(.a(gate164inter12), .b(gate164inter1), .O(N518));
or2 gate165( .a(N130), .b(N492), .O(N519) );
nand2 gate166( .a(N495), .b(N207), .O(N520) );
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
and2 gate170( .a(N451), .b(N171), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );

  xor2  gate706(.a(N189), .b(N451), .O(gate173inter0));
  nand2 gate707(.a(gate173inter0), .b(s_46), .O(gate173inter1));
  and2  gate708(.a(N189), .b(N451), .O(gate173inter2));
  inv1  gate709(.a(s_46), .O(gate173inter3));
  inv1  gate710(.a(s_47), .O(gate173inter4));
  nand2 gate711(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate712(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate713(.a(N451), .O(gate173inter7));
  inv1  gate714(.a(N189), .O(gate173inter8));
  nand2 gate715(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate716(.a(s_47), .b(gate173inter3), .O(gate173inter10));
  nor2  gate717(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate718(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate719(.a(gate173inter12), .b(gate173inter1), .O(N527));

  xor2  gate566(.a(N195), .b(N451), .O(gate174inter0));
  nand2 gate567(.a(gate174inter0), .b(s_26), .O(gate174inter1));
  and2  gate568(.a(N195), .b(N451), .O(gate174inter2));
  inv1  gate569(.a(s_26), .O(gate174inter3));
  inv1  gate570(.a(s_27), .O(gate174inter4));
  nand2 gate571(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate572(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate573(.a(N451), .O(gate174inter7));
  inv1  gate574(.a(N195), .O(gate174inter8));
  nand2 gate575(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate576(.a(s_27), .b(gate174inter3), .O(gate174inter10));
  nor2  gate577(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate578(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate579(.a(gate174inter12), .b(gate174inter1), .O(N528));
nand2 gate175( .a(N451), .b(N201), .O(N529) );
nand2 gate176( .a(N498), .b(N499), .O(N530) );
nand2 gate177( .a(N500), .b(N501), .O(N533) );
nor2 gate178( .a(N309), .b(N502), .O(N536) );
nor2 gate179( .a(N316), .b(N504), .O(N537) );

  xor2  gate580(.a(N506), .b(N317), .O(gate180inter0));
  nand2 gate581(.a(gate180inter0), .b(s_28), .O(gate180inter1));
  and2  gate582(.a(N506), .b(N317), .O(gate180inter2));
  inv1  gate583(.a(s_28), .O(gate180inter3));
  inv1  gate584(.a(s_29), .O(gate180inter4));
  nand2 gate585(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate586(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate587(.a(N317), .O(gate180inter7));
  inv1  gate588(.a(N506), .O(gate180inter8));
  nand2 gate589(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate590(.a(s_29), .b(gate180inter3), .O(gate180inter10));
  nor2  gate591(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate592(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate593(.a(gate180inter12), .b(gate180inter1), .O(N538));

  xor2  gate902(.a(N508), .b(N318), .O(gate181inter0));
  nand2 gate903(.a(gate181inter0), .b(s_74), .O(gate181inter1));
  and2  gate904(.a(N508), .b(N318), .O(gate181inter2));
  inv1  gate905(.a(s_74), .O(gate181inter3));
  inv1  gate906(.a(s_75), .O(gate181inter4));
  nand2 gate907(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate908(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate909(.a(N318), .O(gate181inter7));
  inv1  gate910(.a(N508), .O(gate181inter8));
  nand2 gate911(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate912(.a(s_75), .b(gate181inter3), .O(gate181inter10));
  nor2  gate913(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate914(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate915(.a(gate181inter12), .b(gate181inter1), .O(N539));
nor2 gate182( .a(N510), .b(N511), .O(N540) );
nor2 gate183( .a(N512), .b(N513), .O(N541) );

  xor2  gate440(.a(N515), .b(N514), .O(gate184inter0));
  nand2 gate441(.a(gate184inter0), .b(s_8), .O(gate184inter1));
  and2  gate442(.a(N515), .b(N514), .O(gate184inter2));
  inv1  gate443(.a(s_8), .O(gate184inter3));
  inv1  gate444(.a(s_9), .O(gate184inter4));
  nand2 gate445(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate446(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate447(.a(N514), .O(gate184inter7));
  inv1  gate448(.a(N515), .O(gate184inter8));
  nand2 gate449(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate450(.a(s_9), .b(gate184inter3), .O(gate184inter10));
  nor2  gate451(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate452(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate453(.a(gate184inter12), .b(gate184inter1), .O(N542));

  xor2  gate720(.a(N517), .b(N516), .O(gate185inter0));
  nand2 gate721(.a(gate185inter0), .b(s_48), .O(gate185inter1));
  and2  gate722(.a(N517), .b(N516), .O(gate185inter2));
  inv1  gate723(.a(s_48), .O(gate185inter3));
  inv1  gate724(.a(s_49), .O(gate185inter4));
  nand2 gate725(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate726(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate727(.a(N516), .O(gate185inter7));
  inv1  gate728(.a(N517), .O(gate185inter8));
  nand2 gate729(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate730(.a(s_49), .b(gate185inter3), .O(gate185inter10));
  nor2  gate731(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate732(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate733(.a(gate185inter12), .b(gate185inter1), .O(N543));

  xor2  gate622(.a(N519), .b(N518), .O(gate186inter0));
  nand2 gate623(.a(gate186inter0), .b(s_34), .O(gate186inter1));
  and2  gate624(.a(N519), .b(N518), .O(gate186inter2));
  inv1  gate625(.a(s_34), .O(gate186inter3));
  inv1  gate626(.a(s_35), .O(gate186inter4));
  nand2 gate627(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate628(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate629(.a(N518), .O(gate186inter7));
  inv1  gate630(.a(N519), .O(gate186inter8));
  nand2 gate631(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate632(.a(s_35), .b(gate186inter3), .O(gate186inter10));
  nor2  gate633(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate634(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate635(.a(gate186inter12), .b(gate186inter1), .O(N544));
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );
nand2 gate191( .a(N536), .b(N503), .O(N553) );

  xor2  gate552(.a(N505), .b(N537), .O(gate192inter0));
  nand2 gate553(.a(gate192inter0), .b(s_24), .O(gate192inter1));
  and2  gate554(.a(N505), .b(N537), .O(gate192inter2));
  inv1  gate555(.a(s_24), .O(gate192inter3));
  inv1  gate556(.a(s_25), .O(gate192inter4));
  nand2 gate557(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate558(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate559(.a(N537), .O(gate192inter7));
  inv1  gate560(.a(N505), .O(gate192inter8));
  nand2 gate561(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate562(.a(s_25), .b(gate192inter3), .O(gate192inter10));
  nor2  gate563(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate564(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate565(.a(gate192inter12), .b(gate192inter1), .O(N557));
nand2 gate193( .a(N538), .b(N507), .O(N561) );
nand2 gate194( .a(N539), .b(N509), .O(N565) );

  xor2  gate776(.a(N540), .b(N488), .O(gate195inter0));
  nand2 gate777(.a(gate195inter0), .b(s_56), .O(gate195inter1));
  and2  gate778(.a(N540), .b(N488), .O(gate195inter2));
  inv1  gate779(.a(s_56), .O(gate195inter3));
  inv1  gate780(.a(s_57), .O(gate195inter4));
  nand2 gate781(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate782(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate783(.a(N488), .O(gate195inter7));
  inv1  gate784(.a(N540), .O(gate195inter8));
  nand2 gate785(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate786(.a(s_57), .b(gate195inter3), .O(gate195inter10));
  nor2  gate787(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate788(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate789(.a(gate195inter12), .b(gate195inter1), .O(N569));
nand2 gate196( .a(N489), .b(N541), .O(N573) );
nand2 gate197( .a(N490), .b(N542), .O(N577) );

  xor2  gate650(.a(N543), .b(N491), .O(gate198inter0));
  nand2 gate651(.a(gate198inter0), .b(s_38), .O(gate198inter1));
  and2  gate652(.a(N543), .b(N491), .O(gate198inter2));
  inv1  gate653(.a(s_38), .O(gate198inter3));
  inv1  gate654(.a(s_39), .O(gate198inter4));
  nand2 gate655(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate656(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate657(.a(N491), .O(gate198inter7));
  inv1  gate658(.a(N543), .O(gate198inter8));
  nand2 gate659(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate660(.a(s_39), .b(gate198inter3), .O(gate198inter10));
  nor2  gate661(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate662(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate663(.a(gate198inter12), .b(gate198inter1), .O(N581));
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );
nand2 gate204( .a(N553), .b(N159), .O(N590) );
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );

  xor2  gate804(.a(N165), .b(N557), .O(gate207inter0));
  nand2 gate805(.a(gate207inter0), .b(s_60), .O(gate207inter1));
  and2  gate806(.a(N165), .b(N557), .O(gate207inter2));
  inv1  gate807(.a(s_60), .O(gate207inter3));
  inv1  gate808(.a(s_61), .O(gate207inter4));
  nand2 gate809(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate810(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate811(.a(N557), .O(gate207inter7));
  inv1  gate812(.a(N165), .O(gate207inter8));
  nand2 gate813(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate814(.a(s_61), .b(gate207inter3), .O(gate207inter10));
  nor2  gate815(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate816(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate817(.a(gate207inter12), .b(gate207inter1), .O(N597));
or2 gate208( .a(N557), .b(N165), .O(N600) );
and2 gate209( .a(N246), .b(N557), .O(N605) );
nand2 gate210( .a(N561), .b(N171), .O(N606) );
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );

  xor2  gate916(.a(N177), .b(N565), .O(gate213inter0));
  nand2 gate917(.a(gate213inter0), .b(s_76), .O(gate213inter1));
  and2  gate918(.a(N177), .b(N565), .O(gate213inter2));
  inv1  gate919(.a(s_76), .O(gate213inter3));
  inv1  gate920(.a(s_77), .O(gate213inter4));
  nand2 gate921(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate922(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate923(.a(N565), .O(gate213inter7));
  inv1  gate924(.a(N177), .O(gate213inter8));
  nand2 gate925(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate926(.a(s_77), .b(gate213inter3), .O(gate213inter10));
  nor2  gate927(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate928(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate929(.a(gate213inter12), .b(gate213inter1), .O(N616));
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );
nand2 gate216( .a(N569), .b(N183), .O(N625) );
or2 gate217( .a(N569), .b(N183), .O(N628) );
and2 gate218( .a(N246), .b(N569), .O(N631) );

  xor2  gate678(.a(N189), .b(N573), .O(gate219inter0));
  nand2 gate679(.a(gate219inter0), .b(s_42), .O(gate219inter1));
  and2  gate680(.a(N189), .b(N573), .O(gate219inter2));
  inv1  gate681(.a(s_42), .O(gate219inter3));
  inv1  gate682(.a(s_43), .O(gate219inter4));
  nand2 gate683(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate684(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate685(.a(N573), .O(gate219inter7));
  inv1  gate686(.a(N189), .O(gate219inter8));
  nand2 gate687(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate688(.a(s_43), .b(gate219inter3), .O(gate219inter10));
  nor2  gate689(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate690(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate691(.a(gate219inter12), .b(gate219inter1), .O(N632));
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );

  xor2  gate846(.a(N195), .b(N577), .O(gate222inter0));
  nand2 gate847(.a(gate222inter0), .b(s_66), .O(gate222inter1));
  and2  gate848(.a(N195), .b(N577), .O(gate222inter2));
  inv1  gate849(.a(s_66), .O(gate222inter3));
  inv1  gate850(.a(s_67), .O(gate222inter4));
  nand2 gate851(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate852(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate853(.a(N577), .O(gate222inter7));
  inv1  gate854(.a(N195), .O(gate222inter8));
  nand2 gate855(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate856(.a(s_67), .b(gate222inter3), .O(gate222inter10));
  nor2  gate857(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate858(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate859(.a(gate222inter12), .b(gate222inter1), .O(N641));
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );
nand2 gate225( .a(N581), .b(N201), .O(N651) );
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );

  xor2  gate468(.a(N588), .b(N552), .O(gate228inter0));
  nand2 gate469(.a(gate228inter0), .b(s_12), .O(gate228inter1));
  and2  gate470(.a(N588), .b(N552), .O(gate228inter2));
  inv1  gate471(.a(s_12), .O(gate228inter3));
  inv1  gate472(.a(s_13), .O(gate228inter4));
  nand2 gate473(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate474(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate475(.a(N552), .O(gate228inter7));
  inv1  gate476(.a(N588), .O(gate228inter8));
  nand2 gate477(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate478(.a(s_13), .b(gate228inter3), .O(gate228inter10));
  nor2  gate479(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate480(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate481(.a(gate228inter12), .b(gate228inter1), .O(N660));
nor2 gate229( .a(N587), .b(N589), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
and2 gate231( .a(N593), .b(N590), .O(N665) );
nor2 gate232( .a(N596), .b(N522), .O(N669) );
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );
nor2 gate235( .a(N605), .b(N523), .O(N677) );
inv1 gate236( .a(N606), .O(N678) );
and2 gate237( .a(N609), .b(N606), .O(N682) );

  xor2  gate832(.a(N524), .b(N615), .O(gate238inter0));
  nand2 gate833(.a(gate238inter0), .b(s_64), .O(gate238inter1));
  and2  gate834(.a(N524), .b(N615), .O(gate238inter2));
  inv1  gate835(.a(s_64), .O(gate238inter3));
  inv1  gate836(.a(s_65), .O(gate238inter4));
  nand2 gate837(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate838(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate839(.a(N615), .O(gate238inter7));
  inv1  gate840(.a(N524), .O(gate238inter8));
  nand2 gate841(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate842(.a(s_65), .b(gate238inter3), .O(gate238inter10));
  nor2  gate843(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate844(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate845(.a(gate238inter12), .b(gate238inter1), .O(N686));
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );

  xor2  gate482(.a(N525), .b(N624), .O(gate241inter0));
  nand2 gate483(.a(gate241inter0), .b(s_14), .O(gate241inter1));
  and2  gate484(.a(N525), .b(N624), .O(gate241inter2));
  inv1  gate485(.a(s_14), .O(gate241inter3));
  inv1  gate486(.a(s_15), .O(gate241inter4));
  nand2 gate487(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate488(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate489(.a(N624), .O(gate241inter7));
  inv1  gate490(.a(N525), .O(gate241inter8));
  nand2 gate491(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate492(.a(s_15), .b(gate241inter3), .O(gate241inter10));
  nor2  gate493(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate494(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate495(.a(gate241inter12), .b(gate241inter1), .O(N696));
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );
nor2 gate244( .a(N631), .b(N526), .O(N704) );
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );
nor2 gate247( .a(N337), .b(N640), .O(N712) );
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );
nor2 gate250( .a(N339), .b(N650), .O(N721) );
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );
nor2 gate253( .a(N341), .b(N659), .O(N731) );
nand2 gate254( .a(N654), .b(N261), .O(N732) );
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
and2 gate273( .a(N228), .b(N708), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );
nor2 gate279( .a(N727), .b(N261), .O(N757) );
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );

  xor2  gate762(.a(N713), .b(N635), .O(gate284inter0));
  nand2 gate763(.a(gate284inter0), .b(s_54), .O(gate284inter1));
  and2  gate764(.a(N713), .b(N635), .O(gate284inter2));
  inv1  gate765(.a(s_54), .O(gate284inter3));
  inv1  gate766(.a(s_55), .O(gate284inter4));
  nand2 gate767(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate768(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate769(.a(N635), .O(gate284inter7));
  inv1  gate770(.a(N713), .O(gate284inter8));
  nand2 gate771(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate772(.a(s_55), .b(gate284inter3), .O(gate284inter10));
  nor2  gate773(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate774(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate775(.a(gate284inter12), .b(gate284inter1), .O(N762));
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );
nor2 gate291( .a(N736), .b(N737), .O(N769) );

  xor2  gate874(.a(N740), .b(N739), .O(gate292inter0));
  nand2 gate875(.a(gate292inter0), .b(s_70), .O(gate292inter1));
  and2  gate876(.a(N740), .b(N739), .O(gate292inter2));
  inv1  gate877(.a(s_70), .O(gate292inter3));
  inv1  gate878(.a(s_71), .O(gate292inter4));
  nand2 gate879(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate880(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate881(.a(N739), .O(gate292inter7));
  inv1  gate882(.a(N740), .O(gate292inter8));
  nand2 gate883(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate884(.a(s_71), .b(gate292inter3), .O(gate292inter10));
  nor2  gate885(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate886(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate887(.a(gate292inter12), .b(gate292inter1), .O(N770));
nor2 gate293( .a(N742), .b(N743), .O(N771) );
nor2 gate294( .a(N745), .b(N746), .O(N772) );
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );
nor2 gate296( .a(N748), .b(N749), .O(N777) );
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );
nor2 gate298( .a(N751), .b(N752), .O(N781) );
nand2 gate299( .a(N756), .b(N732), .O(N782) );

  xor2  gate860(.a(N755), .b(N754), .O(gate300inter0));
  nand2 gate861(.a(gate300inter0), .b(s_68), .O(gate300inter1));
  and2  gate862(.a(N755), .b(N754), .O(gate300inter2));
  inv1  gate863(.a(s_68), .O(gate300inter3));
  inv1  gate864(.a(s_69), .O(gate300inter4));
  nand2 gate865(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate866(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate867(.a(N754), .O(gate300inter7));
  inv1  gate868(.a(N755), .O(gate300inter8));
  nand2 gate869(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate870(.a(s_69), .b(gate300inter3), .O(gate300inter10));
  nor2  gate871(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate872(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate873(.a(gate300inter12), .b(gate300inter1), .O(N785));
nor2 gate301( .a(N757), .b(N758), .O(N786) );

  xor2  gate734(.a(N760), .b(N759), .O(gate302inter0));
  nand2 gate735(.a(gate302inter0), .b(s_50), .O(gate302inter1));
  and2  gate736(.a(N760), .b(N759), .O(gate302inter2));
  inv1  gate737(.a(s_50), .O(gate302inter3));
  inv1  gate738(.a(s_51), .O(gate302inter4));
  nand2 gate739(.a(gate302inter4), .b(gate302inter3), .O(gate302inter5));
  nor2  gate740(.a(gate302inter5), .b(gate302inter2), .O(gate302inter6));
  inv1  gate741(.a(N759), .O(gate302inter7));
  inv1  gate742(.a(N760), .O(gate302inter8));
  nand2 gate743(.a(gate302inter8), .b(gate302inter7), .O(gate302inter9));
  nand2 gate744(.a(s_51), .b(gate302inter3), .O(gate302inter10));
  nor2  gate745(.a(gate302inter10), .b(gate302inter9), .O(gate302inter11));
  nor2  gate746(.a(gate302inter11), .b(gate302inter6), .O(gate302inter12));
  nand2 gate747(.a(gate302inter12), .b(gate302inter1), .O(N787));
nor2 gate303( .a(N700), .b(N773), .O(N788) );
and2 gate304( .a(N700), .b(N773), .O(N789) );
nor2 gate305( .a(N708), .b(N778), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );

  xor2  gate692(.a(N782), .b(N717), .O(gate307inter0));
  nand2 gate693(.a(gate307inter0), .b(s_44), .O(gate307inter1));
  and2  gate694(.a(N782), .b(N717), .O(gate307inter2));
  inv1  gate695(.a(s_44), .O(gate307inter3));
  inv1  gate696(.a(s_45), .O(gate307inter4));
  nand2 gate697(.a(gate307inter4), .b(gate307inter3), .O(gate307inter5));
  nor2  gate698(.a(gate307inter5), .b(gate307inter2), .O(gate307inter6));
  inv1  gate699(.a(N717), .O(gate307inter7));
  inv1  gate700(.a(N782), .O(gate307inter8));
  nand2 gate701(.a(gate307inter8), .b(gate307inter7), .O(gate307inter9));
  nand2 gate702(.a(s_45), .b(gate307inter3), .O(gate307inter10));
  nor2  gate703(.a(gate307inter10), .b(gate307inter9), .O(gate307inter11));
  nor2  gate704(.a(gate307inter11), .b(gate307inter6), .O(gate307inter12));
  nand2 gate705(.a(gate307inter12), .b(gate307inter1), .O(N792));
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );
nand2 gate310( .a(N628), .b(N773), .O(N795) );

  xor2  gate454(.a(N747), .b(N795), .O(gate311inter0));
  nand2 gate455(.a(gate311inter0), .b(s_10), .O(gate311inter1));
  and2  gate456(.a(N747), .b(N795), .O(gate311inter2));
  inv1  gate457(.a(s_10), .O(gate311inter3));
  inv1  gate458(.a(s_11), .O(gate311inter4));
  nand2 gate459(.a(gate311inter4), .b(gate311inter3), .O(gate311inter5));
  nor2  gate460(.a(gate311inter5), .b(gate311inter2), .O(gate311inter6));
  inv1  gate461(.a(N795), .O(gate311inter7));
  inv1  gate462(.a(N747), .O(gate311inter8));
  nand2 gate463(.a(gate311inter8), .b(gate311inter7), .O(gate311inter9));
  nand2 gate464(.a(s_11), .b(gate311inter3), .O(gate311inter10));
  nor2  gate465(.a(gate311inter10), .b(gate311inter9), .O(gate311inter11));
  nor2  gate466(.a(gate311inter11), .b(gate311inter6), .O(gate311inter12));
  nand2 gate467(.a(gate311inter12), .b(gate311inter1), .O(N796));
nor2 gate312( .a(N788), .b(N789), .O(N802) );
nor2 gate313( .a(N790), .b(N791), .O(N803) );
nor2 gate314( .a(N792), .b(N793), .O(N804) );

  xor2  gate594(.a(N794), .b(N340), .O(gate315inter0));
  nand2 gate595(.a(gate315inter0), .b(s_30), .O(gate315inter1));
  and2  gate596(.a(N794), .b(N340), .O(gate315inter2));
  inv1  gate597(.a(s_30), .O(gate315inter3));
  inv1  gate598(.a(s_31), .O(gate315inter4));
  nand2 gate599(.a(gate315inter4), .b(gate315inter3), .O(gate315inter5));
  nor2  gate600(.a(gate315inter5), .b(gate315inter2), .O(gate315inter6));
  inv1  gate601(.a(N340), .O(gate315inter7));
  inv1  gate602(.a(N794), .O(gate315inter8));
  nand2 gate603(.a(gate315inter8), .b(gate315inter7), .O(gate315inter9));
  nand2 gate604(.a(s_31), .b(gate315inter3), .O(gate315inter10));
  nor2  gate605(.a(gate315inter10), .b(gate315inter9), .O(gate315inter11));
  nor2  gate606(.a(gate315inter11), .b(gate315inter6), .O(gate315inter12));
  nand2 gate607(.a(gate315inter12), .b(gate315inter1), .O(N805));

  xor2  gate538(.a(N796), .b(N692), .O(gate316inter0));
  nand2 gate539(.a(gate316inter0), .b(s_22), .O(gate316inter1));
  and2  gate540(.a(N796), .b(N692), .O(gate316inter2));
  inv1  gate541(.a(s_22), .O(gate316inter3));
  inv1  gate542(.a(s_23), .O(gate316inter4));
  nand2 gate543(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate544(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate545(.a(N692), .O(gate316inter7));
  inv1  gate546(.a(N796), .O(gate316inter8));
  nand2 gate547(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate548(.a(s_23), .b(gate316inter3), .O(gate316inter10));
  nor2  gate549(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate550(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate551(.a(gate316inter12), .b(gate316inter1), .O(N806));
and2 gate317( .a(N692), .b(N796), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );

  xor2  gate664(.a(N796), .b(N619), .O(gate322inter0));
  nand2 gate665(.a(gate322inter0), .b(s_40), .O(gate322inter1));
  and2  gate666(.a(N796), .b(N619), .O(gate322inter2));
  inv1  gate667(.a(s_40), .O(gate322inter3));
  inv1  gate668(.a(s_41), .O(gate322inter4));
  nand2 gate669(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate670(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate671(.a(N619), .O(gate322inter7));
  inv1  gate672(.a(N796), .O(gate322inter8));
  nand2 gate673(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate674(.a(s_41), .b(gate322inter3), .O(gate322inter10));
  nor2  gate675(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate676(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate677(.a(gate322inter12), .b(gate322inter1), .O(N812));
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );

  xor2  gate636(.a(N812), .b(N744), .O(gate327inter0));
  nand2 gate637(.a(gate327inter0), .b(s_36), .O(gate327inter1));
  and2  gate638(.a(N812), .b(N744), .O(gate327inter2));
  inv1  gate639(.a(s_36), .O(gate327inter3));
  inv1  gate640(.a(s_37), .O(gate327inter4));
  nand2 gate641(.a(gate327inter4), .b(gate327inter3), .O(gate327inter5));
  nor2  gate642(.a(gate327inter5), .b(gate327inter2), .O(gate327inter6));
  inv1  gate643(.a(N744), .O(gate327inter7));
  inv1  gate644(.a(N812), .O(gate327inter8));
  nand2 gate645(.a(gate327inter8), .b(gate327inter7), .O(gate327inter9));
  nand2 gate646(.a(s_37), .b(gate327inter3), .O(gate327inter10));
  nor2  gate647(.a(gate327inter10), .b(gate327inter9), .O(gate327inter11));
  nor2  gate648(.a(gate327inter11), .b(gate327inter6), .O(gate327inter12));
  nand2 gate649(.a(gate327inter12), .b(gate327inter1), .O(N822));

  xor2  gate748(.a(N807), .b(N806), .O(gate328inter0));
  nand2 gate749(.a(gate328inter0), .b(s_52), .O(gate328inter1));
  and2  gate750(.a(N807), .b(N806), .O(gate328inter2));
  inv1  gate751(.a(s_52), .O(gate328inter3));
  inv1  gate752(.a(s_53), .O(gate328inter4));
  nand2 gate753(.a(gate328inter4), .b(gate328inter3), .O(gate328inter5));
  nor2  gate754(.a(gate328inter5), .b(gate328inter2), .O(gate328inter6));
  inv1  gate755(.a(N806), .O(gate328inter7));
  inv1  gate756(.a(N807), .O(gate328inter8));
  nand2 gate757(.a(gate328inter8), .b(gate328inter7), .O(gate328inter9));
  nand2 gate758(.a(s_53), .b(gate328inter3), .O(gate328inter10));
  nor2  gate759(.a(gate328inter10), .b(gate328inter9), .O(gate328inter11));
  nor2  gate760(.a(gate328inter11), .b(gate328inter6), .O(gate328inter12));
  nand2 gate761(.a(gate328inter12), .b(gate328inter1), .O(N825));
nor2 gate329( .a(N335), .b(N808), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );
nor2 gate333( .a(N665), .b(N815), .O(N830) );
and2 gate334( .a(N665), .b(N815), .O(N831) );
nor2 gate335( .a(N673), .b(N819), .O(N832) );
and2 gate336( .a(N673), .b(N819), .O(N833) );
nor2 gate337( .a(N682), .b(N822), .O(N834) );
and2 gate338( .a(N682), .b(N822), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );

  xor2  gate398(.a(N593), .b(N815), .O(gate344inter0));
  nand2 gate399(.a(gate344inter0), .b(s_2), .O(gate344inter1));
  and2  gate400(.a(N593), .b(N815), .O(gate344inter2));
  inv1  gate401(.a(s_2), .O(gate344inter3));
  inv1  gate402(.a(s_3), .O(gate344inter4));
  nand2 gate403(.a(gate344inter4), .b(gate344inter3), .O(gate344inter5));
  nor2  gate404(.a(gate344inter5), .b(gate344inter2), .O(gate344inter6));
  inv1  gate405(.a(N815), .O(gate344inter7));
  inv1  gate406(.a(N593), .O(gate344inter8));
  nand2 gate407(.a(gate344inter8), .b(gate344inter7), .O(gate344inter9));
  nand2 gate408(.a(s_3), .b(gate344inter3), .O(gate344inter10));
  nor2  gate409(.a(gate344inter10), .b(gate344inter9), .O(gate344inter11));
  nor2  gate410(.a(gate344inter11), .b(gate344inter6), .O(gate344inter12));
  nand2 gate411(.a(gate344inter12), .b(gate344inter1), .O(N841));
nor2 gate345( .a(N830), .b(N831), .O(N842) );
nor2 gate346( .a(N832), .b(N833), .O(N843) );

  xor2  gate790(.a(N835), .b(N834), .O(gate347inter0));
  nand2 gate791(.a(gate347inter0), .b(s_58), .O(gate347inter1));
  and2  gate792(.a(N835), .b(N834), .O(gate347inter2));
  inv1  gate793(.a(s_58), .O(gate347inter3));
  inv1  gate794(.a(s_59), .O(gate347inter4));
  nand2 gate795(.a(gate347inter4), .b(gate347inter3), .O(gate347inter5));
  nor2  gate796(.a(gate347inter5), .b(gate347inter2), .O(gate347inter6));
  inv1  gate797(.a(N834), .O(gate347inter7));
  inv1  gate798(.a(N835), .O(gate347inter8));
  nand2 gate799(.a(gate347inter8), .b(gate347inter7), .O(gate347inter9));
  nand2 gate800(.a(s_59), .b(gate347inter3), .O(gate347inter10));
  nor2  gate801(.a(gate347inter10), .b(gate347inter9), .O(gate347inter11));
  nor2  gate802(.a(gate347inter11), .b(gate347inter6), .O(gate347inter12));
  nand2 gate803(.a(gate347inter12), .b(gate347inter1), .O(N844));

  xor2  gate384(.a(N836), .b(N334), .O(gate348inter0));
  nand2 gate385(.a(gate348inter0), .b(s_0), .O(gate348inter1));
  and2  gate386(.a(N836), .b(N334), .O(gate348inter2));
  inv1  gate387(.a(s_0), .O(gate348inter3));
  inv1  gate388(.a(s_1), .O(gate348inter4));
  nand2 gate389(.a(gate348inter4), .b(gate348inter3), .O(gate348inter5));
  nor2  gate390(.a(gate348inter5), .b(gate348inter2), .O(gate348inter6));
  inv1  gate391(.a(N334), .O(gate348inter7));
  inv1  gate392(.a(N836), .O(gate348inter8));
  nand2 gate393(.a(gate348inter8), .b(gate348inter7), .O(gate348inter9));
  nand2 gate394(.a(s_1), .b(gate348inter3), .O(gate348inter10));
  nor2  gate395(.a(gate348inter10), .b(gate348inter9), .O(gate348inter11));
  nor2  gate396(.a(gate348inter11), .b(gate348inter6), .O(gate348inter12));
  nand2 gate397(.a(gate348inter12), .b(gate348inter1), .O(N845));
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
and2 gate354( .a(N219), .b(N842), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );
nor2 gate362( .a(N417), .b(N851), .O(N859) );
nor2 gate363( .a(N332), .b(N852), .O(N860) );
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

endmodule