module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1135(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1136(.a(gate12inter0), .b(s_84), .O(gate12inter1));
  and2  gate1137(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1138(.a(s_84), .O(gate12inter3));
  inv1  gate1139(.a(s_85), .O(gate12inter4));
  nand2 gate1140(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1141(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1142(.a(G7), .O(gate12inter7));
  inv1  gate1143(.a(G8), .O(gate12inter8));
  nand2 gate1144(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1145(.a(s_85), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1146(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1147(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1148(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1919(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1920(.a(gate20inter0), .b(s_196), .O(gate20inter1));
  and2  gate1921(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1922(.a(s_196), .O(gate20inter3));
  inv1  gate1923(.a(s_197), .O(gate20inter4));
  nand2 gate1924(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1925(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1926(.a(G23), .O(gate20inter7));
  inv1  gate1927(.a(G24), .O(gate20inter8));
  nand2 gate1928(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1929(.a(s_197), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1930(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1931(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1932(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate855(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate856(.a(gate21inter0), .b(s_44), .O(gate21inter1));
  and2  gate857(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate858(.a(s_44), .O(gate21inter3));
  inv1  gate859(.a(s_45), .O(gate21inter4));
  nand2 gate860(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate861(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate862(.a(G25), .O(gate21inter7));
  inv1  gate863(.a(G26), .O(gate21inter8));
  nand2 gate864(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate865(.a(s_45), .b(gate21inter3), .O(gate21inter10));
  nor2  gate866(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate867(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate868(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate589(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate590(.a(gate23inter0), .b(s_6), .O(gate23inter1));
  and2  gate591(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate592(.a(s_6), .O(gate23inter3));
  inv1  gate593(.a(s_7), .O(gate23inter4));
  nand2 gate594(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate595(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate596(.a(G29), .O(gate23inter7));
  inv1  gate597(.a(G30), .O(gate23inter8));
  nand2 gate598(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate599(.a(s_7), .b(gate23inter3), .O(gate23inter10));
  nor2  gate600(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate601(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate602(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1527(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1528(.a(gate24inter0), .b(s_140), .O(gate24inter1));
  and2  gate1529(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1530(.a(s_140), .O(gate24inter3));
  inv1  gate1531(.a(s_141), .O(gate24inter4));
  nand2 gate1532(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1533(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1534(.a(G31), .O(gate24inter7));
  inv1  gate1535(.a(G32), .O(gate24inter8));
  nand2 gate1536(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1537(.a(s_141), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1538(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1539(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1540(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate2059(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2060(.a(gate25inter0), .b(s_216), .O(gate25inter1));
  and2  gate2061(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2062(.a(s_216), .O(gate25inter3));
  inv1  gate2063(.a(s_217), .O(gate25inter4));
  nand2 gate2064(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2065(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2066(.a(G1), .O(gate25inter7));
  inv1  gate2067(.a(G5), .O(gate25inter8));
  nand2 gate2068(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2069(.a(s_217), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2070(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2071(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2072(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate967(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate968(.a(gate26inter0), .b(s_60), .O(gate26inter1));
  and2  gate969(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate970(.a(s_60), .O(gate26inter3));
  inv1  gate971(.a(s_61), .O(gate26inter4));
  nand2 gate972(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate973(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate974(.a(G9), .O(gate26inter7));
  inv1  gate975(.a(G13), .O(gate26inter8));
  nand2 gate976(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate977(.a(s_61), .b(gate26inter3), .O(gate26inter10));
  nor2  gate978(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate979(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate980(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1989(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1990(.a(gate29inter0), .b(s_206), .O(gate29inter1));
  and2  gate1991(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1992(.a(s_206), .O(gate29inter3));
  inv1  gate1993(.a(s_207), .O(gate29inter4));
  nand2 gate1994(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1995(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1996(.a(G3), .O(gate29inter7));
  inv1  gate1997(.a(G7), .O(gate29inter8));
  nand2 gate1998(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1999(.a(s_207), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2000(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2001(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2002(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1933(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1934(.a(gate33inter0), .b(s_198), .O(gate33inter1));
  and2  gate1935(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1936(.a(s_198), .O(gate33inter3));
  inv1  gate1937(.a(s_199), .O(gate33inter4));
  nand2 gate1938(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1939(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1940(.a(G17), .O(gate33inter7));
  inv1  gate1941(.a(G21), .O(gate33inter8));
  nand2 gate1942(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1943(.a(s_199), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1944(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1945(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1946(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1303(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1304(.a(gate35inter0), .b(s_108), .O(gate35inter1));
  and2  gate1305(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1306(.a(s_108), .O(gate35inter3));
  inv1  gate1307(.a(s_109), .O(gate35inter4));
  nand2 gate1308(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1309(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1310(.a(G18), .O(gate35inter7));
  inv1  gate1311(.a(G22), .O(gate35inter8));
  nand2 gate1312(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1313(.a(s_109), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1314(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1315(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1316(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1233(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1234(.a(gate38inter0), .b(s_98), .O(gate38inter1));
  and2  gate1235(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1236(.a(s_98), .O(gate38inter3));
  inv1  gate1237(.a(s_99), .O(gate38inter4));
  nand2 gate1238(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1239(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1240(.a(G27), .O(gate38inter7));
  inv1  gate1241(.a(G31), .O(gate38inter8));
  nand2 gate1242(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1243(.a(s_99), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1244(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1245(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1246(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate701(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate702(.a(gate39inter0), .b(s_22), .O(gate39inter1));
  and2  gate703(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate704(.a(s_22), .O(gate39inter3));
  inv1  gate705(.a(s_23), .O(gate39inter4));
  nand2 gate706(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate707(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate708(.a(G20), .O(gate39inter7));
  inv1  gate709(.a(G24), .O(gate39inter8));
  nand2 gate710(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate711(.a(s_23), .b(gate39inter3), .O(gate39inter10));
  nor2  gate712(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate713(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate714(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate687(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate688(.a(gate40inter0), .b(s_20), .O(gate40inter1));
  and2  gate689(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate690(.a(s_20), .O(gate40inter3));
  inv1  gate691(.a(s_21), .O(gate40inter4));
  nand2 gate692(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate693(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate694(.a(G28), .O(gate40inter7));
  inv1  gate695(.a(G32), .O(gate40inter8));
  nand2 gate696(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate697(.a(s_21), .b(gate40inter3), .O(gate40inter10));
  nor2  gate698(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate699(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate700(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate995(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate996(.a(gate43inter0), .b(s_64), .O(gate43inter1));
  and2  gate997(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate998(.a(s_64), .O(gate43inter3));
  inv1  gate999(.a(s_65), .O(gate43inter4));
  nand2 gate1000(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1001(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1002(.a(G3), .O(gate43inter7));
  inv1  gate1003(.a(G269), .O(gate43inter8));
  nand2 gate1004(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1005(.a(s_65), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1006(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1007(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1008(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1023(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1024(.a(gate44inter0), .b(s_68), .O(gate44inter1));
  and2  gate1025(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1026(.a(s_68), .O(gate44inter3));
  inv1  gate1027(.a(s_69), .O(gate44inter4));
  nand2 gate1028(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1029(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1030(.a(G4), .O(gate44inter7));
  inv1  gate1031(.a(G269), .O(gate44inter8));
  nand2 gate1032(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1033(.a(s_69), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1034(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1035(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1036(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1037(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1038(.a(gate45inter0), .b(s_70), .O(gate45inter1));
  and2  gate1039(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1040(.a(s_70), .O(gate45inter3));
  inv1  gate1041(.a(s_71), .O(gate45inter4));
  nand2 gate1042(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1043(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1044(.a(G5), .O(gate45inter7));
  inv1  gate1045(.a(G272), .O(gate45inter8));
  nand2 gate1046(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1047(.a(s_71), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1048(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1049(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1050(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2311(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2312(.a(gate48inter0), .b(s_252), .O(gate48inter1));
  and2  gate2313(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2314(.a(s_252), .O(gate48inter3));
  inv1  gate2315(.a(s_253), .O(gate48inter4));
  nand2 gate2316(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2317(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2318(.a(G8), .O(gate48inter7));
  inv1  gate2319(.a(G275), .O(gate48inter8));
  nand2 gate2320(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2321(.a(s_253), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2322(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2323(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2324(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate603(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate604(.a(gate50inter0), .b(s_8), .O(gate50inter1));
  and2  gate605(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate606(.a(s_8), .O(gate50inter3));
  inv1  gate607(.a(s_9), .O(gate50inter4));
  nand2 gate608(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate609(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate610(.a(G10), .O(gate50inter7));
  inv1  gate611(.a(G278), .O(gate50inter8));
  nand2 gate612(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate613(.a(s_9), .b(gate50inter3), .O(gate50inter10));
  nor2  gate614(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate615(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate616(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2199(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2200(.a(gate56inter0), .b(s_236), .O(gate56inter1));
  and2  gate2201(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2202(.a(s_236), .O(gate56inter3));
  inv1  gate2203(.a(s_237), .O(gate56inter4));
  nand2 gate2204(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2205(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2206(.a(G16), .O(gate56inter7));
  inv1  gate2207(.a(G287), .O(gate56inter8));
  nand2 gate2208(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2209(.a(s_237), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2210(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2211(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2212(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1275(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1276(.a(gate61inter0), .b(s_104), .O(gate61inter1));
  and2  gate1277(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1278(.a(s_104), .O(gate61inter3));
  inv1  gate1279(.a(s_105), .O(gate61inter4));
  nand2 gate1280(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1281(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1282(.a(G21), .O(gate61inter7));
  inv1  gate1283(.a(G296), .O(gate61inter8));
  nand2 gate1284(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1285(.a(s_105), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1286(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1287(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1288(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1443(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1444(.a(gate62inter0), .b(s_128), .O(gate62inter1));
  and2  gate1445(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1446(.a(s_128), .O(gate62inter3));
  inv1  gate1447(.a(s_129), .O(gate62inter4));
  nand2 gate1448(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1449(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1450(.a(G22), .O(gate62inter7));
  inv1  gate1451(.a(G296), .O(gate62inter8));
  nand2 gate1452(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1453(.a(s_129), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1454(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1455(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1456(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate743(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate744(.a(gate64inter0), .b(s_28), .O(gate64inter1));
  and2  gate745(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate746(.a(s_28), .O(gate64inter3));
  inv1  gate747(.a(s_29), .O(gate64inter4));
  nand2 gate748(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate749(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate750(.a(G24), .O(gate64inter7));
  inv1  gate751(.a(G299), .O(gate64inter8));
  nand2 gate752(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate753(.a(s_29), .b(gate64inter3), .O(gate64inter10));
  nor2  gate754(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate755(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate756(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2185(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2186(.a(gate67inter0), .b(s_234), .O(gate67inter1));
  and2  gate2187(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2188(.a(s_234), .O(gate67inter3));
  inv1  gate2189(.a(s_235), .O(gate67inter4));
  nand2 gate2190(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2191(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2192(.a(G27), .O(gate67inter7));
  inv1  gate2193(.a(G305), .O(gate67inter8));
  nand2 gate2194(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2195(.a(s_235), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2196(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2197(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2198(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1611(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1612(.a(gate79inter0), .b(s_152), .O(gate79inter1));
  and2  gate1613(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1614(.a(s_152), .O(gate79inter3));
  inv1  gate1615(.a(s_153), .O(gate79inter4));
  nand2 gate1616(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1617(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1618(.a(G10), .O(gate79inter7));
  inv1  gate1619(.a(G323), .O(gate79inter8));
  nand2 gate1620(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1621(.a(s_153), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1622(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1623(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1624(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate575(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate576(.a(gate80inter0), .b(s_4), .O(gate80inter1));
  and2  gate577(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate578(.a(s_4), .O(gate80inter3));
  inv1  gate579(.a(s_5), .O(gate80inter4));
  nand2 gate580(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate581(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate582(.a(G14), .O(gate80inter7));
  inv1  gate583(.a(G323), .O(gate80inter8));
  nand2 gate584(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate585(.a(s_5), .b(gate80inter3), .O(gate80inter10));
  nor2  gate586(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate587(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate588(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2129(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2130(.a(gate82inter0), .b(s_226), .O(gate82inter1));
  and2  gate2131(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2132(.a(s_226), .O(gate82inter3));
  inv1  gate2133(.a(s_227), .O(gate82inter4));
  nand2 gate2134(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2135(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2136(.a(G7), .O(gate82inter7));
  inv1  gate2137(.a(G326), .O(gate82inter8));
  nand2 gate2138(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2139(.a(s_227), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2140(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2141(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2142(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1163(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1164(.a(gate83inter0), .b(s_88), .O(gate83inter1));
  and2  gate1165(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1166(.a(s_88), .O(gate83inter3));
  inv1  gate1167(.a(s_89), .O(gate83inter4));
  nand2 gate1168(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1169(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1170(.a(G11), .O(gate83inter7));
  inv1  gate1171(.a(G329), .O(gate83inter8));
  nand2 gate1172(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1173(.a(s_89), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1174(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1175(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1176(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1807(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1808(.a(gate88inter0), .b(s_180), .O(gate88inter1));
  and2  gate1809(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1810(.a(s_180), .O(gate88inter3));
  inv1  gate1811(.a(s_181), .O(gate88inter4));
  nand2 gate1812(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1813(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1814(.a(G16), .O(gate88inter7));
  inv1  gate1815(.a(G335), .O(gate88inter8));
  nand2 gate1816(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1817(.a(s_181), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1818(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1819(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1820(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2115(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2116(.a(gate89inter0), .b(s_224), .O(gate89inter1));
  and2  gate2117(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2118(.a(s_224), .O(gate89inter3));
  inv1  gate2119(.a(s_225), .O(gate89inter4));
  nand2 gate2120(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2121(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2122(.a(G17), .O(gate89inter7));
  inv1  gate2123(.a(G338), .O(gate89inter8));
  nand2 gate2124(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2125(.a(s_225), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2126(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2127(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2128(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate1681(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1682(.a(gate90inter0), .b(s_162), .O(gate90inter1));
  and2  gate1683(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1684(.a(s_162), .O(gate90inter3));
  inv1  gate1685(.a(s_163), .O(gate90inter4));
  nand2 gate1686(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1687(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1688(.a(G21), .O(gate90inter7));
  inv1  gate1689(.a(G338), .O(gate90inter8));
  nand2 gate1690(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1691(.a(s_163), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1692(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1693(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1694(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate715(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate716(.a(gate91inter0), .b(s_24), .O(gate91inter1));
  and2  gate717(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate718(.a(s_24), .O(gate91inter3));
  inv1  gate719(.a(s_25), .O(gate91inter4));
  nand2 gate720(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate721(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate722(.a(G25), .O(gate91inter7));
  inv1  gate723(.a(G341), .O(gate91inter8));
  nand2 gate724(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate725(.a(s_25), .b(gate91inter3), .O(gate91inter10));
  nor2  gate726(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate727(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate728(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1065(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1066(.a(gate92inter0), .b(s_74), .O(gate92inter1));
  and2  gate1067(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1068(.a(s_74), .O(gate92inter3));
  inv1  gate1069(.a(s_75), .O(gate92inter4));
  nand2 gate1070(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1071(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1072(.a(G29), .O(gate92inter7));
  inv1  gate1073(.a(G341), .O(gate92inter8));
  nand2 gate1074(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1075(.a(s_75), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1076(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1077(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1078(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2339(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2340(.a(gate94inter0), .b(s_256), .O(gate94inter1));
  and2  gate2341(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2342(.a(s_256), .O(gate94inter3));
  inv1  gate2343(.a(s_257), .O(gate94inter4));
  nand2 gate2344(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2345(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2346(.a(G22), .O(gate94inter7));
  inv1  gate2347(.a(G344), .O(gate94inter8));
  nand2 gate2348(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2349(.a(s_257), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2350(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2351(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2352(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1513(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1514(.a(gate95inter0), .b(s_138), .O(gate95inter1));
  and2  gate1515(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1516(.a(s_138), .O(gate95inter3));
  inv1  gate1517(.a(s_139), .O(gate95inter4));
  nand2 gate1518(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1519(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1520(.a(G26), .O(gate95inter7));
  inv1  gate1521(.a(G347), .O(gate95inter8));
  nand2 gate1522(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1523(.a(s_139), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1524(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1525(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1526(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1877(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1878(.a(gate98inter0), .b(s_190), .O(gate98inter1));
  and2  gate1879(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1880(.a(s_190), .O(gate98inter3));
  inv1  gate1881(.a(s_191), .O(gate98inter4));
  nand2 gate1882(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1883(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1884(.a(G23), .O(gate98inter7));
  inv1  gate1885(.a(G350), .O(gate98inter8));
  nand2 gate1886(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1887(.a(s_191), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1888(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1889(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1890(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1849(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1850(.a(gate103inter0), .b(s_186), .O(gate103inter1));
  and2  gate1851(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1852(.a(s_186), .O(gate103inter3));
  inv1  gate1853(.a(s_187), .O(gate103inter4));
  nand2 gate1854(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1855(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1856(.a(G28), .O(gate103inter7));
  inv1  gate1857(.a(G359), .O(gate103inter8));
  nand2 gate1858(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1859(.a(s_187), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1860(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1861(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1862(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate869(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate870(.a(gate104inter0), .b(s_46), .O(gate104inter1));
  and2  gate871(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate872(.a(s_46), .O(gate104inter3));
  inv1  gate873(.a(s_47), .O(gate104inter4));
  nand2 gate874(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate875(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate876(.a(G32), .O(gate104inter7));
  inv1  gate877(.a(G359), .O(gate104inter8));
  nand2 gate878(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate879(.a(s_47), .b(gate104inter3), .O(gate104inter10));
  nor2  gate880(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate881(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate882(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2017(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2018(.a(gate106inter0), .b(s_210), .O(gate106inter1));
  and2  gate2019(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2020(.a(s_210), .O(gate106inter3));
  inv1  gate2021(.a(s_211), .O(gate106inter4));
  nand2 gate2022(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2023(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2024(.a(G364), .O(gate106inter7));
  inv1  gate2025(.a(G365), .O(gate106inter8));
  nand2 gate2026(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2027(.a(s_211), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2028(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2029(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2030(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1191(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1192(.a(gate108inter0), .b(s_92), .O(gate108inter1));
  and2  gate1193(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1194(.a(s_92), .O(gate108inter3));
  inv1  gate1195(.a(s_93), .O(gate108inter4));
  nand2 gate1196(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1197(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1198(.a(G368), .O(gate108inter7));
  inv1  gate1199(.a(G369), .O(gate108inter8));
  nand2 gate1200(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1201(.a(s_93), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1202(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1203(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1204(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1821(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1822(.a(gate109inter0), .b(s_182), .O(gate109inter1));
  and2  gate1823(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1824(.a(s_182), .O(gate109inter3));
  inv1  gate1825(.a(s_183), .O(gate109inter4));
  nand2 gate1826(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1827(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1828(.a(G370), .O(gate109inter7));
  inv1  gate1829(.a(G371), .O(gate109inter8));
  nand2 gate1830(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1831(.a(s_183), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1832(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1833(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1834(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate631(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate632(.a(gate116inter0), .b(s_12), .O(gate116inter1));
  and2  gate633(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate634(.a(s_12), .O(gate116inter3));
  inv1  gate635(.a(s_13), .O(gate116inter4));
  nand2 gate636(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate637(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate638(.a(G384), .O(gate116inter7));
  inv1  gate639(.a(G385), .O(gate116inter8));
  nand2 gate640(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate641(.a(s_13), .b(gate116inter3), .O(gate116inter10));
  nor2  gate642(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate643(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate644(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1471(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1472(.a(gate126inter0), .b(s_132), .O(gate126inter1));
  and2  gate1473(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1474(.a(s_132), .O(gate126inter3));
  inv1  gate1475(.a(s_133), .O(gate126inter4));
  nand2 gate1476(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1477(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1478(.a(G404), .O(gate126inter7));
  inv1  gate1479(.a(G405), .O(gate126inter8));
  nand2 gate1480(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1481(.a(s_133), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1482(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1483(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1484(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1947(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1948(.a(gate134inter0), .b(s_200), .O(gate134inter1));
  and2  gate1949(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1950(.a(s_200), .O(gate134inter3));
  inv1  gate1951(.a(s_201), .O(gate134inter4));
  nand2 gate1952(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1953(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1954(.a(G420), .O(gate134inter7));
  inv1  gate1955(.a(G421), .O(gate134inter8));
  nand2 gate1956(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1957(.a(s_201), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1958(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1959(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1960(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2171(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2172(.a(gate136inter0), .b(s_232), .O(gate136inter1));
  and2  gate2173(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2174(.a(s_232), .O(gate136inter3));
  inv1  gate2175(.a(s_233), .O(gate136inter4));
  nand2 gate2176(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2177(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2178(.a(G424), .O(gate136inter7));
  inv1  gate2179(.a(G425), .O(gate136inter8));
  nand2 gate2180(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2181(.a(s_233), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2182(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2183(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2184(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1289(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1290(.a(gate141inter0), .b(s_106), .O(gate141inter1));
  and2  gate1291(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1292(.a(s_106), .O(gate141inter3));
  inv1  gate1293(.a(s_107), .O(gate141inter4));
  nand2 gate1294(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1295(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1296(.a(G450), .O(gate141inter7));
  inv1  gate1297(.a(G453), .O(gate141inter8));
  nand2 gate1298(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1299(.a(s_107), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1300(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1301(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1302(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2073(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2074(.a(gate153inter0), .b(s_218), .O(gate153inter1));
  and2  gate2075(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2076(.a(s_218), .O(gate153inter3));
  inv1  gate2077(.a(s_219), .O(gate153inter4));
  nand2 gate2078(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2079(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2080(.a(G426), .O(gate153inter7));
  inv1  gate2081(.a(G522), .O(gate153inter8));
  nand2 gate2082(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2083(.a(s_219), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2084(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2085(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2086(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate911(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate912(.a(gate154inter0), .b(s_52), .O(gate154inter1));
  and2  gate913(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate914(.a(s_52), .O(gate154inter3));
  inv1  gate915(.a(s_53), .O(gate154inter4));
  nand2 gate916(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate917(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate918(.a(G429), .O(gate154inter7));
  inv1  gate919(.a(G522), .O(gate154inter8));
  nand2 gate920(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate921(.a(s_53), .b(gate154inter3), .O(gate154inter10));
  nor2  gate922(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate923(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate924(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1079(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1080(.a(gate156inter0), .b(s_76), .O(gate156inter1));
  and2  gate1081(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1082(.a(s_76), .O(gate156inter3));
  inv1  gate1083(.a(s_77), .O(gate156inter4));
  nand2 gate1084(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1085(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1086(.a(G435), .O(gate156inter7));
  inv1  gate1087(.a(G525), .O(gate156inter8));
  nand2 gate1088(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1089(.a(s_77), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1090(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1091(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1092(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1387(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1388(.a(gate158inter0), .b(s_120), .O(gate158inter1));
  and2  gate1389(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1390(.a(s_120), .O(gate158inter3));
  inv1  gate1391(.a(s_121), .O(gate158inter4));
  nand2 gate1392(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1393(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1394(.a(G441), .O(gate158inter7));
  inv1  gate1395(.a(G528), .O(gate158inter8));
  nand2 gate1396(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1397(.a(s_121), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1398(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1399(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1400(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2325(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2326(.a(gate165inter0), .b(s_254), .O(gate165inter1));
  and2  gate2327(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2328(.a(s_254), .O(gate165inter3));
  inv1  gate2329(.a(s_255), .O(gate165inter4));
  nand2 gate2330(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2331(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2332(.a(G462), .O(gate165inter7));
  inv1  gate2333(.a(G540), .O(gate165inter8));
  nand2 gate2334(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2335(.a(s_255), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2336(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2337(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2338(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1793(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1794(.a(gate169inter0), .b(s_178), .O(gate169inter1));
  and2  gate1795(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1796(.a(s_178), .O(gate169inter3));
  inv1  gate1797(.a(s_179), .O(gate169inter4));
  nand2 gate1798(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1799(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1800(.a(G474), .O(gate169inter7));
  inv1  gate1801(.a(G546), .O(gate169inter8));
  nand2 gate1802(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1803(.a(s_179), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1804(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1805(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1806(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1051(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1052(.a(gate170inter0), .b(s_72), .O(gate170inter1));
  and2  gate1053(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1054(.a(s_72), .O(gate170inter3));
  inv1  gate1055(.a(s_73), .O(gate170inter4));
  nand2 gate1056(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1057(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1058(.a(G477), .O(gate170inter7));
  inv1  gate1059(.a(G546), .O(gate170inter8));
  nand2 gate1060(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1061(.a(s_73), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1062(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1063(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1064(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate659(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate660(.a(gate175inter0), .b(s_16), .O(gate175inter1));
  and2  gate661(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate662(.a(s_16), .O(gate175inter3));
  inv1  gate663(.a(s_17), .O(gate175inter4));
  nand2 gate664(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate665(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate666(.a(G492), .O(gate175inter7));
  inv1  gate667(.a(G555), .O(gate175inter8));
  nand2 gate668(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate669(.a(s_17), .b(gate175inter3), .O(gate175inter10));
  nor2  gate670(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate671(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate672(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate2045(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2046(.a(gate176inter0), .b(s_214), .O(gate176inter1));
  and2  gate2047(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2048(.a(s_214), .O(gate176inter3));
  inv1  gate2049(.a(s_215), .O(gate176inter4));
  nand2 gate2050(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2051(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2052(.a(G495), .O(gate176inter7));
  inv1  gate2053(.a(G555), .O(gate176inter8));
  nand2 gate2054(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2055(.a(s_215), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2056(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2057(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2058(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate1695(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1696(.a(gate177inter0), .b(s_164), .O(gate177inter1));
  and2  gate1697(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1698(.a(s_164), .O(gate177inter3));
  inv1  gate1699(.a(s_165), .O(gate177inter4));
  nand2 gate1700(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1701(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1702(.a(G498), .O(gate177inter7));
  inv1  gate1703(.a(G558), .O(gate177inter8));
  nand2 gate1704(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1705(.a(s_165), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1706(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1707(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1708(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1569(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1570(.a(gate181inter0), .b(s_146), .O(gate181inter1));
  and2  gate1571(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1572(.a(s_146), .O(gate181inter3));
  inv1  gate1573(.a(s_147), .O(gate181inter4));
  nand2 gate1574(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1575(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1576(.a(G510), .O(gate181inter7));
  inv1  gate1577(.a(G564), .O(gate181inter8));
  nand2 gate1578(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1579(.a(s_147), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1580(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1581(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1582(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2003(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2004(.a(gate182inter0), .b(s_208), .O(gate182inter1));
  and2  gate2005(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2006(.a(s_208), .O(gate182inter3));
  inv1  gate2007(.a(s_209), .O(gate182inter4));
  nand2 gate2008(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2009(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2010(.a(G513), .O(gate182inter7));
  inv1  gate2011(.a(G564), .O(gate182inter8));
  nand2 gate2012(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2013(.a(s_209), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2014(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2015(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2016(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate841(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate842(.a(gate183inter0), .b(s_42), .O(gate183inter1));
  and2  gate843(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate844(.a(s_42), .O(gate183inter3));
  inv1  gate845(.a(s_43), .O(gate183inter4));
  nand2 gate846(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate847(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate848(.a(G516), .O(gate183inter7));
  inv1  gate849(.a(G567), .O(gate183inter8));
  nand2 gate850(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate851(.a(s_43), .b(gate183inter3), .O(gate183inter10));
  nor2  gate852(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate853(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate854(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1597(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1598(.a(gate189inter0), .b(s_150), .O(gate189inter1));
  and2  gate1599(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1600(.a(s_150), .O(gate189inter3));
  inv1  gate1601(.a(s_151), .O(gate189inter4));
  nand2 gate1602(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1603(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1604(.a(G578), .O(gate189inter7));
  inv1  gate1605(.a(G579), .O(gate189inter8));
  nand2 gate1606(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1607(.a(s_151), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1608(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1609(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1610(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1373(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1374(.a(gate191inter0), .b(s_118), .O(gate191inter1));
  and2  gate1375(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1376(.a(s_118), .O(gate191inter3));
  inv1  gate1377(.a(s_119), .O(gate191inter4));
  nand2 gate1378(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1379(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1380(.a(G582), .O(gate191inter7));
  inv1  gate1381(.a(G583), .O(gate191inter8));
  nand2 gate1382(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1383(.a(s_119), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1384(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1385(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1386(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1765(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1766(.a(gate193inter0), .b(s_174), .O(gate193inter1));
  and2  gate1767(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1768(.a(s_174), .O(gate193inter3));
  inv1  gate1769(.a(s_175), .O(gate193inter4));
  nand2 gate1770(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1771(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1772(.a(G586), .O(gate193inter7));
  inv1  gate1773(.a(G587), .O(gate193inter8));
  nand2 gate1774(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1775(.a(s_175), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1776(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1777(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1778(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate813(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate814(.a(gate200inter0), .b(s_38), .O(gate200inter1));
  and2  gate815(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate816(.a(s_38), .O(gate200inter3));
  inv1  gate817(.a(s_39), .O(gate200inter4));
  nand2 gate818(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate819(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate820(.a(G600), .O(gate200inter7));
  inv1  gate821(.a(G601), .O(gate200inter8));
  nand2 gate822(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate823(.a(s_39), .b(gate200inter3), .O(gate200inter10));
  nor2  gate824(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate825(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate826(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2367(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2368(.a(gate203inter0), .b(s_260), .O(gate203inter1));
  and2  gate2369(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2370(.a(s_260), .O(gate203inter3));
  inv1  gate2371(.a(s_261), .O(gate203inter4));
  nand2 gate2372(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2373(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2374(.a(G602), .O(gate203inter7));
  inv1  gate2375(.a(G612), .O(gate203inter8));
  nand2 gate2376(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2377(.a(s_261), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2378(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2379(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2380(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1121(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1122(.a(gate206inter0), .b(s_82), .O(gate206inter1));
  and2  gate1123(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1124(.a(s_82), .O(gate206inter3));
  inv1  gate1125(.a(s_83), .O(gate206inter4));
  nand2 gate1126(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1127(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1128(.a(G632), .O(gate206inter7));
  inv1  gate1129(.a(G637), .O(gate206inter8));
  nand2 gate1130(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1131(.a(s_83), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1132(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1133(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1134(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1751(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1752(.a(gate210inter0), .b(s_172), .O(gate210inter1));
  and2  gate1753(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1754(.a(s_172), .O(gate210inter3));
  inv1  gate1755(.a(s_173), .O(gate210inter4));
  nand2 gate1756(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1757(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1758(.a(G607), .O(gate210inter7));
  inv1  gate1759(.a(G666), .O(gate210inter8));
  nand2 gate1760(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1761(.a(s_173), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1762(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1763(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1764(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1583(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1584(.a(gate216inter0), .b(s_148), .O(gate216inter1));
  and2  gate1585(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1586(.a(s_148), .O(gate216inter3));
  inv1  gate1587(.a(s_149), .O(gate216inter4));
  nand2 gate1588(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1589(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1590(.a(G617), .O(gate216inter7));
  inv1  gate1591(.a(G675), .O(gate216inter8));
  nand2 gate1592(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1593(.a(s_149), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1594(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1595(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1596(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1667(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1668(.a(gate218inter0), .b(s_160), .O(gate218inter1));
  and2  gate1669(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1670(.a(s_160), .O(gate218inter3));
  inv1  gate1671(.a(s_161), .O(gate218inter4));
  nand2 gate1672(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1673(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1674(.a(G627), .O(gate218inter7));
  inv1  gate1675(.a(G678), .O(gate218inter8));
  nand2 gate1676(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1677(.a(s_161), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1678(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1679(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1680(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1345(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1346(.a(gate221inter0), .b(s_114), .O(gate221inter1));
  and2  gate1347(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1348(.a(s_114), .O(gate221inter3));
  inv1  gate1349(.a(s_115), .O(gate221inter4));
  nand2 gate1350(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1351(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1352(.a(G622), .O(gate221inter7));
  inv1  gate1353(.a(G684), .O(gate221inter8));
  nand2 gate1354(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1355(.a(s_115), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1356(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1357(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1358(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1219(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1220(.a(gate222inter0), .b(s_96), .O(gate222inter1));
  and2  gate1221(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1222(.a(s_96), .O(gate222inter3));
  inv1  gate1223(.a(s_97), .O(gate222inter4));
  nand2 gate1224(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1225(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1226(.a(G632), .O(gate222inter7));
  inv1  gate1227(.a(G684), .O(gate222inter8));
  nand2 gate1228(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1229(.a(s_97), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1230(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1231(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1232(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1961(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1962(.a(gate225inter0), .b(s_202), .O(gate225inter1));
  and2  gate1963(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1964(.a(s_202), .O(gate225inter3));
  inv1  gate1965(.a(s_203), .O(gate225inter4));
  nand2 gate1966(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1967(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1968(.a(G690), .O(gate225inter7));
  inv1  gate1969(.a(G691), .O(gate225inter8));
  nand2 gate1970(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1971(.a(s_203), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1972(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1973(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1974(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2213(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2214(.a(gate231inter0), .b(s_238), .O(gate231inter1));
  and2  gate2215(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2216(.a(s_238), .O(gate231inter3));
  inv1  gate2217(.a(s_239), .O(gate231inter4));
  nand2 gate2218(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2219(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2220(.a(G702), .O(gate231inter7));
  inv1  gate2221(.a(G703), .O(gate231inter8));
  nand2 gate2222(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2223(.a(s_239), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2224(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2225(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2226(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate2241(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2242(.a(gate237inter0), .b(s_242), .O(gate237inter1));
  and2  gate2243(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2244(.a(s_242), .O(gate237inter3));
  inv1  gate2245(.a(s_243), .O(gate237inter4));
  nand2 gate2246(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2247(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2248(.a(G254), .O(gate237inter7));
  inv1  gate2249(.a(G706), .O(gate237inter8));
  nand2 gate2250(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2251(.a(s_243), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2252(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2253(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2254(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1331(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1332(.a(gate242inter0), .b(s_112), .O(gate242inter1));
  and2  gate1333(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1334(.a(s_112), .O(gate242inter3));
  inv1  gate1335(.a(s_113), .O(gate242inter4));
  nand2 gate1336(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1337(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1338(.a(G718), .O(gate242inter7));
  inv1  gate1339(.a(G730), .O(gate242inter8));
  nand2 gate1340(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1341(.a(s_113), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1342(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1343(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1344(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1625(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1626(.a(gate245inter0), .b(s_154), .O(gate245inter1));
  and2  gate1627(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1628(.a(s_154), .O(gate245inter3));
  inv1  gate1629(.a(s_155), .O(gate245inter4));
  nand2 gate1630(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1631(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1632(.a(G248), .O(gate245inter7));
  inv1  gate1633(.a(G736), .O(gate245inter8));
  nand2 gate1634(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1635(.a(s_155), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1636(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1637(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1638(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1009(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1010(.a(gate247inter0), .b(s_66), .O(gate247inter1));
  and2  gate1011(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1012(.a(s_66), .O(gate247inter3));
  inv1  gate1013(.a(s_67), .O(gate247inter4));
  nand2 gate1014(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1015(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1016(.a(G251), .O(gate247inter7));
  inv1  gate1017(.a(G739), .O(gate247inter8));
  nand2 gate1018(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1019(.a(s_67), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1020(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1021(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1022(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1905(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1906(.a(gate251inter0), .b(s_194), .O(gate251inter1));
  and2  gate1907(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1908(.a(s_194), .O(gate251inter3));
  inv1  gate1909(.a(s_195), .O(gate251inter4));
  nand2 gate1910(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1911(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1912(.a(G257), .O(gate251inter7));
  inv1  gate1913(.a(G745), .O(gate251inter8));
  nand2 gate1914(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1915(.a(s_195), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1916(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1917(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1918(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1107(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1108(.a(gate254inter0), .b(s_80), .O(gate254inter1));
  and2  gate1109(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1110(.a(s_80), .O(gate254inter3));
  inv1  gate1111(.a(s_81), .O(gate254inter4));
  nand2 gate1112(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1113(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1114(.a(G712), .O(gate254inter7));
  inv1  gate1115(.a(G748), .O(gate254inter8));
  nand2 gate1116(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1117(.a(s_81), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1118(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1119(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1120(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1247(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1248(.a(gate257inter0), .b(s_100), .O(gate257inter1));
  and2  gate1249(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1250(.a(s_100), .O(gate257inter3));
  inv1  gate1251(.a(s_101), .O(gate257inter4));
  nand2 gate1252(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1253(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1254(.a(G754), .O(gate257inter7));
  inv1  gate1255(.a(G755), .O(gate257inter8));
  nand2 gate1256(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1257(.a(s_101), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1258(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1259(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1260(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1779(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1780(.a(gate258inter0), .b(s_176), .O(gate258inter1));
  and2  gate1781(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1782(.a(s_176), .O(gate258inter3));
  inv1  gate1783(.a(s_177), .O(gate258inter4));
  nand2 gate1784(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1785(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1786(.a(G756), .O(gate258inter7));
  inv1  gate1787(.a(G757), .O(gate258inter8));
  nand2 gate1788(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1789(.a(s_177), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1790(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1791(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1792(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate827(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate828(.a(gate259inter0), .b(s_40), .O(gate259inter1));
  and2  gate829(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate830(.a(s_40), .O(gate259inter3));
  inv1  gate831(.a(s_41), .O(gate259inter4));
  nand2 gate832(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate833(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate834(.a(G758), .O(gate259inter7));
  inv1  gate835(.a(G759), .O(gate259inter8));
  nand2 gate836(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate837(.a(s_41), .b(gate259inter3), .O(gate259inter10));
  nor2  gate838(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate839(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate840(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate547(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate548(.a(gate268inter0), .b(s_0), .O(gate268inter1));
  and2  gate549(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate550(.a(s_0), .O(gate268inter3));
  inv1  gate551(.a(s_1), .O(gate268inter4));
  nand2 gate552(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate553(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate554(.a(G651), .O(gate268inter7));
  inv1  gate555(.a(G779), .O(gate268inter8));
  nand2 gate556(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate557(.a(s_1), .b(gate268inter3), .O(gate268inter10));
  nor2  gate558(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate559(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate560(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1835(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1836(.a(gate274inter0), .b(s_184), .O(gate274inter1));
  and2  gate1837(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1838(.a(s_184), .O(gate274inter3));
  inv1  gate1839(.a(s_185), .O(gate274inter4));
  nand2 gate1840(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1841(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1842(.a(G770), .O(gate274inter7));
  inv1  gate1843(.a(G794), .O(gate274inter8));
  nand2 gate1844(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1845(.a(s_185), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1846(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1847(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1848(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2297(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2298(.a(gate277inter0), .b(s_250), .O(gate277inter1));
  and2  gate2299(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2300(.a(s_250), .O(gate277inter3));
  inv1  gate2301(.a(s_251), .O(gate277inter4));
  nand2 gate2302(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2303(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2304(.a(G648), .O(gate277inter7));
  inv1  gate2305(.a(G800), .O(gate277inter8));
  nand2 gate2306(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2307(.a(s_251), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2308(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2309(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2310(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1723(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1724(.a(gate278inter0), .b(s_168), .O(gate278inter1));
  and2  gate1725(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1726(.a(s_168), .O(gate278inter3));
  inv1  gate1727(.a(s_169), .O(gate278inter4));
  nand2 gate1728(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1729(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1730(.a(G776), .O(gate278inter7));
  inv1  gate1731(.a(G800), .O(gate278inter8));
  nand2 gate1732(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1733(.a(s_169), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1734(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1735(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1736(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate799(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate800(.a(gate279inter0), .b(s_36), .O(gate279inter1));
  and2  gate801(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate802(.a(s_36), .O(gate279inter3));
  inv1  gate803(.a(s_37), .O(gate279inter4));
  nand2 gate804(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate805(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate806(.a(G651), .O(gate279inter7));
  inv1  gate807(.a(G803), .O(gate279inter8));
  nand2 gate808(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate809(.a(s_37), .b(gate279inter3), .O(gate279inter10));
  nor2  gate810(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate811(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate812(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate771(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate772(.a(gate280inter0), .b(s_32), .O(gate280inter1));
  and2  gate773(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate774(.a(s_32), .O(gate280inter3));
  inv1  gate775(.a(s_33), .O(gate280inter4));
  nand2 gate776(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate777(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate778(.a(G779), .O(gate280inter7));
  inv1  gate779(.a(G803), .O(gate280inter8));
  nand2 gate780(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate781(.a(s_33), .b(gate280inter3), .O(gate280inter10));
  nor2  gate782(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate783(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate784(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate757(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate758(.a(gate281inter0), .b(s_30), .O(gate281inter1));
  and2  gate759(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate760(.a(s_30), .O(gate281inter3));
  inv1  gate761(.a(s_31), .O(gate281inter4));
  nand2 gate762(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate763(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate764(.a(G654), .O(gate281inter7));
  inv1  gate765(.a(G806), .O(gate281inter8));
  nand2 gate766(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate767(.a(s_31), .b(gate281inter3), .O(gate281inter10));
  nor2  gate768(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate769(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate770(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1653(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1654(.a(gate283inter0), .b(s_158), .O(gate283inter1));
  and2  gate1655(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1656(.a(s_158), .O(gate283inter3));
  inv1  gate1657(.a(s_159), .O(gate283inter4));
  nand2 gate1658(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1659(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1660(.a(G657), .O(gate283inter7));
  inv1  gate1661(.a(G809), .O(gate283inter8));
  nand2 gate1662(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1663(.a(s_159), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1664(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1665(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1666(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate617(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate618(.a(gate284inter0), .b(s_10), .O(gate284inter1));
  and2  gate619(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate620(.a(s_10), .O(gate284inter3));
  inv1  gate621(.a(s_11), .O(gate284inter4));
  nand2 gate622(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate623(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate624(.a(G785), .O(gate284inter7));
  inv1  gate625(.a(G809), .O(gate284inter8));
  nand2 gate626(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate627(.a(s_11), .b(gate284inter3), .O(gate284inter10));
  nor2  gate628(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate629(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate630(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1863(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1864(.a(gate286inter0), .b(s_188), .O(gate286inter1));
  and2  gate1865(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1866(.a(s_188), .O(gate286inter3));
  inv1  gate1867(.a(s_189), .O(gate286inter4));
  nand2 gate1868(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1869(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1870(.a(G788), .O(gate286inter7));
  inv1  gate1871(.a(G812), .O(gate286inter8));
  nand2 gate1872(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1873(.a(s_189), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1874(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1875(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1876(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2143(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2144(.a(gate288inter0), .b(s_228), .O(gate288inter1));
  and2  gate2145(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2146(.a(s_228), .O(gate288inter3));
  inv1  gate2147(.a(s_229), .O(gate288inter4));
  nand2 gate2148(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2149(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2150(.a(G791), .O(gate288inter7));
  inv1  gate2151(.a(G815), .O(gate288inter8));
  nand2 gate2152(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2153(.a(s_229), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2154(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2155(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2156(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2157(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2158(.a(gate295inter0), .b(s_230), .O(gate295inter1));
  and2  gate2159(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2160(.a(s_230), .O(gate295inter3));
  inv1  gate2161(.a(s_231), .O(gate295inter4));
  nand2 gate2162(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2163(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2164(.a(G830), .O(gate295inter7));
  inv1  gate2165(.a(G831), .O(gate295inter8));
  nand2 gate2166(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2167(.a(s_231), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2168(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2169(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2170(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1177(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1178(.a(gate388inter0), .b(s_90), .O(gate388inter1));
  and2  gate1179(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1180(.a(s_90), .O(gate388inter3));
  inv1  gate1181(.a(s_91), .O(gate388inter4));
  nand2 gate1182(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1183(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1184(.a(G2), .O(gate388inter7));
  inv1  gate1185(.a(G1039), .O(gate388inter8));
  nand2 gate1186(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1187(.a(s_91), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1188(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1189(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1190(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1485(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1486(.a(gate393inter0), .b(s_134), .O(gate393inter1));
  and2  gate1487(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1488(.a(s_134), .O(gate393inter3));
  inv1  gate1489(.a(s_135), .O(gate393inter4));
  nand2 gate1490(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1491(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1492(.a(G7), .O(gate393inter7));
  inv1  gate1493(.a(G1054), .O(gate393inter8));
  nand2 gate1494(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1495(.a(s_135), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1496(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1497(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1498(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1359(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1360(.a(gate398inter0), .b(s_116), .O(gate398inter1));
  and2  gate1361(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1362(.a(s_116), .O(gate398inter3));
  inv1  gate1363(.a(s_117), .O(gate398inter4));
  nand2 gate1364(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1365(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1366(.a(G12), .O(gate398inter7));
  inv1  gate1367(.a(G1069), .O(gate398inter8));
  nand2 gate1368(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1369(.a(s_117), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1370(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1371(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1372(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate925(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate926(.a(gate402inter0), .b(s_54), .O(gate402inter1));
  and2  gate927(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate928(.a(s_54), .O(gate402inter3));
  inv1  gate929(.a(s_55), .O(gate402inter4));
  nand2 gate930(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate931(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate932(.a(G16), .O(gate402inter7));
  inv1  gate933(.a(G1081), .O(gate402inter8));
  nand2 gate934(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate935(.a(s_55), .b(gate402inter3), .O(gate402inter10));
  nor2  gate936(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate937(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate938(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2283(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2284(.a(gate406inter0), .b(s_248), .O(gate406inter1));
  and2  gate2285(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2286(.a(s_248), .O(gate406inter3));
  inv1  gate2287(.a(s_249), .O(gate406inter4));
  nand2 gate2288(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2289(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2290(.a(G20), .O(gate406inter7));
  inv1  gate2291(.a(G1093), .O(gate406inter8));
  nand2 gate2292(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2293(.a(s_249), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2294(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2295(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2296(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate645(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate646(.a(gate408inter0), .b(s_14), .O(gate408inter1));
  and2  gate647(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate648(.a(s_14), .O(gate408inter3));
  inv1  gate649(.a(s_15), .O(gate408inter4));
  nand2 gate650(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate651(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate652(.a(G22), .O(gate408inter7));
  inv1  gate653(.a(G1099), .O(gate408inter8));
  nand2 gate654(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate655(.a(s_15), .b(gate408inter3), .O(gate408inter10));
  nor2  gate656(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate657(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate658(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate953(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate954(.a(gate415inter0), .b(s_58), .O(gate415inter1));
  and2  gate955(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate956(.a(s_58), .O(gate415inter3));
  inv1  gate957(.a(s_59), .O(gate415inter4));
  nand2 gate958(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate959(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate960(.a(G29), .O(gate415inter7));
  inv1  gate961(.a(G1120), .O(gate415inter8));
  nand2 gate962(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate963(.a(s_59), .b(gate415inter3), .O(gate415inter10));
  nor2  gate964(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate965(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate966(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate981(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate982(.a(gate419inter0), .b(s_62), .O(gate419inter1));
  and2  gate983(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate984(.a(s_62), .O(gate419inter3));
  inv1  gate985(.a(s_63), .O(gate419inter4));
  nand2 gate986(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate987(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate988(.a(G1), .O(gate419inter7));
  inv1  gate989(.a(G1132), .O(gate419inter8));
  nand2 gate990(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate991(.a(s_63), .b(gate419inter3), .O(gate419inter10));
  nor2  gate992(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate993(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate994(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1401(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1402(.a(gate421inter0), .b(s_122), .O(gate421inter1));
  and2  gate1403(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1404(.a(s_122), .O(gate421inter3));
  inv1  gate1405(.a(s_123), .O(gate421inter4));
  nand2 gate1406(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1407(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1408(.a(G2), .O(gate421inter7));
  inv1  gate1409(.a(G1135), .O(gate421inter8));
  nand2 gate1410(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1411(.a(s_123), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1412(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1413(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1414(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate673(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate674(.a(gate423inter0), .b(s_18), .O(gate423inter1));
  and2  gate675(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate676(.a(s_18), .O(gate423inter3));
  inv1  gate677(.a(s_19), .O(gate423inter4));
  nand2 gate678(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate679(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate680(.a(G3), .O(gate423inter7));
  inv1  gate681(.a(G1138), .O(gate423inter8));
  nand2 gate682(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate683(.a(s_19), .b(gate423inter3), .O(gate423inter10));
  nor2  gate684(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate685(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate686(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2353(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2354(.a(gate424inter0), .b(s_258), .O(gate424inter1));
  and2  gate2355(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2356(.a(s_258), .O(gate424inter3));
  inv1  gate2357(.a(s_259), .O(gate424inter4));
  nand2 gate2358(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2359(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2360(.a(G1042), .O(gate424inter7));
  inv1  gate2361(.a(G1138), .O(gate424inter8));
  nand2 gate2362(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2363(.a(s_259), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2364(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2365(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2366(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2227(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2228(.a(gate432inter0), .b(s_240), .O(gate432inter1));
  and2  gate2229(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2230(.a(s_240), .O(gate432inter3));
  inv1  gate2231(.a(s_241), .O(gate432inter4));
  nand2 gate2232(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2233(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2234(.a(G1054), .O(gate432inter7));
  inv1  gate2235(.a(G1150), .O(gate432inter8));
  nand2 gate2236(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2237(.a(s_241), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2238(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2239(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2240(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1149(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1150(.a(gate434inter0), .b(s_86), .O(gate434inter1));
  and2  gate1151(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1152(.a(s_86), .O(gate434inter3));
  inv1  gate1153(.a(s_87), .O(gate434inter4));
  nand2 gate1154(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1155(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1156(.a(G1057), .O(gate434inter7));
  inv1  gate1157(.a(G1153), .O(gate434inter8));
  nand2 gate1158(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1159(.a(s_87), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1160(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1161(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1162(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1415(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1416(.a(gate435inter0), .b(s_124), .O(gate435inter1));
  and2  gate1417(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1418(.a(s_124), .O(gate435inter3));
  inv1  gate1419(.a(s_125), .O(gate435inter4));
  nand2 gate1420(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1421(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1422(.a(G9), .O(gate435inter7));
  inv1  gate1423(.a(G1156), .O(gate435inter8));
  nand2 gate1424(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1425(.a(s_125), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1426(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1427(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1428(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate785(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate786(.a(gate445inter0), .b(s_34), .O(gate445inter1));
  and2  gate787(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate788(.a(s_34), .O(gate445inter3));
  inv1  gate789(.a(s_35), .O(gate445inter4));
  nand2 gate790(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate791(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate792(.a(G14), .O(gate445inter7));
  inv1  gate793(.a(G1171), .O(gate445inter8));
  nand2 gate794(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate795(.a(s_35), .b(gate445inter3), .O(gate445inter10));
  nor2  gate796(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate797(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate798(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1205(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1206(.a(gate446inter0), .b(s_94), .O(gate446inter1));
  and2  gate1207(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1208(.a(s_94), .O(gate446inter3));
  inv1  gate1209(.a(s_95), .O(gate446inter4));
  nand2 gate1210(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1211(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1212(.a(G1075), .O(gate446inter7));
  inv1  gate1213(.a(G1171), .O(gate446inter8));
  nand2 gate1214(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1215(.a(s_95), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1216(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1217(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1218(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1317(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1318(.a(gate452inter0), .b(s_110), .O(gate452inter1));
  and2  gate1319(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1320(.a(s_110), .O(gate452inter3));
  inv1  gate1321(.a(s_111), .O(gate452inter4));
  nand2 gate1322(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1323(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1324(.a(G1084), .O(gate452inter7));
  inv1  gate1325(.a(G1180), .O(gate452inter8));
  nand2 gate1326(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1327(.a(s_111), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1328(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1329(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1330(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2087(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2088(.a(gate454inter0), .b(s_220), .O(gate454inter1));
  and2  gate2089(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2090(.a(s_220), .O(gate454inter3));
  inv1  gate2091(.a(s_221), .O(gate454inter4));
  nand2 gate2092(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2093(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2094(.a(G1087), .O(gate454inter7));
  inv1  gate2095(.a(G1183), .O(gate454inter8));
  nand2 gate2096(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2097(.a(s_221), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2098(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2099(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2100(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate729(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate730(.a(gate457inter0), .b(s_26), .O(gate457inter1));
  and2  gate731(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate732(.a(s_26), .O(gate457inter3));
  inv1  gate733(.a(s_27), .O(gate457inter4));
  nand2 gate734(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate735(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate736(.a(G20), .O(gate457inter7));
  inv1  gate737(.a(G1189), .O(gate457inter8));
  nand2 gate738(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate739(.a(s_27), .b(gate457inter3), .O(gate457inter10));
  nor2  gate740(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate741(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate742(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate897(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate898(.a(gate460inter0), .b(s_50), .O(gate460inter1));
  and2  gate899(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate900(.a(s_50), .O(gate460inter3));
  inv1  gate901(.a(s_51), .O(gate460inter4));
  nand2 gate902(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate903(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate904(.a(G1096), .O(gate460inter7));
  inv1  gate905(.a(G1192), .O(gate460inter8));
  nand2 gate906(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate907(.a(s_51), .b(gate460inter3), .O(gate460inter10));
  nor2  gate908(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate909(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate910(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate1891(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1892(.a(gate461inter0), .b(s_192), .O(gate461inter1));
  and2  gate1893(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1894(.a(s_192), .O(gate461inter3));
  inv1  gate1895(.a(s_193), .O(gate461inter4));
  nand2 gate1896(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1897(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1898(.a(G22), .O(gate461inter7));
  inv1  gate1899(.a(G1195), .O(gate461inter8));
  nand2 gate1900(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1901(.a(s_193), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1902(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1903(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1904(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1093(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1094(.a(gate464inter0), .b(s_78), .O(gate464inter1));
  and2  gate1095(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1096(.a(s_78), .O(gate464inter3));
  inv1  gate1097(.a(s_79), .O(gate464inter4));
  nand2 gate1098(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1099(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1100(.a(G1102), .O(gate464inter7));
  inv1  gate1101(.a(G1198), .O(gate464inter8));
  nand2 gate1102(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1103(.a(s_79), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1104(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1105(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1106(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2269(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2270(.a(gate465inter0), .b(s_246), .O(gate465inter1));
  and2  gate2271(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2272(.a(s_246), .O(gate465inter3));
  inv1  gate2273(.a(s_247), .O(gate465inter4));
  nand2 gate2274(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2275(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2276(.a(G24), .O(gate465inter7));
  inv1  gate2277(.a(G1201), .O(gate465inter8));
  nand2 gate2278(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2279(.a(s_247), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2280(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2281(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2282(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2031(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2032(.a(gate469inter0), .b(s_212), .O(gate469inter1));
  and2  gate2033(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2034(.a(s_212), .O(gate469inter3));
  inv1  gate2035(.a(s_213), .O(gate469inter4));
  nand2 gate2036(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2037(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2038(.a(G26), .O(gate469inter7));
  inv1  gate2039(.a(G1207), .O(gate469inter8));
  nand2 gate2040(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2041(.a(s_213), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2042(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2043(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2044(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1639(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1640(.a(gate471inter0), .b(s_156), .O(gate471inter1));
  and2  gate1641(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1642(.a(s_156), .O(gate471inter3));
  inv1  gate1643(.a(s_157), .O(gate471inter4));
  nand2 gate1644(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1645(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1646(.a(G27), .O(gate471inter7));
  inv1  gate1647(.a(G1210), .O(gate471inter8));
  nand2 gate1648(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1649(.a(s_157), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1650(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1651(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1652(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate939(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate940(.a(gate472inter0), .b(s_56), .O(gate472inter1));
  and2  gate941(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate942(.a(s_56), .O(gate472inter3));
  inv1  gate943(.a(s_57), .O(gate472inter4));
  nand2 gate944(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate945(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate946(.a(G1114), .O(gate472inter7));
  inv1  gate947(.a(G1210), .O(gate472inter8));
  nand2 gate948(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate949(.a(s_57), .b(gate472inter3), .O(gate472inter10));
  nor2  gate950(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate951(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate952(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate883(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate884(.a(gate477inter0), .b(s_48), .O(gate477inter1));
  and2  gate885(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate886(.a(s_48), .O(gate477inter3));
  inv1  gate887(.a(s_49), .O(gate477inter4));
  nand2 gate888(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate889(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate890(.a(G30), .O(gate477inter7));
  inv1  gate891(.a(G1219), .O(gate477inter8));
  nand2 gate892(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate893(.a(s_49), .b(gate477inter3), .O(gate477inter10));
  nor2  gate894(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate895(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate896(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1429(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1430(.a(gate480inter0), .b(s_126), .O(gate480inter1));
  and2  gate1431(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1432(.a(s_126), .O(gate480inter3));
  inv1  gate1433(.a(s_127), .O(gate480inter4));
  nand2 gate1434(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1435(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1436(.a(G1126), .O(gate480inter7));
  inv1  gate1437(.a(G1222), .O(gate480inter8));
  nand2 gate1438(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1439(.a(s_127), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1440(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1441(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1442(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1541(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1542(.a(gate483inter0), .b(s_142), .O(gate483inter1));
  and2  gate1543(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1544(.a(s_142), .O(gate483inter3));
  inv1  gate1545(.a(s_143), .O(gate483inter4));
  nand2 gate1546(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1547(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1548(.a(G1228), .O(gate483inter7));
  inv1  gate1549(.a(G1229), .O(gate483inter8));
  nand2 gate1550(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1551(.a(s_143), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1552(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1553(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1554(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate561(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate562(.a(gate484inter0), .b(s_2), .O(gate484inter1));
  and2  gate563(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate564(.a(s_2), .O(gate484inter3));
  inv1  gate565(.a(s_3), .O(gate484inter4));
  nand2 gate566(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate567(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate568(.a(G1230), .O(gate484inter7));
  inv1  gate569(.a(G1231), .O(gate484inter8));
  nand2 gate570(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate571(.a(s_3), .b(gate484inter3), .O(gate484inter10));
  nor2  gate572(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate573(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate574(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1975(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1976(.a(gate486inter0), .b(s_204), .O(gate486inter1));
  and2  gate1977(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1978(.a(s_204), .O(gate486inter3));
  inv1  gate1979(.a(s_205), .O(gate486inter4));
  nand2 gate1980(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1981(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1982(.a(G1234), .O(gate486inter7));
  inv1  gate1983(.a(G1235), .O(gate486inter8));
  nand2 gate1984(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1985(.a(s_205), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1986(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1987(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1988(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2101(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2102(.a(gate487inter0), .b(s_222), .O(gate487inter1));
  and2  gate2103(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2104(.a(s_222), .O(gate487inter3));
  inv1  gate2105(.a(s_223), .O(gate487inter4));
  nand2 gate2106(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2107(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2108(.a(G1236), .O(gate487inter7));
  inv1  gate2109(.a(G1237), .O(gate487inter8));
  nand2 gate2110(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2111(.a(s_223), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2112(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2113(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2114(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1499(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1500(.a(gate488inter0), .b(s_136), .O(gate488inter1));
  and2  gate1501(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1502(.a(s_136), .O(gate488inter3));
  inv1  gate1503(.a(s_137), .O(gate488inter4));
  nand2 gate1504(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1505(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1506(.a(G1238), .O(gate488inter7));
  inv1  gate1507(.a(G1239), .O(gate488inter8));
  nand2 gate1508(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1509(.a(s_137), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1510(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1511(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1512(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1555(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1556(.a(gate489inter0), .b(s_144), .O(gate489inter1));
  and2  gate1557(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1558(.a(s_144), .O(gate489inter3));
  inv1  gate1559(.a(s_145), .O(gate489inter4));
  nand2 gate1560(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1561(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1562(.a(G1240), .O(gate489inter7));
  inv1  gate1563(.a(G1241), .O(gate489inter8));
  nand2 gate1564(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1565(.a(s_145), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1566(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1567(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1568(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1709(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1710(.a(gate492inter0), .b(s_166), .O(gate492inter1));
  and2  gate1711(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1712(.a(s_166), .O(gate492inter3));
  inv1  gate1713(.a(s_167), .O(gate492inter4));
  nand2 gate1714(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1715(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1716(.a(G1246), .O(gate492inter7));
  inv1  gate1717(.a(G1247), .O(gate492inter8));
  nand2 gate1718(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1719(.a(s_167), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1720(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1721(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1722(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate2255(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2256(.a(gate502inter0), .b(s_244), .O(gate502inter1));
  and2  gate2257(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2258(.a(s_244), .O(gate502inter3));
  inv1  gate2259(.a(s_245), .O(gate502inter4));
  nand2 gate2260(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2261(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2262(.a(G1266), .O(gate502inter7));
  inv1  gate2263(.a(G1267), .O(gate502inter8));
  nand2 gate2264(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2265(.a(s_245), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2266(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2267(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2268(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1457(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1458(.a(gate508inter0), .b(s_130), .O(gate508inter1));
  and2  gate1459(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1460(.a(s_130), .O(gate508inter3));
  inv1  gate1461(.a(s_131), .O(gate508inter4));
  nand2 gate1462(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1463(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1464(.a(G1278), .O(gate508inter7));
  inv1  gate1465(.a(G1279), .O(gate508inter8));
  nand2 gate1466(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1467(.a(s_131), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1468(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1469(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1470(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1737(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1738(.a(gate513inter0), .b(s_170), .O(gate513inter1));
  and2  gate1739(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1740(.a(s_170), .O(gate513inter3));
  inv1  gate1741(.a(s_171), .O(gate513inter4));
  nand2 gate1742(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1743(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1744(.a(G1288), .O(gate513inter7));
  inv1  gate1745(.a(G1289), .O(gate513inter8));
  nand2 gate1746(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1747(.a(s_171), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1748(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1749(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1750(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1261(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1262(.a(gate514inter0), .b(s_102), .O(gate514inter1));
  and2  gate1263(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1264(.a(s_102), .O(gate514inter3));
  inv1  gate1265(.a(s_103), .O(gate514inter4));
  nand2 gate1266(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1267(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1268(.a(G1290), .O(gate514inter7));
  inv1  gate1269(.a(G1291), .O(gate514inter8));
  nand2 gate1270(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1271(.a(s_103), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1272(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1273(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1274(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule