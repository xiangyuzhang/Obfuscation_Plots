module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate743(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate744(.a(gate15inter0), .b(s_28), .O(gate15inter1));
  and2  gate745(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate746(.a(s_28), .O(gate15inter3));
  inv1  gate747(.a(s_29), .O(gate15inter4));
  nand2 gate748(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate749(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate750(.a(G13), .O(gate15inter7));
  inv1  gate751(.a(G14), .O(gate15inter8));
  nand2 gate752(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate753(.a(s_29), .b(gate15inter3), .O(gate15inter10));
  nor2  gate754(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate755(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate756(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate967(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate968(.a(gate16inter0), .b(s_60), .O(gate16inter1));
  and2  gate969(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate970(.a(s_60), .O(gate16inter3));
  inv1  gate971(.a(s_61), .O(gate16inter4));
  nand2 gate972(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate973(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate974(.a(G15), .O(gate16inter7));
  inv1  gate975(.a(G16), .O(gate16inter8));
  nand2 gate976(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate977(.a(s_61), .b(gate16inter3), .O(gate16inter10));
  nor2  gate978(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate979(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate980(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1023(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1024(.a(gate22inter0), .b(s_68), .O(gate22inter1));
  and2  gate1025(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1026(.a(s_68), .O(gate22inter3));
  inv1  gate1027(.a(s_69), .O(gate22inter4));
  nand2 gate1028(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1029(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1030(.a(G27), .O(gate22inter7));
  inv1  gate1031(.a(G28), .O(gate22inter8));
  nand2 gate1032(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1033(.a(s_69), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1034(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1035(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1036(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1261(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1262(.a(gate27inter0), .b(s_102), .O(gate27inter1));
  and2  gate1263(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1264(.a(s_102), .O(gate27inter3));
  inv1  gate1265(.a(s_103), .O(gate27inter4));
  nand2 gate1266(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1267(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1268(.a(G2), .O(gate27inter7));
  inv1  gate1269(.a(G6), .O(gate27inter8));
  nand2 gate1270(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1271(.a(s_103), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1272(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1273(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1274(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate547(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate548(.a(gate28inter0), .b(s_0), .O(gate28inter1));
  and2  gate549(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate550(.a(s_0), .O(gate28inter3));
  inv1  gate551(.a(s_1), .O(gate28inter4));
  nand2 gate552(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate553(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate554(.a(G10), .O(gate28inter7));
  inv1  gate555(.a(G14), .O(gate28inter8));
  nand2 gate556(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate557(.a(s_1), .b(gate28inter3), .O(gate28inter10));
  nor2  gate558(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate559(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate560(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1205(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1206(.a(gate31inter0), .b(s_94), .O(gate31inter1));
  and2  gate1207(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1208(.a(s_94), .O(gate31inter3));
  inv1  gate1209(.a(s_95), .O(gate31inter4));
  nand2 gate1210(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1211(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1212(.a(G4), .O(gate31inter7));
  inv1  gate1213(.a(G8), .O(gate31inter8));
  nand2 gate1214(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1215(.a(s_95), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1216(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1217(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1218(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate981(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate982(.a(gate35inter0), .b(s_62), .O(gate35inter1));
  and2  gate983(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate984(.a(s_62), .O(gate35inter3));
  inv1  gate985(.a(s_63), .O(gate35inter4));
  nand2 gate986(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate987(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate988(.a(G18), .O(gate35inter7));
  inv1  gate989(.a(G22), .O(gate35inter8));
  nand2 gate990(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate991(.a(s_63), .b(gate35inter3), .O(gate35inter10));
  nor2  gate992(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate993(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate994(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate617(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate618(.a(gate37inter0), .b(s_10), .O(gate37inter1));
  and2  gate619(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate620(.a(s_10), .O(gate37inter3));
  inv1  gate621(.a(s_11), .O(gate37inter4));
  nand2 gate622(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate623(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate624(.a(G19), .O(gate37inter7));
  inv1  gate625(.a(G23), .O(gate37inter8));
  nand2 gate626(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate627(.a(s_11), .b(gate37inter3), .O(gate37inter10));
  nor2  gate628(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate629(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate630(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1345(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1346(.a(gate40inter0), .b(s_114), .O(gate40inter1));
  and2  gate1347(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1348(.a(s_114), .O(gate40inter3));
  inv1  gate1349(.a(s_115), .O(gate40inter4));
  nand2 gate1350(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1351(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1352(.a(G28), .O(gate40inter7));
  inv1  gate1353(.a(G32), .O(gate40inter8));
  nand2 gate1354(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1355(.a(s_115), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1356(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1357(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1358(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1191(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1192(.a(gate41inter0), .b(s_92), .O(gate41inter1));
  and2  gate1193(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1194(.a(s_92), .O(gate41inter3));
  inv1  gate1195(.a(s_93), .O(gate41inter4));
  nand2 gate1196(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1197(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1198(.a(G1), .O(gate41inter7));
  inv1  gate1199(.a(G266), .O(gate41inter8));
  nand2 gate1200(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1201(.a(s_93), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1202(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1203(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1204(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate897(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate898(.a(gate42inter0), .b(s_50), .O(gate42inter1));
  and2  gate899(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate900(.a(s_50), .O(gate42inter3));
  inv1  gate901(.a(s_51), .O(gate42inter4));
  nand2 gate902(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate903(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate904(.a(G2), .O(gate42inter7));
  inv1  gate905(.a(G266), .O(gate42inter8));
  nand2 gate906(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate907(.a(s_51), .b(gate42inter3), .O(gate42inter10));
  nor2  gate908(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate909(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate910(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1065(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1066(.a(gate50inter0), .b(s_74), .O(gate50inter1));
  and2  gate1067(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1068(.a(s_74), .O(gate50inter3));
  inv1  gate1069(.a(s_75), .O(gate50inter4));
  nand2 gate1070(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1071(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1072(.a(G10), .O(gate50inter7));
  inv1  gate1073(.a(G278), .O(gate50inter8));
  nand2 gate1074(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1075(.a(s_75), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1076(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1077(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1078(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate771(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate772(.a(gate67inter0), .b(s_32), .O(gate67inter1));
  and2  gate773(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate774(.a(s_32), .O(gate67inter3));
  inv1  gate775(.a(s_33), .O(gate67inter4));
  nand2 gate776(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate777(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate778(.a(G27), .O(gate67inter7));
  inv1  gate779(.a(G305), .O(gate67inter8));
  nand2 gate780(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate781(.a(s_33), .b(gate67inter3), .O(gate67inter10));
  nor2  gate782(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate783(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate784(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1009(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1010(.a(gate69inter0), .b(s_66), .O(gate69inter1));
  and2  gate1011(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1012(.a(s_66), .O(gate69inter3));
  inv1  gate1013(.a(s_67), .O(gate69inter4));
  nand2 gate1014(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1015(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1016(.a(G29), .O(gate69inter7));
  inv1  gate1017(.a(G308), .O(gate69inter8));
  nand2 gate1018(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1019(.a(s_67), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1020(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1021(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1022(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1163(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1164(.a(gate77inter0), .b(s_88), .O(gate77inter1));
  and2  gate1165(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1166(.a(s_88), .O(gate77inter3));
  inv1  gate1167(.a(s_89), .O(gate77inter4));
  nand2 gate1168(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1169(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1170(.a(G2), .O(gate77inter7));
  inv1  gate1171(.a(G320), .O(gate77inter8));
  nand2 gate1172(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1173(.a(s_89), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1174(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1175(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1176(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1429(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1430(.a(gate81inter0), .b(s_126), .O(gate81inter1));
  and2  gate1431(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1432(.a(s_126), .O(gate81inter3));
  inv1  gate1433(.a(s_127), .O(gate81inter4));
  nand2 gate1434(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1435(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1436(.a(G3), .O(gate81inter7));
  inv1  gate1437(.a(G326), .O(gate81inter8));
  nand2 gate1438(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1439(.a(s_127), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1440(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1441(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1442(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate575(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate576(.a(gate88inter0), .b(s_4), .O(gate88inter1));
  and2  gate577(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate578(.a(s_4), .O(gate88inter3));
  inv1  gate579(.a(s_5), .O(gate88inter4));
  nand2 gate580(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate581(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate582(.a(G16), .O(gate88inter7));
  inv1  gate583(.a(G335), .O(gate88inter8));
  nand2 gate584(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate585(.a(s_5), .b(gate88inter3), .O(gate88inter10));
  nor2  gate586(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate587(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate588(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1107(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1108(.a(gate105inter0), .b(s_80), .O(gate105inter1));
  and2  gate1109(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1110(.a(s_80), .O(gate105inter3));
  inv1  gate1111(.a(s_81), .O(gate105inter4));
  nand2 gate1112(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1113(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1114(.a(G362), .O(gate105inter7));
  inv1  gate1115(.a(G363), .O(gate105inter8));
  nand2 gate1116(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1117(.a(s_81), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1118(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1119(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1120(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate995(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate996(.a(gate109inter0), .b(s_64), .O(gate109inter1));
  and2  gate997(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate998(.a(s_64), .O(gate109inter3));
  inv1  gate999(.a(s_65), .O(gate109inter4));
  nand2 gate1000(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1001(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1002(.a(G370), .O(gate109inter7));
  inv1  gate1003(.a(G371), .O(gate109inter8));
  nand2 gate1004(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1005(.a(s_65), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1006(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1007(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1008(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate757(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate758(.a(gate110inter0), .b(s_30), .O(gate110inter1));
  and2  gate759(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate760(.a(s_30), .O(gate110inter3));
  inv1  gate761(.a(s_31), .O(gate110inter4));
  nand2 gate762(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate763(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate764(.a(G372), .O(gate110inter7));
  inv1  gate765(.a(G373), .O(gate110inter8));
  nand2 gate766(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate767(.a(s_31), .b(gate110inter3), .O(gate110inter10));
  nor2  gate768(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate769(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate770(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1275(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1276(.a(gate117inter0), .b(s_104), .O(gate117inter1));
  and2  gate1277(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1278(.a(s_104), .O(gate117inter3));
  inv1  gate1279(.a(s_105), .O(gate117inter4));
  nand2 gate1280(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1281(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1282(.a(G386), .O(gate117inter7));
  inv1  gate1283(.a(G387), .O(gate117inter8));
  nand2 gate1284(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1285(.a(s_105), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1286(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1287(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1288(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate1093(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1094(.a(gate118inter0), .b(s_78), .O(gate118inter1));
  and2  gate1095(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1096(.a(s_78), .O(gate118inter3));
  inv1  gate1097(.a(s_79), .O(gate118inter4));
  nand2 gate1098(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1099(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1100(.a(G388), .O(gate118inter7));
  inv1  gate1101(.a(G389), .O(gate118inter8));
  nand2 gate1102(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1103(.a(s_79), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1104(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1105(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1106(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1079(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1080(.a(gate121inter0), .b(s_76), .O(gate121inter1));
  and2  gate1081(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1082(.a(s_76), .O(gate121inter3));
  inv1  gate1083(.a(s_77), .O(gate121inter4));
  nand2 gate1084(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1085(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1086(.a(G394), .O(gate121inter7));
  inv1  gate1087(.a(G395), .O(gate121inter8));
  nand2 gate1088(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1089(.a(s_77), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1090(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1091(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1092(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1121(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1122(.a(gate141inter0), .b(s_82), .O(gate141inter1));
  and2  gate1123(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1124(.a(s_82), .O(gate141inter3));
  inv1  gate1125(.a(s_83), .O(gate141inter4));
  nand2 gate1126(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1127(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1128(.a(G450), .O(gate141inter7));
  inv1  gate1129(.a(G453), .O(gate141inter8));
  nand2 gate1130(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1131(.a(s_83), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1132(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1133(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1134(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1219(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1220(.a(gate150inter0), .b(s_96), .O(gate150inter1));
  and2  gate1221(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1222(.a(s_96), .O(gate150inter3));
  inv1  gate1223(.a(s_97), .O(gate150inter4));
  nand2 gate1224(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1225(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1226(.a(G504), .O(gate150inter7));
  inv1  gate1227(.a(G507), .O(gate150inter8));
  nand2 gate1228(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1229(.a(s_97), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1230(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1231(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1232(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate799(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate800(.a(gate151inter0), .b(s_36), .O(gate151inter1));
  and2  gate801(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate802(.a(s_36), .O(gate151inter3));
  inv1  gate803(.a(s_37), .O(gate151inter4));
  nand2 gate804(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate805(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate806(.a(G510), .O(gate151inter7));
  inv1  gate807(.a(G513), .O(gate151inter8));
  nand2 gate808(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate809(.a(s_37), .b(gate151inter3), .O(gate151inter10));
  nor2  gate810(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate811(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate812(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate855(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate856(.a(gate159inter0), .b(s_44), .O(gate159inter1));
  and2  gate857(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate858(.a(s_44), .O(gate159inter3));
  inv1  gate859(.a(s_45), .O(gate159inter4));
  nand2 gate860(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate861(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate862(.a(G444), .O(gate159inter7));
  inv1  gate863(.a(G531), .O(gate159inter8));
  nand2 gate864(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate865(.a(s_45), .b(gate159inter3), .O(gate159inter10));
  nor2  gate866(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate867(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate868(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1373(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1374(.a(gate163inter0), .b(s_118), .O(gate163inter1));
  and2  gate1375(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1376(.a(s_118), .O(gate163inter3));
  inv1  gate1377(.a(s_119), .O(gate163inter4));
  nand2 gate1378(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1379(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1380(.a(G456), .O(gate163inter7));
  inv1  gate1381(.a(G537), .O(gate163inter8));
  nand2 gate1382(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1383(.a(s_119), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1384(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1385(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1386(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate659(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate660(.a(gate166inter0), .b(s_16), .O(gate166inter1));
  and2  gate661(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate662(.a(s_16), .O(gate166inter3));
  inv1  gate663(.a(s_17), .O(gate166inter4));
  nand2 gate664(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate665(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate666(.a(G465), .O(gate166inter7));
  inv1  gate667(.a(G540), .O(gate166inter8));
  nand2 gate668(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate669(.a(s_17), .b(gate166inter3), .O(gate166inter10));
  nor2  gate670(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate671(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate672(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate953(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate954(.a(gate176inter0), .b(s_58), .O(gate176inter1));
  and2  gate955(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate956(.a(s_58), .O(gate176inter3));
  inv1  gate957(.a(s_59), .O(gate176inter4));
  nand2 gate958(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate959(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate960(.a(G495), .O(gate176inter7));
  inv1  gate961(.a(G555), .O(gate176inter8));
  nand2 gate962(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate963(.a(s_59), .b(gate176inter3), .O(gate176inter10));
  nor2  gate964(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate965(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate966(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate925(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate926(.a(gate177inter0), .b(s_54), .O(gate177inter1));
  and2  gate927(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate928(.a(s_54), .O(gate177inter3));
  inv1  gate929(.a(s_55), .O(gate177inter4));
  nand2 gate930(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate931(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate932(.a(G498), .O(gate177inter7));
  inv1  gate933(.a(G558), .O(gate177inter8));
  nand2 gate934(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate935(.a(s_55), .b(gate177inter3), .O(gate177inter10));
  nor2  gate936(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate937(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate938(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1177(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1178(.a(gate178inter0), .b(s_90), .O(gate178inter1));
  and2  gate1179(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1180(.a(s_90), .O(gate178inter3));
  inv1  gate1181(.a(s_91), .O(gate178inter4));
  nand2 gate1182(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1183(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1184(.a(G501), .O(gate178inter7));
  inv1  gate1185(.a(G558), .O(gate178inter8));
  nand2 gate1186(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1187(.a(s_91), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1188(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1189(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1190(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate701(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate702(.a(gate195inter0), .b(s_22), .O(gate195inter1));
  and2  gate703(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate704(.a(s_22), .O(gate195inter3));
  inv1  gate705(.a(s_23), .O(gate195inter4));
  nand2 gate706(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate707(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate708(.a(G590), .O(gate195inter7));
  inv1  gate709(.a(G591), .O(gate195inter8));
  nand2 gate710(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate711(.a(s_23), .b(gate195inter3), .O(gate195inter10));
  nor2  gate712(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate713(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate714(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1317(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1318(.a(gate207inter0), .b(s_110), .O(gate207inter1));
  and2  gate1319(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1320(.a(s_110), .O(gate207inter3));
  inv1  gate1321(.a(s_111), .O(gate207inter4));
  nand2 gate1322(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1323(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1324(.a(G622), .O(gate207inter7));
  inv1  gate1325(.a(G632), .O(gate207inter8));
  nand2 gate1326(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1327(.a(s_111), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1328(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1329(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1330(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1387(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1388(.a(gate210inter0), .b(s_120), .O(gate210inter1));
  and2  gate1389(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1390(.a(s_120), .O(gate210inter3));
  inv1  gate1391(.a(s_121), .O(gate210inter4));
  nand2 gate1392(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1393(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1394(.a(G607), .O(gate210inter7));
  inv1  gate1395(.a(G666), .O(gate210inter8));
  nand2 gate1396(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1397(.a(s_121), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1398(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1399(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1400(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1135(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1136(.a(gate213inter0), .b(s_84), .O(gate213inter1));
  and2  gate1137(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1138(.a(s_84), .O(gate213inter3));
  inv1  gate1139(.a(s_85), .O(gate213inter4));
  nand2 gate1140(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1141(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1142(.a(G602), .O(gate213inter7));
  inv1  gate1143(.a(G672), .O(gate213inter8));
  nand2 gate1144(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1145(.a(s_85), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1146(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1147(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1148(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate883(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate884(.a(gate217inter0), .b(s_48), .O(gate217inter1));
  and2  gate885(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate886(.a(s_48), .O(gate217inter3));
  inv1  gate887(.a(s_49), .O(gate217inter4));
  nand2 gate888(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate889(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate890(.a(G622), .O(gate217inter7));
  inv1  gate891(.a(G678), .O(gate217inter8));
  nand2 gate892(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate893(.a(s_49), .b(gate217inter3), .O(gate217inter10));
  nor2  gate894(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate895(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate896(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate589(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate590(.a(gate226inter0), .b(s_6), .O(gate226inter1));
  and2  gate591(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate592(.a(s_6), .O(gate226inter3));
  inv1  gate593(.a(s_7), .O(gate226inter4));
  nand2 gate594(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate595(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate596(.a(G692), .O(gate226inter7));
  inv1  gate597(.a(G693), .O(gate226inter8));
  nand2 gate598(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate599(.a(s_7), .b(gate226inter3), .O(gate226inter10));
  nor2  gate600(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate601(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate602(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1051(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1052(.a(gate233inter0), .b(s_72), .O(gate233inter1));
  and2  gate1053(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1054(.a(s_72), .O(gate233inter3));
  inv1  gate1055(.a(s_73), .O(gate233inter4));
  nand2 gate1056(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1057(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1058(.a(G242), .O(gate233inter7));
  inv1  gate1059(.a(G718), .O(gate233inter8));
  nand2 gate1060(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1061(.a(s_73), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1062(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1063(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1064(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate673(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate674(.a(gate240inter0), .b(s_18), .O(gate240inter1));
  and2  gate675(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate676(.a(s_18), .O(gate240inter3));
  inv1  gate677(.a(s_19), .O(gate240inter4));
  nand2 gate678(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate679(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate680(.a(G263), .O(gate240inter7));
  inv1  gate681(.a(G715), .O(gate240inter8));
  nand2 gate682(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate683(.a(s_19), .b(gate240inter3), .O(gate240inter10));
  nor2  gate684(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate685(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate686(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1303(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1304(.a(gate242inter0), .b(s_108), .O(gate242inter1));
  and2  gate1305(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1306(.a(s_108), .O(gate242inter3));
  inv1  gate1307(.a(s_109), .O(gate242inter4));
  nand2 gate1308(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1309(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1310(.a(G718), .O(gate242inter7));
  inv1  gate1311(.a(G730), .O(gate242inter8));
  nand2 gate1312(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1313(.a(s_109), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1314(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1315(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1316(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate841(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate842(.a(gate250inter0), .b(s_42), .O(gate250inter1));
  and2  gate843(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate844(.a(s_42), .O(gate250inter3));
  inv1  gate845(.a(s_43), .O(gate250inter4));
  nand2 gate846(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate847(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate848(.a(G706), .O(gate250inter7));
  inv1  gate849(.a(G742), .O(gate250inter8));
  nand2 gate850(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate851(.a(s_43), .b(gate250inter3), .O(gate250inter10));
  nor2  gate852(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate853(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate854(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate645(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate646(.a(gate255inter0), .b(s_14), .O(gate255inter1));
  and2  gate647(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate648(.a(s_14), .O(gate255inter3));
  inv1  gate649(.a(s_15), .O(gate255inter4));
  nand2 gate650(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate651(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate652(.a(G263), .O(gate255inter7));
  inv1  gate653(.a(G751), .O(gate255inter8));
  nand2 gate654(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate655(.a(s_15), .b(gate255inter3), .O(gate255inter10));
  nor2  gate656(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate657(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate658(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1457(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1458(.a(gate256inter0), .b(s_130), .O(gate256inter1));
  and2  gate1459(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1460(.a(s_130), .O(gate256inter3));
  inv1  gate1461(.a(s_131), .O(gate256inter4));
  nand2 gate1462(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1463(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1464(.a(G715), .O(gate256inter7));
  inv1  gate1465(.a(G751), .O(gate256inter8));
  nand2 gate1466(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1467(.a(s_131), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1468(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1469(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1470(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate687(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate688(.a(gate267inter0), .b(s_20), .O(gate267inter1));
  and2  gate689(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate690(.a(s_20), .O(gate267inter3));
  inv1  gate691(.a(s_21), .O(gate267inter4));
  nand2 gate692(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate693(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate694(.a(G648), .O(gate267inter7));
  inv1  gate695(.a(G776), .O(gate267inter8));
  nand2 gate696(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate697(.a(s_21), .b(gate267inter3), .O(gate267inter10));
  nor2  gate698(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate699(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate700(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1401(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1402(.a(gate268inter0), .b(s_122), .O(gate268inter1));
  and2  gate1403(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1404(.a(s_122), .O(gate268inter3));
  inv1  gate1405(.a(s_123), .O(gate268inter4));
  nand2 gate1406(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1407(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1408(.a(G651), .O(gate268inter7));
  inv1  gate1409(.a(G779), .O(gate268inter8));
  nand2 gate1410(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1411(.a(s_123), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1412(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1413(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1414(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1247(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1248(.a(gate269inter0), .b(s_100), .O(gate269inter1));
  and2  gate1249(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1250(.a(s_100), .O(gate269inter3));
  inv1  gate1251(.a(s_101), .O(gate269inter4));
  nand2 gate1252(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1253(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1254(.a(G654), .O(gate269inter7));
  inv1  gate1255(.a(G782), .O(gate269inter8));
  nand2 gate1256(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1257(.a(s_101), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1258(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1259(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1260(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate939(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate940(.a(gate277inter0), .b(s_56), .O(gate277inter1));
  and2  gate941(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate942(.a(s_56), .O(gate277inter3));
  inv1  gate943(.a(s_57), .O(gate277inter4));
  nand2 gate944(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate945(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate946(.a(G648), .O(gate277inter7));
  inv1  gate947(.a(G800), .O(gate277inter8));
  nand2 gate948(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate949(.a(s_57), .b(gate277inter3), .O(gate277inter10));
  nor2  gate950(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate951(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate952(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1359(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1360(.a(gate288inter0), .b(s_116), .O(gate288inter1));
  and2  gate1361(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1362(.a(s_116), .O(gate288inter3));
  inv1  gate1363(.a(s_117), .O(gate288inter4));
  nand2 gate1364(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1365(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1366(.a(G791), .O(gate288inter7));
  inv1  gate1367(.a(G815), .O(gate288inter8));
  nand2 gate1368(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1369(.a(s_117), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1370(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1371(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1372(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1233(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1234(.a(gate293inter0), .b(s_98), .O(gate293inter1));
  and2  gate1235(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1236(.a(s_98), .O(gate293inter3));
  inv1  gate1237(.a(s_99), .O(gate293inter4));
  nand2 gate1238(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1239(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1240(.a(G828), .O(gate293inter7));
  inv1  gate1241(.a(G829), .O(gate293inter8));
  nand2 gate1242(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1243(.a(s_99), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1244(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1245(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1246(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate561(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate562(.a(gate397inter0), .b(s_2), .O(gate397inter1));
  and2  gate563(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate564(.a(s_2), .O(gate397inter3));
  inv1  gate565(.a(s_3), .O(gate397inter4));
  nand2 gate566(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate567(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate568(.a(G11), .O(gate397inter7));
  inv1  gate569(.a(G1066), .O(gate397inter8));
  nand2 gate570(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate571(.a(s_3), .b(gate397inter3), .O(gate397inter10));
  nor2  gate572(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate573(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate574(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate715(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate716(.a(gate398inter0), .b(s_24), .O(gate398inter1));
  and2  gate717(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate718(.a(s_24), .O(gate398inter3));
  inv1  gate719(.a(s_25), .O(gate398inter4));
  nand2 gate720(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate721(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate722(.a(G12), .O(gate398inter7));
  inv1  gate723(.a(G1069), .O(gate398inter8));
  nand2 gate724(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate725(.a(s_25), .b(gate398inter3), .O(gate398inter10));
  nor2  gate726(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate727(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate728(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1037(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1038(.a(gate406inter0), .b(s_70), .O(gate406inter1));
  and2  gate1039(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1040(.a(s_70), .O(gate406inter3));
  inv1  gate1041(.a(s_71), .O(gate406inter4));
  nand2 gate1042(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1043(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1044(.a(G20), .O(gate406inter7));
  inv1  gate1045(.a(G1093), .O(gate406inter8));
  nand2 gate1046(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1047(.a(s_71), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1048(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1049(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1050(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate729(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate730(.a(gate407inter0), .b(s_26), .O(gate407inter1));
  and2  gate731(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate732(.a(s_26), .O(gate407inter3));
  inv1  gate733(.a(s_27), .O(gate407inter4));
  nand2 gate734(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate735(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate736(.a(G21), .O(gate407inter7));
  inv1  gate737(.a(G1096), .O(gate407inter8));
  nand2 gate738(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate739(.a(s_27), .b(gate407inter3), .O(gate407inter10));
  nor2  gate740(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate741(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate742(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1415(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1416(.a(gate416inter0), .b(s_124), .O(gate416inter1));
  and2  gate1417(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1418(.a(s_124), .O(gate416inter3));
  inv1  gate1419(.a(s_125), .O(gate416inter4));
  nand2 gate1420(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1421(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1422(.a(G30), .O(gate416inter7));
  inv1  gate1423(.a(G1123), .O(gate416inter8));
  nand2 gate1424(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1425(.a(s_125), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1426(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1427(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1428(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1149(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1150(.a(gate435inter0), .b(s_86), .O(gate435inter1));
  and2  gate1151(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1152(.a(s_86), .O(gate435inter3));
  inv1  gate1153(.a(s_87), .O(gate435inter4));
  nand2 gate1154(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1155(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1156(.a(G9), .O(gate435inter7));
  inv1  gate1157(.a(G1156), .O(gate435inter8));
  nand2 gate1158(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1159(.a(s_87), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1160(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1161(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1162(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate603(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate604(.a(gate444inter0), .b(s_8), .O(gate444inter1));
  and2  gate605(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate606(.a(s_8), .O(gate444inter3));
  inv1  gate607(.a(s_9), .O(gate444inter4));
  nand2 gate608(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate609(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate610(.a(G1072), .O(gate444inter7));
  inv1  gate611(.a(G1168), .O(gate444inter8));
  nand2 gate612(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate613(.a(s_9), .b(gate444inter3), .O(gate444inter10));
  nor2  gate614(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate615(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate616(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1443(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1444(.a(gate445inter0), .b(s_128), .O(gate445inter1));
  and2  gate1445(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1446(.a(s_128), .O(gate445inter3));
  inv1  gate1447(.a(s_129), .O(gate445inter4));
  nand2 gate1448(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1449(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1450(.a(G14), .O(gate445inter7));
  inv1  gate1451(.a(G1171), .O(gate445inter8));
  nand2 gate1452(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1453(.a(s_129), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1454(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1455(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1456(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1331(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1332(.a(gate455inter0), .b(s_112), .O(gate455inter1));
  and2  gate1333(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1334(.a(s_112), .O(gate455inter3));
  inv1  gate1335(.a(s_113), .O(gate455inter4));
  nand2 gate1336(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1337(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1338(.a(G19), .O(gate455inter7));
  inv1  gate1339(.a(G1186), .O(gate455inter8));
  nand2 gate1340(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1341(.a(s_113), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1342(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1343(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1344(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate785(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate786(.a(gate467inter0), .b(s_34), .O(gate467inter1));
  and2  gate787(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate788(.a(s_34), .O(gate467inter3));
  inv1  gate789(.a(s_35), .O(gate467inter4));
  nand2 gate790(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate791(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate792(.a(G25), .O(gate467inter7));
  inv1  gate793(.a(G1204), .O(gate467inter8));
  nand2 gate794(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate795(.a(s_35), .b(gate467inter3), .O(gate467inter10));
  nor2  gate796(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate797(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate798(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate813(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate814(.a(gate470inter0), .b(s_38), .O(gate470inter1));
  and2  gate815(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate816(.a(s_38), .O(gate470inter3));
  inv1  gate817(.a(s_39), .O(gate470inter4));
  nand2 gate818(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate819(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate820(.a(G1111), .O(gate470inter7));
  inv1  gate821(.a(G1207), .O(gate470inter8));
  nand2 gate822(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate823(.a(s_39), .b(gate470inter3), .O(gate470inter10));
  nor2  gate824(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate825(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate826(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate631(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate632(.a(gate471inter0), .b(s_12), .O(gate471inter1));
  and2  gate633(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate634(.a(s_12), .O(gate471inter3));
  inv1  gate635(.a(s_13), .O(gate471inter4));
  nand2 gate636(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate637(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate638(.a(G27), .O(gate471inter7));
  inv1  gate639(.a(G1210), .O(gate471inter8));
  nand2 gate640(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate641(.a(s_13), .b(gate471inter3), .O(gate471inter10));
  nor2  gate642(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate643(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate644(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate869(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate870(.a(gate472inter0), .b(s_46), .O(gate472inter1));
  and2  gate871(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate872(.a(s_46), .O(gate472inter3));
  inv1  gate873(.a(s_47), .O(gate472inter4));
  nand2 gate874(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate875(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate876(.a(G1114), .O(gate472inter7));
  inv1  gate877(.a(G1210), .O(gate472inter8));
  nand2 gate878(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate879(.a(s_47), .b(gate472inter3), .O(gate472inter10));
  nor2  gate880(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate881(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate882(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1289(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1290(.a(gate473inter0), .b(s_106), .O(gate473inter1));
  and2  gate1291(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1292(.a(s_106), .O(gate473inter3));
  inv1  gate1293(.a(s_107), .O(gate473inter4));
  nand2 gate1294(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1295(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1296(.a(G28), .O(gate473inter7));
  inv1  gate1297(.a(G1213), .O(gate473inter8));
  nand2 gate1298(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1299(.a(s_107), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1300(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1301(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1302(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate911(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate912(.a(gate497inter0), .b(s_52), .O(gate497inter1));
  and2  gate913(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate914(.a(s_52), .O(gate497inter3));
  inv1  gate915(.a(s_53), .O(gate497inter4));
  nand2 gate916(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate917(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate918(.a(G1256), .O(gate497inter7));
  inv1  gate919(.a(G1257), .O(gate497inter8));
  nand2 gate920(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate921(.a(s_53), .b(gate497inter3), .O(gate497inter10));
  nor2  gate922(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate923(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate924(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate827(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate828(.a(gate502inter0), .b(s_40), .O(gate502inter1));
  and2  gate829(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate830(.a(s_40), .O(gate502inter3));
  inv1  gate831(.a(s_41), .O(gate502inter4));
  nand2 gate832(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate833(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate834(.a(G1266), .O(gate502inter7));
  inv1  gate835(.a(G1267), .O(gate502inter8));
  nand2 gate836(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate837(.a(s_41), .b(gate502inter3), .O(gate502inter10));
  nor2  gate838(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate839(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate840(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule