module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate827(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate828(.a(gate9inter0), .b(s_40), .O(gate9inter1));
  and2  gate829(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate830(.a(s_40), .O(gate9inter3));
  inv1  gate831(.a(s_41), .O(gate9inter4));
  nand2 gate832(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate833(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate834(.a(G1), .O(gate9inter7));
  inv1  gate835(.a(G2), .O(gate9inter8));
  nand2 gate836(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate837(.a(s_41), .b(gate9inter3), .O(gate9inter10));
  nor2  gate838(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate839(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate840(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate939(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate940(.a(gate10inter0), .b(s_56), .O(gate10inter1));
  and2  gate941(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate942(.a(s_56), .O(gate10inter3));
  inv1  gate943(.a(s_57), .O(gate10inter4));
  nand2 gate944(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate945(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate946(.a(G3), .O(gate10inter7));
  inv1  gate947(.a(G4), .O(gate10inter8));
  nand2 gate948(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate949(.a(s_57), .b(gate10inter3), .O(gate10inter10));
  nor2  gate950(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate951(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate952(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1009(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1010(.a(gate12inter0), .b(s_66), .O(gate12inter1));
  and2  gate1011(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1012(.a(s_66), .O(gate12inter3));
  inv1  gate1013(.a(s_67), .O(gate12inter4));
  nand2 gate1014(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1015(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1016(.a(G7), .O(gate12inter7));
  inv1  gate1017(.a(G8), .O(gate12inter8));
  nand2 gate1018(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1019(.a(s_67), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1020(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1021(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1022(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate981(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate982(.a(gate17inter0), .b(s_62), .O(gate17inter1));
  and2  gate983(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate984(.a(s_62), .O(gate17inter3));
  inv1  gate985(.a(s_63), .O(gate17inter4));
  nand2 gate986(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate987(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate988(.a(G17), .O(gate17inter7));
  inv1  gate989(.a(G18), .O(gate17inter8));
  nand2 gate990(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate991(.a(s_63), .b(gate17inter3), .O(gate17inter10));
  nor2  gate992(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate993(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate994(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1135(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1136(.a(gate18inter0), .b(s_84), .O(gate18inter1));
  and2  gate1137(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1138(.a(s_84), .O(gate18inter3));
  inv1  gate1139(.a(s_85), .O(gate18inter4));
  nand2 gate1140(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1141(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1142(.a(G19), .O(gate18inter7));
  inv1  gate1143(.a(G20), .O(gate18inter8));
  nand2 gate1144(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1145(.a(s_85), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1146(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1147(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1148(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate841(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate842(.a(gate24inter0), .b(s_42), .O(gate24inter1));
  and2  gate843(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate844(.a(s_42), .O(gate24inter3));
  inv1  gate845(.a(s_43), .O(gate24inter4));
  nand2 gate846(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate847(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate848(.a(G31), .O(gate24inter7));
  inv1  gate849(.a(G32), .O(gate24inter8));
  nand2 gate850(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate851(.a(s_43), .b(gate24inter3), .O(gate24inter10));
  nor2  gate852(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate853(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate854(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate673(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate674(.a(gate26inter0), .b(s_18), .O(gate26inter1));
  and2  gate675(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate676(.a(s_18), .O(gate26inter3));
  inv1  gate677(.a(s_19), .O(gate26inter4));
  nand2 gate678(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate679(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate680(.a(G9), .O(gate26inter7));
  inv1  gate681(.a(G13), .O(gate26inter8));
  nand2 gate682(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate683(.a(s_19), .b(gate26inter3), .O(gate26inter10));
  nor2  gate684(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate685(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate686(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate1205(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1206(.a(gate27inter0), .b(s_94), .O(gate27inter1));
  and2  gate1207(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1208(.a(s_94), .O(gate27inter3));
  inv1  gate1209(.a(s_95), .O(gate27inter4));
  nand2 gate1210(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1211(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1212(.a(G2), .O(gate27inter7));
  inv1  gate1213(.a(G6), .O(gate27inter8));
  nand2 gate1214(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1215(.a(s_95), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1216(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1217(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1218(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate589(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate590(.a(gate28inter0), .b(s_6), .O(gate28inter1));
  and2  gate591(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate592(.a(s_6), .O(gate28inter3));
  inv1  gate593(.a(s_7), .O(gate28inter4));
  nand2 gate594(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate595(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate596(.a(G10), .O(gate28inter7));
  inv1  gate597(.a(G14), .O(gate28inter8));
  nand2 gate598(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate599(.a(s_7), .b(gate28inter3), .O(gate28inter10));
  nor2  gate600(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate601(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate602(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1261(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1262(.a(gate33inter0), .b(s_102), .O(gate33inter1));
  and2  gate1263(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1264(.a(s_102), .O(gate33inter3));
  inv1  gate1265(.a(s_103), .O(gate33inter4));
  nand2 gate1266(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1267(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1268(.a(G17), .O(gate33inter7));
  inv1  gate1269(.a(G21), .O(gate33inter8));
  nand2 gate1270(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1271(.a(s_103), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1272(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1273(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1274(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate869(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate870(.a(gate36inter0), .b(s_46), .O(gate36inter1));
  and2  gate871(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate872(.a(s_46), .O(gate36inter3));
  inv1  gate873(.a(s_47), .O(gate36inter4));
  nand2 gate874(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate875(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate876(.a(G26), .O(gate36inter7));
  inv1  gate877(.a(G30), .O(gate36inter8));
  nand2 gate878(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate879(.a(s_47), .b(gate36inter3), .O(gate36inter10));
  nor2  gate880(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate881(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate882(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1023(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1024(.a(gate38inter0), .b(s_68), .O(gate38inter1));
  and2  gate1025(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1026(.a(s_68), .O(gate38inter3));
  inv1  gate1027(.a(s_69), .O(gate38inter4));
  nand2 gate1028(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1029(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1030(.a(G27), .O(gate38inter7));
  inv1  gate1031(.a(G31), .O(gate38inter8));
  nand2 gate1032(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1033(.a(s_69), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1034(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1035(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1036(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate561(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate562(.a(gate39inter0), .b(s_2), .O(gate39inter1));
  and2  gate563(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate564(.a(s_2), .O(gate39inter3));
  inv1  gate565(.a(s_3), .O(gate39inter4));
  nand2 gate566(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate567(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate568(.a(G20), .O(gate39inter7));
  inv1  gate569(.a(G24), .O(gate39inter8));
  nand2 gate570(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate571(.a(s_3), .b(gate39inter3), .O(gate39inter10));
  nor2  gate572(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate573(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate574(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1499(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1500(.a(gate43inter0), .b(s_136), .O(gate43inter1));
  and2  gate1501(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1502(.a(s_136), .O(gate43inter3));
  inv1  gate1503(.a(s_137), .O(gate43inter4));
  nand2 gate1504(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1505(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1506(.a(G3), .O(gate43inter7));
  inv1  gate1507(.a(G269), .O(gate43inter8));
  nand2 gate1508(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1509(.a(s_137), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1510(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1511(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1512(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate2073(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2074(.a(gate45inter0), .b(s_218), .O(gate45inter1));
  and2  gate2075(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2076(.a(s_218), .O(gate45inter3));
  inv1  gate2077(.a(s_219), .O(gate45inter4));
  nand2 gate2078(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2079(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2080(.a(G5), .O(gate45inter7));
  inv1  gate2081(.a(G272), .O(gate45inter8));
  nand2 gate2082(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2083(.a(s_219), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2084(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2085(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2086(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate953(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate954(.a(gate46inter0), .b(s_58), .O(gate46inter1));
  and2  gate955(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate956(.a(s_58), .O(gate46inter3));
  inv1  gate957(.a(s_59), .O(gate46inter4));
  nand2 gate958(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate959(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate960(.a(G6), .O(gate46inter7));
  inv1  gate961(.a(G272), .O(gate46inter8));
  nand2 gate962(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate963(.a(s_59), .b(gate46inter3), .O(gate46inter10));
  nor2  gate964(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate965(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate966(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1247(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1248(.a(gate48inter0), .b(s_100), .O(gate48inter1));
  and2  gate1249(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1250(.a(s_100), .O(gate48inter3));
  inv1  gate1251(.a(s_101), .O(gate48inter4));
  nand2 gate1252(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1253(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1254(.a(G8), .O(gate48inter7));
  inv1  gate1255(.a(G275), .O(gate48inter8));
  nand2 gate1256(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1257(.a(s_101), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1258(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1259(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1260(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1723(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1724(.a(gate55inter0), .b(s_168), .O(gate55inter1));
  and2  gate1725(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1726(.a(s_168), .O(gate55inter3));
  inv1  gate1727(.a(s_169), .O(gate55inter4));
  nand2 gate1728(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1729(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1730(.a(G15), .O(gate55inter7));
  inv1  gate1731(.a(G287), .O(gate55inter8));
  nand2 gate1732(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1733(.a(s_169), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1734(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1735(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1736(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1667(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1668(.a(gate57inter0), .b(s_160), .O(gate57inter1));
  and2  gate1669(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1670(.a(s_160), .O(gate57inter3));
  inv1  gate1671(.a(s_161), .O(gate57inter4));
  nand2 gate1672(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1673(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1674(.a(G17), .O(gate57inter7));
  inv1  gate1675(.a(G290), .O(gate57inter8));
  nand2 gate1676(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1677(.a(s_161), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1678(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1679(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1680(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1555(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1556(.a(gate60inter0), .b(s_144), .O(gate60inter1));
  and2  gate1557(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1558(.a(s_144), .O(gate60inter3));
  inv1  gate1559(.a(s_145), .O(gate60inter4));
  nand2 gate1560(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1561(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1562(.a(G20), .O(gate60inter7));
  inv1  gate1563(.a(G293), .O(gate60inter8));
  nand2 gate1564(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1565(.a(s_145), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1566(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1567(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1568(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1037(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1038(.a(gate63inter0), .b(s_70), .O(gate63inter1));
  and2  gate1039(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1040(.a(s_70), .O(gate63inter3));
  inv1  gate1041(.a(s_71), .O(gate63inter4));
  nand2 gate1042(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1043(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1044(.a(G23), .O(gate63inter7));
  inv1  gate1045(.a(G299), .O(gate63inter8));
  nand2 gate1046(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1047(.a(s_71), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1048(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1049(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1050(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1387(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1388(.a(gate64inter0), .b(s_120), .O(gate64inter1));
  and2  gate1389(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1390(.a(s_120), .O(gate64inter3));
  inv1  gate1391(.a(s_121), .O(gate64inter4));
  nand2 gate1392(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1393(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1394(.a(G24), .O(gate64inter7));
  inv1  gate1395(.a(G299), .O(gate64inter8));
  nand2 gate1396(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1397(.a(s_121), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1398(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1399(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1400(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1905(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1906(.a(gate65inter0), .b(s_194), .O(gate65inter1));
  and2  gate1907(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1908(.a(s_194), .O(gate65inter3));
  inv1  gate1909(.a(s_195), .O(gate65inter4));
  nand2 gate1910(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1911(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1912(.a(G25), .O(gate65inter7));
  inv1  gate1913(.a(G302), .O(gate65inter8));
  nand2 gate1914(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1915(.a(s_195), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1916(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1917(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1918(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1457(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1458(.a(gate69inter0), .b(s_130), .O(gate69inter1));
  and2  gate1459(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1460(.a(s_130), .O(gate69inter3));
  inv1  gate1461(.a(s_131), .O(gate69inter4));
  nand2 gate1462(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1463(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1464(.a(G29), .O(gate69inter7));
  inv1  gate1465(.a(G308), .O(gate69inter8));
  nand2 gate1466(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1467(.a(s_131), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1468(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1469(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1470(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1359(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1360(.a(gate70inter0), .b(s_116), .O(gate70inter1));
  and2  gate1361(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1362(.a(s_116), .O(gate70inter3));
  inv1  gate1363(.a(s_117), .O(gate70inter4));
  nand2 gate1364(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1365(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1366(.a(G30), .O(gate70inter7));
  inv1  gate1367(.a(G308), .O(gate70inter8));
  nand2 gate1368(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1369(.a(s_117), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1370(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1371(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1372(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2059(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2060(.a(gate74inter0), .b(s_216), .O(gate74inter1));
  and2  gate2061(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2062(.a(s_216), .O(gate74inter3));
  inv1  gate2063(.a(s_217), .O(gate74inter4));
  nand2 gate2064(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2065(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2066(.a(G5), .O(gate74inter7));
  inv1  gate2067(.a(G314), .O(gate74inter8));
  nand2 gate2068(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2069(.a(s_217), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2070(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2071(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2072(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate617(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate618(.a(gate76inter0), .b(s_10), .O(gate76inter1));
  and2  gate619(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate620(.a(s_10), .O(gate76inter3));
  inv1  gate621(.a(s_11), .O(gate76inter4));
  nand2 gate622(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate623(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate624(.a(G13), .O(gate76inter7));
  inv1  gate625(.a(G317), .O(gate76inter8));
  nand2 gate626(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate627(.a(s_11), .b(gate76inter3), .O(gate76inter10));
  nor2  gate628(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate629(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate630(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate701(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate702(.a(gate102inter0), .b(s_22), .O(gate102inter1));
  and2  gate703(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate704(.a(s_22), .O(gate102inter3));
  inv1  gate705(.a(s_23), .O(gate102inter4));
  nand2 gate706(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate707(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate708(.a(G24), .O(gate102inter7));
  inv1  gate709(.a(G356), .O(gate102inter8));
  nand2 gate710(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate711(.a(s_23), .b(gate102inter3), .O(gate102inter10));
  nor2  gate712(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate713(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate714(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1765(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1766(.a(gate113inter0), .b(s_174), .O(gate113inter1));
  and2  gate1767(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1768(.a(s_174), .O(gate113inter3));
  inv1  gate1769(.a(s_175), .O(gate113inter4));
  nand2 gate1770(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1771(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1772(.a(G378), .O(gate113inter7));
  inv1  gate1773(.a(G379), .O(gate113inter8));
  nand2 gate1774(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1775(.a(s_175), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1776(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1777(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1778(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate1079(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1080(.a(gate114inter0), .b(s_76), .O(gate114inter1));
  and2  gate1081(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1082(.a(s_76), .O(gate114inter3));
  inv1  gate1083(.a(s_77), .O(gate114inter4));
  nand2 gate1084(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1085(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1086(.a(G380), .O(gate114inter7));
  inv1  gate1087(.a(G381), .O(gate114inter8));
  nand2 gate1088(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1089(.a(s_77), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1090(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1091(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1092(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate855(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate856(.a(gate126inter0), .b(s_44), .O(gate126inter1));
  and2  gate857(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate858(.a(s_44), .O(gate126inter3));
  inv1  gate859(.a(s_45), .O(gate126inter4));
  nand2 gate860(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate861(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate862(.a(G404), .O(gate126inter7));
  inv1  gate863(.a(G405), .O(gate126inter8));
  nand2 gate864(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate865(.a(s_45), .b(gate126inter3), .O(gate126inter10));
  nor2  gate866(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate867(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate868(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1989(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1990(.a(gate131inter0), .b(s_206), .O(gate131inter1));
  and2  gate1991(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1992(.a(s_206), .O(gate131inter3));
  inv1  gate1993(.a(s_207), .O(gate131inter4));
  nand2 gate1994(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1995(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1996(.a(G414), .O(gate131inter7));
  inv1  gate1997(.a(G415), .O(gate131inter8));
  nand2 gate1998(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1999(.a(s_207), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2000(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2001(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2002(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate645(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate646(.a(gate138inter0), .b(s_14), .O(gate138inter1));
  and2  gate647(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate648(.a(s_14), .O(gate138inter3));
  inv1  gate649(.a(s_15), .O(gate138inter4));
  nand2 gate650(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate651(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate652(.a(G432), .O(gate138inter7));
  inv1  gate653(.a(G435), .O(gate138inter8));
  nand2 gate654(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate655(.a(s_15), .b(gate138inter3), .O(gate138inter10));
  nor2  gate656(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate657(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate658(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate967(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate968(.a(gate139inter0), .b(s_60), .O(gate139inter1));
  and2  gate969(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate970(.a(s_60), .O(gate139inter3));
  inv1  gate971(.a(s_61), .O(gate139inter4));
  nand2 gate972(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate973(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate974(.a(G438), .O(gate139inter7));
  inv1  gate975(.a(G441), .O(gate139inter8));
  nand2 gate976(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate977(.a(s_61), .b(gate139inter3), .O(gate139inter10));
  nor2  gate978(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate979(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate980(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1303(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1304(.a(gate140inter0), .b(s_108), .O(gate140inter1));
  and2  gate1305(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1306(.a(s_108), .O(gate140inter3));
  inv1  gate1307(.a(s_109), .O(gate140inter4));
  nand2 gate1308(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1309(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1310(.a(G444), .O(gate140inter7));
  inv1  gate1311(.a(G447), .O(gate140inter8));
  nand2 gate1312(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1313(.a(s_109), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1314(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1315(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1316(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1569(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1570(.a(gate154inter0), .b(s_146), .O(gate154inter1));
  and2  gate1571(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1572(.a(s_146), .O(gate154inter3));
  inv1  gate1573(.a(s_147), .O(gate154inter4));
  nand2 gate1574(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1575(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1576(.a(G429), .O(gate154inter7));
  inv1  gate1577(.a(G522), .O(gate154inter8));
  nand2 gate1578(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1579(.a(s_147), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1580(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1581(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1582(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1527(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1528(.a(gate164inter0), .b(s_140), .O(gate164inter1));
  and2  gate1529(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1530(.a(s_140), .O(gate164inter3));
  inv1  gate1531(.a(s_141), .O(gate164inter4));
  nand2 gate1532(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1533(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1534(.a(G459), .O(gate164inter7));
  inv1  gate1535(.a(G537), .O(gate164inter8));
  nand2 gate1536(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1537(.a(s_141), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1538(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1539(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1540(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1485(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1486(.a(gate179inter0), .b(s_134), .O(gate179inter1));
  and2  gate1487(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1488(.a(s_134), .O(gate179inter3));
  inv1  gate1489(.a(s_135), .O(gate179inter4));
  nand2 gate1490(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1491(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1492(.a(G504), .O(gate179inter7));
  inv1  gate1493(.a(G561), .O(gate179inter8));
  nand2 gate1494(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1495(.a(s_135), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1496(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1497(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1498(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate2087(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2088(.a(gate182inter0), .b(s_220), .O(gate182inter1));
  and2  gate2089(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2090(.a(s_220), .O(gate182inter3));
  inv1  gate2091(.a(s_221), .O(gate182inter4));
  nand2 gate2092(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2093(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2094(.a(G513), .O(gate182inter7));
  inv1  gate2095(.a(G564), .O(gate182inter8));
  nand2 gate2096(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2097(.a(s_221), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2098(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2099(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2100(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1541(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1542(.a(gate183inter0), .b(s_142), .O(gate183inter1));
  and2  gate1543(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1544(.a(s_142), .O(gate183inter3));
  inv1  gate1545(.a(s_143), .O(gate183inter4));
  nand2 gate1546(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1547(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1548(.a(G516), .O(gate183inter7));
  inv1  gate1549(.a(G567), .O(gate183inter8));
  nand2 gate1550(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1551(.a(s_143), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1552(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1553(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1554(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate757(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate758(.a(gate184inter0), .b(s_30), .O(gate184inter1));
  and2  gate759(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate760(.a(s_30), .O(gate184inter3));
  inv1  gate761(.a(s_31), .O(gate184inter4));
  nand2 gate762(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate763(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate764(.a(G519), .O(gate184inter7));
  inv1  gate765(.a(G567), .O(gate184inter8));
  nand2 gate766(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate767(.a(s_31), .b(gate184inter3), .O(gate184inter10));
  nor2  gate768(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate769(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate770(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1947(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1948(.a(gate185inter0), .b(s_200), .O(gate185inter1));
  and2  gate1949(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1950(.a(s_200), .O(gate185inter3));
  inv1  gate1951(.a(s_201), .O(gate185inter4));
  nand2 gate1952(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1953(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1954(.a(G570), .O(gate185inter7));
  inv1  gate1955(.a(G571), .O(gate185inter8));
  nand2 gate1956(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1957(.a(s_201), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1958(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1959(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1960(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate743(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate744(.a(gate189inter0), .b(s_28), .O(gate189inter1));
  and2  gate745(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate746(.a(s_28), .O(gate189inter3));
  inv1  gate747(.a(s_29), .O(gate189inter4));
  nand2 gate748(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate749(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate750(.a(G578), .O(gate189inter7));
  inv1  gate751(.a(G579), .O(gate189inter8));
  nand2 gate752(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate753(.a(s_29), .b(gate189inter3), .O(gate189inter10));
  nor2  gate754(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate755(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate756(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1289(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1290(.a(gate190inter0), .b(s_106), .O(gate190inter1));
  and2  gate1291(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1292(.a(s_106), .O(gate190inter3));
  inv1  gate1293(.a(s_107), .O(gate190inter4));
  nand2 gate1294(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1295(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1296(.a(G580), .O(gate190inter7));
  inv1  gate1297(.a(G581), .O(gate190inter8));
  nand2 gate1298(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1299(.a(s_107), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1300(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1301(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1302(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate631(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate632(.a(gate191inter0), .b(s_12), .O(gate191inter1));
  and2  gate633(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate634(.a(s_12), .O(gate191inter3));
  inv1  gate635(.a(s_13), .O(gate191inter4));
  nand2 gate636(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate637(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate638(.a(G582), .O(gate191inter7));
  inv1  gate639(.a(G583), .O(gate191inter8));
  nand2 gate640(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate641(.a(s_13), .b(gate191inter3), .O(gate191inter10));
  nor2  gate642(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate643(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate644(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1429(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1430(.a(gate195inter0), .b(s_126), .O(gate195inter1));
  and2  gate1431(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1432(.a(s_126), .O(gate195inter3));
  inv1  gate1433(.a(s_127), .O(gate195inter4));
  nand2 gate1434(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1435(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1436(.a(G590), .O(gate195inter7));
  inv1  gate1437(.a(G591), .O(gate195inter8));
  nand2 gate1438(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1439(.a(s_127), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1440(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1441(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1442(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1051(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1052(.a(gate197inter0), .b(s_72), .O(gate197inter1));
  and2  gate1053(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1054(.a(s_72), .O(gate197inter3));
  inv1  gate1055(.a(s_73), .O(gate197inter4));
  nand2 gate1056(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1057(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1058(.a(G594), .O(gate197inter7));
  inv1  gate1059(.a(G595), .O(gate197inter8));
  nand2 gate1060(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1061(.a(s_73), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1062(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1063(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1064(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate883(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate884(.a(gate199inter0), .b(s_48), .O(gate199inter1));
  and2  gate885(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate886(.a(s_48), .O(gate199inter3));
  inv1  gate887(.a(s_49), .O(gate199inter4));
  nand2 gate888(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate889(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate890(.a(G598), .O(gate199inter7));
  inv1  gate891(.a(G599), .O(gate199inter8));
  nand2 gate892(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate893(.a(s_49), .b(gate199inter3), .O(gate199inter10));
  nor2  gate894(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate895(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate896(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1933(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1934(.a(gate201inter0), .b(s_198), .O(gate201inter1));
  and2  gate1935(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1936(.a(s_198), .O(gate201inter3));
  inv1  gate1937(.a(s_199), .O(gate201inter4));
  nand2 gate1938(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1939(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1940(.a(G602), .O(gate201inter7));
  inv1  gate1941(.a(G607), .O(gate201inter8));
  nand2 gate1942(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1943(.a(s_199), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1944(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1945(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1946(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1975(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1976(.a(gate212inter0), .b(s_204), .O(gate212inter1));
  and2  gate1977(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1978(.a(s_204), .O(gate212inter3));
  inv1  gate1979(.a(s_205), .O(gate212inter4));
  nand2 gate1980(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1981(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1982(.a(G617), .O(gate212inter7));
  inv1  gate1983(.a(G669), .O(gate212inter8));
  nand2 gate1984(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1985(.a(s_205), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1986(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1987(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1988(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1751(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1752(.a(gate223inter0), .b(s_172), .O(gate223inter1));
  and2  gate1753(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1754(.a(s_172), .O(gate223inter3));
  inv1  gate1755(.a(s_173), .O(gate223inter4));
  nand2 gate1756(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1757(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1758(.a(G627), .O(gate223inter7));
  inv1  gate1759(.a(G687), .O(gate223inter8));
  nand2 gate1760(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1761(.a(s_173), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1762(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1763(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1764(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1401(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1402(.a(gate226inter0), .b(s_122), .O(gate226inter1));
  and2  gate1403(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1404(.a(s_122), .O(gate226inter3));
  inv1  gate1405(.a(s_123), .O(gate226inter4));
  nand2 gate1406(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1407(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1408(.a(G692), .O(gate226inter7));
  inv1  gate1409(.a(G693), .O(gate226inter8));
  nand2 gate1410(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1411(.a(s_123), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1412(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1413(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1414(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate785(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate786(.a(gate227inter0), .b(s_34), .O(gate227inter1));
  and2  gate787(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate788(.a(s_34), .O(gate227inter3));
  inv1  gate789(.a(s_35), .O(gate227inter4));
  nand2 gate790(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate791(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate792(.a(G694), .O(gate227inter7));
  inv1  gate793(.a(G695), .O(gate227inter8));
  nand2 gate794(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate795(.a(s_35), .b(gate227inter3), .O(gate227inter10));
  nor2  gate796(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate797(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate798(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1065(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1066(.a(gate234inter0), .b(s_74), .O(gate234inter1));
  and2  gate1067(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1068(.a(s_74), .O(gate234inter3));
  inv1  gate1069(.a(s_75), .O(gate234inter4));
  nand2 gate1070(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1071(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1072(.a(G245), .O(gate234inter7));
  inv1  gate1073(.a(G721), .O(gate234inter8));
  nand2 gate1074(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1075(.a(s_75), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1076(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1077(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1078(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1373(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1374(.a(gate235inter0), .b(s_118), .O(gate235inter1));
  and2  gate1375(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1376(.a(s_118), .O(gate235inter3));
  inv1  gate1377(.a(s_119), .O(gate235inter4));
  nand2 gate1378(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1379(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1380(.a(G248), .O(gate235inter7));
  inv1  gate1381(.a(G724), .O(gate235inter8));
  nand2 gate1382(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1383(.a(s_119), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1384(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1385(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1386(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate1345(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1346(.a(gate236inter0), .b(s_114), .O(gate236inter1));
  and2  gate1347(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1348(.a(s_114), .O(gate236inter3));
  inv1  gate1349(.a(s_115), .O(gate236inter4));
  nand2 gate1350(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1351(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1352(.a(G251), .O(gate236inter7));
  inv1  gate1353(.a(G727), .O(gate236inter8));
  nand2 gate1354(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1355(.a(s_115), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1356(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1357(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1358(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1849(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1850(.a(gate239inter0), .b(s_186), .O(gate239inter1));
  and2  gate1851(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1852(.a(s_186), .O(gate239inter3));
  inv1  gate1853(.a(s_187), .O(gate239inter4));
  nand2 gate1854(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1855(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1856(.a(G260), .O(gate239inter7));
  inv1  gate1857(.a(G712), .O(gate239inter8));
  nand2 gate1858(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1859(.a(s_187), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1860(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1861(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1862(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1149(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1150(.a(gate243inter0), .b(s_86), .O(gate243inter1));
  and2  gate1151(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1152(.a(s_86), .O(gate243inter3));
  inv1  gate1153(.a(s_87), .O(gate243inter4));
  nand2 gate1154(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1155(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1156(.a(G245), .O(gate243inter7));
  inv1  gate1157(.a(G733), .O(gate243inter8));
  nand2 gate1158(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1159(.a(s_87), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1160(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1161(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1162(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1639(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1640(.a(gate246inter0), .b(s_156), .O(gate246inter1));
  and2  gate1641(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1642(.a(s_156), .O(gate246inter3));
  inv1  gate1643(.a(s_157), .O(gate246inter4));
  nand2 gate1644(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1645(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1646(.a(G724), .O(gate246inter7));
  inv1  gate1647(.a(G736), .O(gate246inter8));
  nand2 gate1648(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1649(.a(s_157), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1650(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1651(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1652(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate547(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate548(.a(gate247inter0), .b(s_0), .O(gate247inter1));
  and2  gate549(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate550(.a(s_0), .O(gate247inter3));
  inv1  gate551(.a(s_1), .O(gate247inter4));
  nand2 gate552(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate553(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate554(.a(G251), .O(gate247inter7));
  inv1  gate555(.a(G739), .O(gate247inter8));
  nand2 gate556(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate557(.a(s_1), .b(gate247inter3), .O(gate247inter10));
  nor2  gate558(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate559(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate560(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1779(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1780(.a(gate249inter0), .b(s_176), .O(gate249inter1));
  and2  gate1781(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1782(.a(s_176), .O(gate249inter3));
  inv1  gate1783(.a(s_177), .O(gate249inter4));
  nand2 gate1784(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1785(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1786(.a(G254), .O(gate249inter7));
  inv1  gate1787(.a(G742), .O(gate249inter8));
  nand2 gate1788(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1789(.a(s_177), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1790(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1791(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1792(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1163(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1164(.a(gate253inter0), .b(s_88), .O(gate253inter1));
  and2  gate1165(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1166(.a(s_88), .O(gate253inter3));
  inv1  gate1167(.a(s_89), .O(gate253inter4));
  nand2 gate1168(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1169(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1170(.a(G260), .O(gate253inter7));
  inv1  gate1171(.a(G748), .O(gate253inter8));
  nand2 gate1172(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1173(.a(s_89), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1174(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1175(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1176(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1093(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1094(.a(gate254inter0), .b(s_78), .O(gate254inter1));
  and2  gate1095(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1096(.a(s_78), .O(gate254inter3));
  inv1  gate1097(.a(s_79), .O(gate254inter4));
  nand2 gate1098(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1099(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1100(.a(G712), .O(gate254inter7));
  inv1  gate1101(.a(G748), .O(gate254inter8));
  nand2 gate1102(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1103(.a(s_79), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1104(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1105(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1106(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate911(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate912(.a(gate255inter0), .b(s_52), .O(gate255inter1));
  and2  gate913(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate914(.a(s_52), .O(gate255inter3));
  inv1  gate915(.a(s_53), .O(gate255inter4));
  nand2 gate916(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate917(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate918(.a(G263), .O(gate255inter7));
  inv1  gate919(.a(G751), .O(gate255inter8));
  nand2 gate920(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate921(.a(s_53), .b(gate255inter3), .O(gate255inter10));
  nor2  gate922(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate923(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate924(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1695(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1696(.a(gate260inter0), .b(s_164), .O(gate260inter1));
  and2  gate1697(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1698(.a(s_164), .O(gate260inter3));
  inv1  gate1699(.a(s_165), .O(gate260inter4));
  nand2 gate1700(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1701(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1702(.a(G760), .O(gate260inter7));
  inv1  gate1703(.a(G761), .O(gate260inter8));
  nand2 gate1704(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1705(.a(s_165), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1706(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1707(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1708(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1443(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1444(.a(gate263inter0), .b(s_128), .O(gate263inter1));
  and2  gate1445(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1446(.a(s_128), .O(gate263inter3));
  inv1  gate1447(.a(s_129), .O(gate263inter4));
  nand2 gate1448(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1449(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1450(.a(G766), .O(gate263inter7));
  inv1  gate1451(.a(G767), .O(gate263inter8));
  nand2 gate1452(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1453(.a(s_129), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1454(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1455(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1456(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1177(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1178(.a(gate271inter0), .b(s_90), .O(gate271inter1));
  and2  gate1179(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1180(.a(s_90), .O(gate271inter3));
  inv1  gate1181(.a(s_91), .O(gate271inter4));
  nand2 gate1182(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1183(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1184(.a(G660), .O(gate271inter7));
  inv1  gate1185(.a(G788), .O(gate271inter8));
  nand2 gate1186(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1187(.a(s_91), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1188(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1189(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1190(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate729(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate730(.a(gate274inter0), .b(s_26), .O(gate274inter1));
  and2  gate731(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate732(.a(s_26), .O(gate274inter3));
  inv1  gate733(.a(s_27), .O(gate274inter4));
  nand2 gate734(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate735(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate736(.a(G770), .O(gate274inter7));
  inv1  gate737(.a(G794), .O(gate274inter8));
  nand2 gate738(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate739(.a(s_27), .b(gate274inter3), .O(gate274inter10));
  nor2  gate740(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate741(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate742(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1863(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1864(.a(gate275inter0), .b(s_188), .O(gate275inter1));
  and2  gate1865(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1866(.a(s_188), .O(gate275inter3));
  inv1  gate1867(.a(s_189), .O(gate275inter4));
  nand2 gate1868(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1869(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1870(.a(G645), .O(gate275inter7));
  inv1  gate1871(.a(G797), .O(gate275inter8));
  nand2 gate1872(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1873(.a(s_189), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1874(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1875(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1876(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1807(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1808(.a(gate276inter0), .b(s_180), .O(gate276inter1));
  and2  gate1809(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1810(.a(s_180), .O(gate276inter3));
  inv1  gate1811(.a(s_181), .O(gate276inter4));
  nand2 gate1812(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1813(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1814(.a(G773), .O(gate276inter7));
  inv1  gate1815(.a(G797), .O(gate276inter8));
  nand2 gate1816(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1817(.a(s_181), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1818(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1819(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1820(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate575(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate576(.a(gate279inter0), .b(s_4), .O(gate279inter1));
  and2  gate577(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate578(.a(s_4), .O(gate279inter3));
  inv1  gate579(.a(s_5), .O(gate279inter4));
  nand2 gate580(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate581(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate582(.a(G651), .O(gate279inter7));
  inv1  gate583(.a(G803), .O(gate279inter8));
  nand2 gate584(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate585(.a(s_5), .b(gate279inter3), .O(gate279inter10));
  nor2  gate586(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate587(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate588(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate715(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate716(.a(gate282inter0), .b(s_24), .O(gate282inter1));
  and2  gate717(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate718(.a(s_24), .O(gate282inter3));
  inv1  gate719(.a(s_25), .O(gate282inter4));
  nand2 gate720(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate721(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate722(.a(G782), .O(gate282inter7));
  inv1  gate723(.a(G806), .O(gate282inter8));
  nand2 gate724(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate725(.a(s_25), .b(gate282inter3), .O(gate282inter10));
  nor2  gate726(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate727(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate728(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate925(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate926(.a(gate285inter0), .b(s_54), .O(gate285inter1));
  and2  gate927(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate928(.a(s_54), .O(gate285inter3));
  inv1  gate929(.a(s_55), .O(gate285inter4));
  nand2 gate930(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate931(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate932(.a(G660), .O(gate285inter7));
  inv1  gate933(.a(G812), .O(gate285inter8));
  nand2 gate934(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate935(.a(s_55), .b(gate285inter3), .O(gate285inter10));
  nor2  gate936(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate937(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate938(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1961(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1962(.a(gate287inter0), .b(s_202), .O(gate287inter1));
  and2  gate1963(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1964(.a(s_202), .O(gate287inter3));
  inv1  gate1965(.a(s_203), .O(gate287inter4));
  nand2 gate1966(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1967(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1968(.a(G663), .O(gate287inter7));
  inv1  gate1969(.a(G815), .O(gate287inter8));
  nand2 gate1970(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1971(.a(s_203), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1972(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1973(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1974(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate2003(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2004(.a(gate288inter0), .b(s_208), .O(gate288inter1));
  and2  gate2005(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2006(.a(s_208), .O(gate288inter3));
  inv1  gate2007(.a(s_209), .O(gate288inter4));
  nand2 gate2008(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2009(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2010(.a(G791), .O(gate288inter7));
  inv1  gate2011(.a(G815), .O(gate288inter8));
  nand2 gate2012(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2013(.a(s_209), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2014(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2015(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2016(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate687(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate688(.a(gate290inter0), .b(s_20), .O(gate290inter1));
  and2  gate689(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate690(.a(s_20), .O(gate290inter3));
  inv1  gate691(.a(s_21), .O(gate290inter4));
  nand2 gate692(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate693(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate694(.a(G820), .O(gate290inter7));
  inv1  gate695(.a(G821), .O(gate290inter8));
  nand2 gate696(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate697(.a(s_21), .b(gate290inter3), .O(gate290inter10));
  nor2  gate698(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate699(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate700(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1919(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1920(.a(gate295inter0), .b(s_196), .O(gate295inter1));
  and2  gate1921(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1922(.a(s_196), .O(gate295inter3));
  inv1  gate1923(.a(s_197), .O(gate295inter4));
  nand2 gate1924(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1925(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1926(.a(G830), .O(gate295inter7));
  inv1  gate1927(.a(G831), .O(gate295inter8));
  nand2 gate1928(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1929(.a(s_197), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1930(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1931(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1932(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1107(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1108(.a(gate296inter0), .b(s_80), .O(gate296inter1));
  and2  gate1109(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1110(.a(s_80), .O(gate296inter3));
  inv1  gate1111(.a(s_81), .O(gate296inter4));
  nand2 gate1112(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1113(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1114(.a(G826), .O(gate296inter7));
  inv1  gate1115(.a(G827), .O(gate296inter8));
  nand2 gate1116(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1117(.a(s_81), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1118(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1119(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1120(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1821(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1822(.a(gate389inter0), .b(s_182), .O(gate389inter1));
  and2  gate1823(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1824(.a(s_182), .O(gate389inter3));
  inv1  gate1825(.a(s_183), .O(gate389inter4));
  nand2 gate1826(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1827(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1828(.a(G3), .O(gate389inter7));
  inv1  gate1829(.a(G1042), .O(gate389inter8));
  nand2 gate1830(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1831(.a(s_183), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1832(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1833(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1834(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1891(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1892(.a(gate397inter0), .b(s_192), .O(gate397inter1));
  and2  gate1893(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1894(.a(s_192), .O(gate397inter3));
  inv1  gate1895(.a(s_193), .O(gate397inter4));
  nand2 gate1896(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1897(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1898(.a(G11), .O(gate397inter7));
  inv1  gate1899(.a(G1066), .O(gate397inter8));
  nand2 gate1900(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1901(.a(s_193), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1902(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1903(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1904(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate995(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate996(.a(gate404inter0), .b(s_64), .O(gate404inter1));
  and2  gate997(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate998(.a(s_64), .O(gate404inter3));
  inv1  gate999(.a(s_65), .O(gate404inter4));
  nand2 gate1000(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1001(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1002(.a(G18), .O(gate404inter7));
  inv1  gate1003(.a(G1087), .O(gate404inter8));
  nand2 gate1004(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1005(.a(s_65), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1006(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1007(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1008(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1415(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1416(.a(gate407inter0), .b(s_124), .O(gate407inter1));
  and2  gate1417(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1418(.a(s_124), .O(gate407inter3));
  inv1  gate1419(.a(s_125), .O(gate407inter4));
  nand2 gate1420(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1421(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1422(.a(G21), .O(gate407inter7));
  inv1  gate1423(.a(G1096), .O(gate407inter8));
  nand2 gate1424(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1425(.a(s_125), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1426(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1427(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1428(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1471(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1472(.a(gate420inter0), .b(s_132), .O(gate420inter1));
  and2  gate1473(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1474(.a(s_132), .O(gate420inter3));
  inv1  gate1475(.a(s_133), .O(gate420inter4));
  nand2 gate1476(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1477(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1478(.a(G1036), .O(gate420inter7));
  inv1  gate1479(.a(G1132), .O(gate420inter8));
  nand2 gate1480(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1481(.a(s_133), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1482(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1483(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1484(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1121(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1122(.a(gate422inter0), .b(s_82), .O(gate422inter1));
  and2  gate1123(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1124(.a(s_82), .O(gate422inter3));
  inv1  gate1125(.a(s_83), .O(gate422inter4));
  nand2 gate1126(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1127(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1128(.a(G1039), .O(gate422inter7));
  inv1  gate1129(.a(G1135), .O(gate422inter8));
  nand2 gate1130(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1131(.a(s_83), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1132(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1133(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1134(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2031(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2032(.a(gate425inter0), .b(s_212), .O(gate425inter1));
  and2  gate2033(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2034(.a(s_212), .O(gate425inter3));
  inv1  gate2035(.a(s_213), .O(gate425inter4));
  nand2 gate2036(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2037(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2038(.a(G4), .O(gate425inter7));
  inv1  gate2039(.a(G1141), .O(gate425inter8));
  nand2 gate2040(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2041(.a(s_213), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2042(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2043(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2044(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate897(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate898(.a(gate427inter0), .b(s_50), .O(gate427inter1));
  and2  gate899(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate900(.a(s_50), .O(gate427inter3));
  inv1  gate901(.a(s_51), .O(gate427inter4));
  nand2 gate902(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate903(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate904(.a(G5), .O(gate427inter7));
  inv1  gate905(.a(G1144), .O(gate427inter8));
  nand2 gate906(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate907(.a(s_51), .b(gate427inter3), .O(gate427inter10));
  nor2  gate908(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate909(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate910(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1233(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1234(.a(gate430inter0), .b(s_98), .O(gate430inter1));
  and2  gate1235(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1236(.a(s_98), .O(gate430inter3));
  inv1  gate1237(.a(s_99), .O(gate430inter4));
  nand2 gate1238(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1239(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1240(.a(G1051), .O(gate430inter7));
  inv1  gate1241(.a(G1147), .O(gate430inter8));
  nand2 gate1242(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1243(.a(s_99), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1244(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1245(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1246(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1317(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1318(.a(gate431inter0), .b(s_110), .O(gate431inter1));
  and2  gate1319(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1320(.a(s_110), .O(gate431inter3));
  inv1  gate1321(.a(s_111), .O(gate431inter4));
  nand2 gate1322(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1323(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1324(.a(G7), .O(gate431inter7));
  inv1  gate1325(.a(G1150), .O(gate431inter8));
  nand2 gate1326(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1327(.a(s_111), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1328(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1329(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1330(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1219(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1220(.a(gate434inter0), .b(s_96), .O(gate434inter1));
  and2  gate1221(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1222(.a(s_96), .O(gate434inter3));
  inv1  gate1223(.a(s_97), .O(gate434inter4));
  nand2 gate1224(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1225(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1226(.a(G1057), .O(gate434inter7));
  inv1  gate1227(.a(G1153), .O(gate434inter8));
  nand2 gate1228(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1229(.a(s_97), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1230(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1231(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1232(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1191(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1192(.a(gate439inter0), .b(s_92), .O(gate439inter1));
  and2  gate1193(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1194(.a(s_92), .O(gate439inter3));
  inv1  gate1195(.a(s_93), .O(gate439inter4));
  nand2 gate1196(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1197(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1198(.a(G11), .O(gate439inter7));
  inv1  gate1199(.a(G1162), .O(gate439inter8));
  nand2 gate1200(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1201(.a(s_93), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1202(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1203(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1204(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1331(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1332(.a(gate445inter0), .b(s_112), .O(gate445inter1));
  and2  gate1333(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1334(.a(s_112), .O(gate445inter3));
  inv1  gate1335(.a(s_113), .O(gate445inter4));
  nand2 gate1336(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1337(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1338(.a(G14), .O(gate445inter7));
  inv1  gate1339(.a(G1171), .O(gate445inter8));
  nand2 gate1340(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1341(.a(s_113), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1342(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1343(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1344(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate799(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate800(.a(gate446inter0), .b(s_36), .O(gate446inter1));
  and2  gate801(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate802(.a(s_36), .O(gate446inter3));
  inv1  gate803(.a(s_37), .O(gate446inter4));
  nand2 gate804(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate805(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate806(.a(G1075), .O(gate446inter7));
  inv1  gate807(.a(G1171), .O(gate446inter8));
  nand2 gate808(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate809(.a(s_37), .b(gate446inter3), .O(gate446inter10));
  nor2  gate810(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate811(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate812(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1275(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1276(.a(gate448inter0), .b(s_104), .O(gate448inter1));
  and2  gate1277(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1278(.a(s_104), .O(gate448inter3));
  inv1  gate1279(.a(s_105), .O(gate448inter4));
  nand2 gate1280(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1281(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1282(.a(G1078), .O(gate448inter7));
  inv1  gate1283(.a(G1174), .O(gate448inter8));
  nand2 gate1284(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1285(.a(s_105), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1286(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1287(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1288(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate603(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate604(.a(gate460inter0), .b(s_8), .O(gate460inter1));
  and2  gate605(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate606(.a(s_8), .O(gate460inter3));
  inv1  gate607(.a(s_9), .O(gate460inter4));
  nand2 gate608(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate609(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate610(.a(G1096), .O(gate460inter7));
  inv1  gate611(.a(G1192), .O(gate460inter8));
  nand2 gate612(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate613(.a(s_9), .b(gate460inter3), .O(gate460inter10));
  nor2  gate614(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate615(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate616(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1681(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1682(.a(gate462inter0), .b(s_162), .O(gate462inter1));
  and2  gate1683(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1684(.a(s_162), .O(gate462inter3));
  inv1  gate1685(.a(s_163), .O(gate462inter4));
  nand2 gate1686(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1687(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1688(.a(G1099), .O(gate462inter7));
  inv1  gate1689(.a(G1195), .O(gate462inter8));
  nand2 gate1690(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1691(.a(s_163), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1692(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1693(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1694(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate771(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate772(.a(gate464inter0), .b(s_32), .O(gate464inter1));
  and2  gate773(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate774(.a(s_32), .O(gate464inter3));
  inv1  gate775(.a(s_33), .O(gate464inter4));
  nand2 gate776(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate777(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate778(.a(G1102), .O(gate464inter7));
  inv1  gate779(.a(G1198), .O(gate464inter8));
  nand2 gate780(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate781(.a(s_33), .b(gate464inter3), .O(gate464inter10));
  nor2  gate782(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate783(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate784(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1653(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1654(.a(gate466inter0), .b(s_158), .O(gate466inter1));
  and2  gate1655(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1656(.a(s_158), .O(gate466inter3));
  inv1  gate1657(.a(s_159), .O(gate466inter4));
  nand2 gate1658(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1659(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1660(.a(G1105), .O(gate466inter7));
  inv1  gate1661(.a(G1201), .O(gate466inter8));
  nand2 gate1662(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1663(.a(s_159), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1664(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1665(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1666(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2017(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2018(.a(gate467inter0), .b(s_210), .O(gate467inter1));
  and2  gate2019(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2020(.a(s_210), .O(gate467inter3));
  inv1  gate2021(.a(s_211), .O(gate467inter4));
  nand2 gate2022(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2023(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2024(.a(G25), .O(gate467inter7));
  inv1  gate2025(.a(G1204), .O(gate467inter8));
  nand2 gate2026(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2027(.a(s_211), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2028(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2029(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2030(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1793(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1794(.a(gate469inter0), .b(s_178), .O(gate469inter1));
  and2  gate1795(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1796(.a(s_178), .O(gate469inter3));
  inv1  gate1797(.a(s_179), .O(gate469inter4));
  nand2 gate1798(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1799(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1800(.a(G26), .O(gate469inter7));
  inv1  gate1801(.a(G1207), .O(gate469inter8));
  nand2 gate1802(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1803(.a(s_179), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1804(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1805(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1806(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate659(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate660(.a(gate472inter0), .b(s_16), .O(gate472inter1));
  and2  gate661(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate662(.a(s_16), .O(gate472inter3));
  inv1  gate663(.a(s_17), .O(gate472inter4));
  nand2 gate664(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate665(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate666(.a(G1114), .O(gate472inter7));
  inv1  gate667(.a(G1210), .O(gate472inter8));
  nand2 gate668(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate669(.a(s_17), .b(gate472inter3), .O(gate472inter10));
  nor2  gate670(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate671(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate672(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1611(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1612(.a(gate474inter0), .b(s_152), .O(gate474inter1));
  and2  gate1613(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1614(.a(s_152), .O(gate474inter3));
  inv1  gate1615(.a(s_153), .O(gate474inter4));
  nand2 gate1616(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1617(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1618(.a(G1117), .O(gate474inter7));
  inv1  gate1619(.a(G1213), .O(gate474inter8));
  nand2 gate1620(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1621(.a(s_153), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1622(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1623(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1624(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1597(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1598(.a(gate480inter0), .b(s_150), .O(gate480inter1));
  and2  gate1599(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1600(.a(s_150), .O(gate480inter3));
  inv1  gate1601(.a(s_151), .O(gate480inter4));
  nand2 gate1602(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1603(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1604(.a(G1126), .O(gate480inter7));
  inv1  gate1605(.a(G1222), .O(gate480inter8));
  nand2 gate1606(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1607(.a(s_151), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1608(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1609(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1610(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1513(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1514(.a(gate481inter0), .b(s_138), .O(gate481inter1));
  and2  gate1515(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1516(.a(s_138), .O(gate481inter3));
  inv1  gate1517(.a(s_139), .O(gate481inter4));
  nand2 gate1518(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1519(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1520(.a(G32), .O(gate481inter7));
  inv1  gate1521(.a(G1225), .O(gate481inter8));
  nand2 gate1522(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1523(.a(s_139), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1524(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1525(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1526(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate813(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate814(.a(gate484inter0), .b(s_38), .O(gate484inter1));
  and2  gate815(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate816(.a(s_38), .O(gate484inter3));
  inv1  gate817(.a(s_39), .O(gate484inter4));
  nand2 gate818(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate819(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate820(.a(G1230), .O(gate484inter7));
  inv1  gate821(.a(G1231), .O(gate484inter8));
  nand2 gate822(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate823(.a(s_39), .b(gate484inter3), .O(gate484inter10));
  nor2  gate824(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate825(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate826(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1625(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1626(.a(gate485inter0), .b(s_154), .O(gate485inter1));
  and2  gate1627(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1628(.a(s_154), .O(gate485inter3));
  inv1  gate1629(.a(s_155), .O(gate485inter4));
  nand2 gate1630(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1631(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1632(.a(G1232), .O(gate485inter7));
  inv1  gate1633(.a(G1233), .O(gate485inter8));
  nand2 gate1634(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1635(.a(s_155), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1636(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1637(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1638(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1877(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1878(.a(gate486inter0), .b(s_190), .O(gate486inter1));
  and2  gate1879(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1880(.a(s_190), .O(gate486inter3));
  inv1  gate1881(.a(s_191), .O(gate486inter4));
  nand2 gate1882(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1883(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1884(.a(G1234), .O(gate486inter7));
  inv1  gate1885(.a(G1235), .O(gate486inter8));
  nand2 gate1886(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1887(.a(s_191), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1888(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1889(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1890(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1709(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1710(.a(gate490inter0), .b(s_166), .O(gate490inter1));
  and2  gate1711(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1712(.a(s_166), .O(gate490inter3));
  inv1  gate1713(.a(s_167), .O(gate490inter4));
  nand2 gate1714(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1715(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1716(.a(G1242), .O(gate490inter7));
  inv1  gate1717(.a(G1243), .O(gate490inter8));
  nand2 gate1718(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1719(.a(s_167), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1720(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1721(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1722(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1737(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1738(.a(gate495inter0), .b(s_170), .O(gate495inter1));
  and2  gate1739(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1740(.a(s_170), .O(gate495inter3));
  inv1  gate1741(.a(s_171), .O(gate495inter4));
  nand2 gate1742(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1743(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1744(.a(G1252), .O(gate495inter7));
  inv1  gate1745(.a(G1253), .O(gate495inter8));
  nand2 gate1746(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1747(.a(s_171), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1748(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1749(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1750(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate2045(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2046(.a(gate496inter0), .b(s_214), .O(gate496inter1));
  and2  gate2047(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2048(.a(s_214), .O(gate496inter3));
  inv1  gate2049(.a(s_215), .O(gate496inter4));
  nand2 gate2050(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2051(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2052(.a(G1254), .O(gate496inter7));
  inv1  gate2053(.a(G1255), .O(gate496inter8));
  nand2 gate2054(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2055(.a(s_215), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2056(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2057(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2058(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1583(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1584(.a(gate500inter0), .b(s_148), .O(gate500inter1));
  and2  gate1585(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1586(.a(s_148), .O(gate500inter3));
  inv1  gate1587(.a(s_149), .O(gate500inter4));
  nand2 gate1588(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1589(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1590(.a(G1262), .O(gate500inter7));
  inv1  gate1591(.a(G1263), .O(gate500inter8));
  nand2 gate1592(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1593(.a(s_149), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1594(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1595(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1596(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1835(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1836(.a(gate510inter0), .b(s_184), .O(gate510inter1));
  and2  gate1837(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1838(.a(s_184), .O(gate510inter3));
  inv1  gate1839(.a(s_185), .O(gate510inter4));
  nand2 gate1840(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1841(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1842(.a(G1282), .O(gate510inter7));
  inv1  gate1843(.a(G1283), .O(gate510inter8));
  nand2 gate1844(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1845(.a(s_185), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1846(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1847(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1848(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule