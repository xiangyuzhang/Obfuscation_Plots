module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1723(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1724(.a(gate12inter0), .b(s_168), .O(gate12inter1));
  and2  gate1725(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1726(.a(s_168), .O(gate12inter3));
  inv1  gate1727(.a(s_169), .O(gate12inter4));
  nand2 gate1728(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1729(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1730(.a(G7), .O(gate12inter7));
  inv1  gate1731(.a(G8), .O(gate12inter8));
  nand2 gate1732(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1733(.a(s_169), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1734(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1735(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1736(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1583(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1584(.a(gate16inter0), .b(s_148), .O(gate16inter1));
  and2  gate1585(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1586(.a(s_148), .O(gate16inter3));
  inv1  gate1587(.a(s_149), .O(gate16inter4));
  nand2 gate1588(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1589(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1590(.a(G15), .O(gate16inter7));
  inv1  gate1591(.a(G16), .O(gate16inter8));
  nand2 gate1592(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1593(.a(s_149), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1594(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1595(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1596(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate631(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate632(.a(gate18inter0), .b(s_12), .O(gate18inter1));
  and2  gate633(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate634(.a(s_12), .O(gate18inter3));
  inv1  gate635(.a(s_13), .O(gate18inter4));
  nand2 gate636(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate637(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate638(.a(G19), .O(gate18inter7));
  inv1  gate639(.a(G20), .O(gate18inter8));
  nand2 gate640(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate641(.a(s_13), .b(gate18inter3), .O(gate18inter10));
  nor2  gate642(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate643(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate644(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate855(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate856(.a(gate24inter0), .b(s_44), .O(gate24inter1));
  and2  gate857(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate858(.a(s_44), .O(gate24inter3));
  inv1  gate859(.a(s_45), .O(gate24inter4));
  nand2 gate860(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate861(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate862(.a(G31), .O(gate24inter7));
  inv1  gate863(.a(G32), .O(gate24inter8));
  nand2 gate864(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate865(.a(s_45), .b(gate24inter3), .O(gate24inter10));
  nor2  gate866(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate867(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate868(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1793(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1794(.a(gate32inter0), .b(s_178), .O(gate32inter1));
  and2  gate1795(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1796(.a(s_178), .O(gate32inter3));
  inv1  gate1797(.a(s_179), .O(gate32inter4));
  nand2 gate1798(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1799(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1800(.a(G12), .O(gate32inter7));
  inv1  gate1801(.a(G16), .O(gate32inter8));
  nand2 gate1802(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1803(.a(s_179), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1804(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1805(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1806(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1121(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1122(.a(gate33inter0), .b(s_82), .O(gate33inter1));
  and2  gate1123(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1124(.a(s_82), .O(gate33inter3));
  inv1  gate1125(.a(s_83), .O(gate33inter4));
  nand2 gate1126(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1127(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1128(.a(G17), .O(gate33inter7));
  inv1  gate1129(.a(G21), .O(gate33inter8));
  nand2 gate1130(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1131(.a(s_83), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1132(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1133(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1134(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1387(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1388(.a(gate39inter0), .b(s_120), .O(gate39inter1));
  and2  gate1389(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1390(.a(s_120), .O(gate39inter3));
  inv1  gate1391(.a(s_121), .O(gate39inter4));
  nand2 gate1392(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1393(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1394(.a(G20), .O(gate39inter7));
  inv1  gate1395(.a(G24), .O(gate39inter8));
  nand2 gate1396(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1397(.a(s_121), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1398(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1399(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1400(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1233(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1234(.a(gate41inter0), .b(s_98), .O(gate41inter1));
  and2  gate1235(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1236(.a(s_98), .O(gate41inter3));
  inv1  gate1237(.a(s_99), .O(gate41inter4));
  nand2 gate1238(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1239(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1240(.a(G1), .O(gate41inter7));
  inv1  gate1241(.a(G266), .O(gate41inter8));
  nand2 gate1242(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1243(.a(s_99), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1244(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1245(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1246(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1625(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1626(.a(gate43inter0), .b(s_154), .O(gate43inter1));
  and2  gate1627(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1628(.a(s_154), .O(gate43inter3));
  inv1  gate1629(.a(s_155), .O(gate43inter4));
  nand2 gate1630(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1631(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1632(.a(G3), .O(gate43inter7));
  inv1  gate1633(.a(G269), .O(gate43inter8));
  nand2 gate1634(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1635(.a(s_155), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1636(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1637(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1638(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate939(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate940(.a(gate46inter0), .b(s_56), .O(gate46inter1));
  and2  gate941(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate942(.a(s_56), .O(gate46inter3));
  inv1  gate943(.a(s_57), .O(gate46inter4));
  nand2 gate944(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate945(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate946(.a(G6), .O(gate46inter7));
  inv1  gate947(.a(G272), .O(gate46inter8));
  nand2 gate948(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate949(.a(s_57), .b(gate46inter3), .O(gate46inter10));
  nor2  gate950(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate951(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate952(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate883(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate884(.a(gate47inter0), .b(s_48), .O(gate47inter1));
  and2  gate885(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate886(.a(s_48), .O(gate47inter3));
  inv1  gate887(.a(s_49), .O(gate47inter4));
  nand2 gate888(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate889(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate890(.a(G7), .O(gate47inter7));
  inv1  gate891(.a(G275), .O(gate47inter8));
  nand2 gate892(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate893(.a(s_49), .b(gate47inter3), .O(gate47inter10));
  nor2  gate894(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate895(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate896(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate897(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate898(.a(gate50inter0), .b(s_50), .O(gate50inter1));
  and2  gate899(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate900(.a(s_50), .O(gate50inter3));
  inv1  gate901(.a(s_51), .O(gate50inter4));
  nand2 gate902(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate903(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate904(.a(G10), .O(gate50inter7));
  inv1  gate905(.a(G278), .O(gate50inter8));
  nand2 gate906(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate907(.a(s_51), .b(gate50inter3), .O(gate50inter10));
  nor2  gate908(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate909(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate910(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1821(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1822(.a(gate51inter0), .b(s_182), .O(gate51inter1));
  and2  gate1823(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1824(.a(s_182), .O(gate51inter3));
  inv1  gate1825(.a(s_183), .O(gate51inter4));
  nand2 gate1826(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1827(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1828(.a(G11), .O(gate51inter7));
  inv1  gate1829(.a(G281), .O(gate51inter8));
  nand2 gate1830(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1831(.a(s_183), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1832(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1833(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1834(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1471(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1472(.a(gate53inter0), .b(s_132), .O(gate53inter1));
  and2  gate1473(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1474(.a(s_132), .O(gate53inter3));
  inv1  gate1475(.a(s_133), .O(gate53inter4));
  nand2 gate1476(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1477(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1478(.a(G13), .O(gate53inter7));
  inv1  gate1479(.a(G284), .O(gate53inter8));
  nand2 gate1480(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1481(.a(s_133), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1482(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1483(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1484(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1611(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1612(.a(gate55inter0), .b(s_152), .O(gate55inter1));
  and2  gate1613(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1614(.a(s_152), .O(gate55inter3));
  inv1  gate1615(.a(s_153), .O(gate55inter4));
  nand2 gate1616(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1617(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1618(.a(G15), .O(gate55inter7));
  inv1  gate1619(.a(G287), .O(gate55inter8));
  nand2 gate1620(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1621(.a(s_153), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1622(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1623(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1624(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1107(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1108(.a(gate63inter0), .b(s_80), .O(gate63inter1));
  and2  gate1109(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1110(.a(s_80), .O(gate63inter3));
  inv1  gate1111(.a(s_81), .O(gate63inter4));
  nand2 gate1112(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1113(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1114(.a(G23), .O(gate63inter7));
  inv1  gate1115(.a(G299), .O(gate63inter8));
  nand2 gate1116(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1117(.a(s_81), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1118(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1119(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1120(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1065(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1066(.a(gate68inter0), .b(s_74), .O(gate68inter1));
  and2  gate1067(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1068(.a(s_74), .O(gate68inter3));
  inv1  gate1069(.a(s_75), .O(gate68inter4));
  nand2 gate1070(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1071(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1072(.a(G28), .O(gate68inter7));
  inv1  gate1073(.a(G305), .O(gate68inter8));
  nand2 gate1074(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1075(.a(s_75), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1076(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1077(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1078(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1737(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1738(.a(gate70inter0), .b(s_170), .O(gate70inter1));
  and2  gate1739(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1740(.a(s_170), .O(gate70inter3));
  inv1  gate1741(.a(s_171), .O(gate70inter4));
  nand2 gate1742(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1743(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1744(.a(G30), .O(gate70inter7));
  inv1  gate1745(.a(G308), .O(gate70inter8));
  nand2 gate1746(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1747(.a(s_171), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1748(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1749(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1750(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate827(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate828(.a(gate71inter0), .b(s_40), .O(gate71inter1));
  and2  gate829(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate830(.a(s_40), .O(gate71inter3));
  inv1  gate831(.a(s_41), .O(gate71inter4));
  nand2 gate832(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate833(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate834(.a(G31), .O(gate71inter7));
  inv1  gate835(.a(G311), .O(gate71inter8));
  nand2 gate836(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate837(.a(s_41), .b(gate71inter3), .O(gate71inter10));
  nor2  gate838(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate839(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate840(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate981(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate982(.a(gate80inter0), .b(s_62), .O(gate80inter1));
  and2  gate983(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate984(.a(s_62), .O(gate80inter3));
  inv1  gate985(.a(s_63), .O(gate80inter4));
  nand2 gate986(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate987(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate988(.a(G14), .O(gate80inter7));
  inv1  gate989(.a(G323), .O(gate80inter8));
  nand2 gate990(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate991(.a(s_63), .b(gate80inter3), .O(gate80inter10));
  nor2  gate992(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate993(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate994(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate617(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate618(.a(gate81inter0), .b(s_10), .O(gate81inter1));
  and2  gate619(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate620(.a(s_10), .O(gate81inter3));
  inv1  gate621(.a(s_11), .O(gate81inter4));
  nand2 gate622(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate623(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate624(.a(G3), .O(gate81inter7));
  inv1  gate625(.a(G326), .O(gate81inter8));
  nand2 gate626(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate627(.a(s_11), .b(gate81inter3), .O(gate81inter10));
  nor2  gate628(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate629(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate630(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1569(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1570(.a(gate83inter0), .b(s_146), .O(gate83inter1));
  and2  gate1571(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1572(.a(s_146), .O(gate83inter3));
  inv1  gate1573(.a(s_147), .O(gate83inter4));
  nand2 gate1574(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1575(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1576(.a(G11), .O(gate83inter7));
  inv1  gate1577(.a(G329), .O(gate83inter8));
  nand2 gate1578(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1579(.a(s_147), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1580(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1581(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1582(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1219(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1220(.a(gate86inter0), .b(s_96), .O(gate86inter1));
  and2  gate1221(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1222(.a(s_96), .O(gate86inter3));
  inv1  gate1223(.a(s_97), .O(gate86inter4));
  nand2 gate1224(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1225(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1226(.a(G8), .O(gate86inter7));
  inv1  gate1227(.a(G332), .O(gate86inter8));
  nand2 gate1228(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1229(.a(s_97), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1230(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1231(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1232(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1779(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1780(.a(gate87inter0), .b(s_176), .O(gate87inter1));
  and2  gate1781(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1782(.a(s_176), .O(gate87inter3));
  inv1  gate1783(.a(s_177), .O(gate87inter4));
  nand2 gate1784(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1785(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1786(.a(G12), .O(gate87inter7));
  inv1  gate1787(.a(G335), .O(gate87inter8));
  nand2 gate1788(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1789(.a(s_177), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1790(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1791(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1792(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1499(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1500(.a(gate97inter0), .b(s_136), .O(gate97inter1));
  and2  gate1501(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1502(.a(s_136), .O(gate97inter3));
  inv1  gate1503(.a(s_137), .O(gate97inter4));
  nand2 gate1504(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1505(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1506(.a(G19), .O(gate97inter7));
  inv1  gate1507(.a(G350), .O(gate97inter8));
  nand2 gate1508(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1509(.a(s_137), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1510(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1511(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1512(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1835(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1836(.a(gate98inter0), .b(s_184), .O(gate98inter1));
  and2  gate1837(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1838(.a(s_184), .O(gate98inter3));
  inv1  gate1839(.a(s_185), .O(gate98inter4));
  nand2 gate1840(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1841(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1842(.a(G23), .O(gate98inter7));
  inv1  gate1843(.a(G350), .O(gate98inter8));
  nand2 gate1844(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1845(.a(s_185), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1846(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1847(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1848(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1415(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1416(.a(gate103inter0), .b(s_124), .O(gate103inter1));
  and2  gate1417(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1418(.a(s_124), .O(gate103inter3));
  inv1  gate1419(.a(s_125), .O(gate103inter4));
  nand2 gate1420(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1421(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1422(.a(G28), .O(gate103inter7));
  inv1  gate1423(.a(G359), .O(gate103inter8));
  nand2 gate1424(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1425(.a(s_125), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1426(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1427(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1428(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1079(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1080(.a(gate104inter0), .b(s_76), .O(gate104inter1));
  and2  gate1081(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1082(.a(s_76), .O(gate104inter3));
  inv1  gate1083(.a(s_77), .O(gate104inter4));
  nand2 gate1084(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1085(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1086(.a(G32), .O(gate104inter7));
  inv1  gate1087(.a(G359), .O(gate104inter8));
  nand2 gate1088(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1089(.a(s_77), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1090(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1091(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1092(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1373(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1374(.a(gate107inter0), .b(s_118), .O(gate107inter1));
  and2  gate1375(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1376(.a(s_118), .O(gate107inter3));
  inv1  gate1377(.a(s_119), .O(gate107inter4));
  nand2 gate1378(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1379(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1380(.a(G366), .O(gate107inter7));
  inv1  gate1381(.a(G367), .O(gate107inter8));
  nand2 gate1382(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1383(.a(s_119), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1384(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1385(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1386(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate673(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate674(.a(gate110inter0), .b(s_18), .O(gate110inter1));
  and2  gate675(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate676(.a(s_18), .O(gate110inter3));
  inv1  gate677(.a(s_19), .O(gate110inter4));
  nand2 gate678(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate679(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate680(.a(G372), .O(gate110inter7));
  inv1  gate681(.a(G373), .O(gate110inter8));
  nand2 gate682(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate683(.a(s_19), .b(gate110inter3), .O(gate110inter10));
  nor2  gate684(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate685(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate686(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate575(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate576(.a(gate122inter0), .b(s_4), .O(gate122inter1));
  and2  gate577(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate578(.a(s_4), .O(gate122inter3));
  inv1  gate579(.a(s_5), .O(gate122inter4));
  nand2 gate580(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate581(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate582(.a(G396), .O(gate122inter7));
  inv1  gate583(.a(G397), .O(gate122inter8));
  nand2 gate584(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate585(.a(s_5), .b(gate122inter3), .O(gate122inter10));
  nor2  gate586(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate587(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate588(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1597(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1598(.a(gate126inter0), .b(s_150), .O(gate126inter1));
  and2  gate1599(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1600(.a(s_150), .O(gate126inter3));
  inv1  gate1601(.a(s_151), .O(gate126inter4));
  nand2 gate1602(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1603(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1604(.a(G404), .O(gate126inter7));
  inv1  gate1605(.a(G405), .O(gate126inter8));
  nand2 gate1606(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1607(.a(s_151), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1608(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1609(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1610(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1457(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1458(.a(gate127inter0), .b(s_130), .O(gate127inter1));
  and2  gate1459(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1460(.a(s_130), .O(gate127inter3));
  inv1  gate1461(.a(s_131), .O(gate127inter4));
  nand2 gate1462(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1463(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1464(.a(G406), .O(gate127inter7));
  inv1  gate1465(.a(G407), .O(gate127inter8));
  nand2 gate1466(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1467(.a(s_131), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1468(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1469(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1470(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1359(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1360(.a(gate136inter0), .b(s_116), .O(gate136inter1));
  and2  gate1361(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1362(.a(s_116), .O(gate136inter3));
  inv1  gate1363(.a(s_117), .O(gate136inter4));
  nand2 gate1364(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1365(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1366(.a(G424), .O(gate136inter7));
  inv1  gate1367(.a(G425), .O(gate136inter8));
  nand2 gate1368(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1369(.a(s_117), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1370(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1371(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1372(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate547(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate548(.a(gate137inter0), .b(s_0), .O(gate137inter1));
  and2  gate549(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate550(.a(s_0), .O(gate137inter3));
  inv1  gate551(.a(s_1), .O(gate137inter4));
  nand2 gate552(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate553(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate554(.a(G426), .O(gate137inter7));
  inv1  gate555(.a(G429), .O(gate137inter8));
  nand2 gate556(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate557(.a(s_1), .b(gate137inter3), .O(gate137inter10));
  nor2  gate558(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate559(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate560(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate729(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate730(.a(gate150inter0), .b(s_26), .O(gate150inter1));
  and2  gate731(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate732(.a(s_26), .O(gate150inter3));
  inv1  gate733(.a(s_27), .O(gate150inter4));
  nand2 gate734(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate735(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate736(.a(G504), .O(gate150inter7));
  inv1  gate737(.a(G507), .O(gate150inter8));
  nand2 gate738(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate739(.a(s_27), .b(gate150inter3), .O(gate150inter10));
  nor2  gate740(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate741(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate742(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate701(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate702(.a(gate151inter0), .b(s_22), .O(gate151inter1));
  and2  gate703(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate704(.a(s_22), .O(gate151inter3));
  inv1  gate705(.a(s_23), .O(gate151inter4));
  nand2 gate706(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate707(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate708(.a(G510), .O(gate151inter7));
  inv1  gate709(.a(G513), .O(gate151inter8));
  nand2 gate710(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate711(.a(s_23), .b(gate151inter3), .O(gate151inter10));
  nor2  gate712(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate713(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate714(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1527(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1528(.a(gate155inter0), .b(s_140), .O(gate155inter1));
  and2  gate1529(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1530(.a(s_140), .O(gate155inter3));
  inv1  gate1531(.a(s_141), .O(gate155inter4));
  nand2 gate1532(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1533(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1534(.a(G432), .O(gate155inter7));
  inv1  gate1535(.a(G525), .O(gate155inter8));
  nand2 gate1536(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1537(.a(s_141), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1538(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1539(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1540(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1345(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1346(.a(gate157inter0), .b(s_114), .O(gate157inter1));
  and2  gate1347(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1348(.a(s_114), .O(gate157inter3));
  inv1  gate1349(.a(s_115), .O(gate157inter4));
  nand2 gate1350(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1351(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1352(.a(G438), .O(gate157inter7));
  inv1  gate1353(.a(G528), .O(gate157inter8));
  nand2 gate1354(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1355(.a(s_115), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1356(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1357(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1358(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1947(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1948(.a(gate160inter0), .b(s_200), .O(gate160inter1));
  and2  gate1949(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1950(.a(s_200), .O(gate160inter3));
  inv1  gate1951(.a(s_201), .O(gate160inter4));
  nand2 gate1952(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1953(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1954(.a(G447), .O(gate160inter7));
  inv1  gate1955(.a(G531), .O(gate160inter8));
  nand2 gate1956(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1957(.a(s_201), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1958(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1959(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1960(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1653(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1654(.a(gate161inter0), .b(s_158), .O(gate161inter1));
  and2  gate1655(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1656(.a(s_158), .O(gate161inter3));
  inv1  gate1657(.a(s_159), .O(gate161inter4));
  nand2 gate1658(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1659(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1660(.a(G450), .O(gate161inter7));
  inv1  gate1661(.a(G534), .O(gate161inter8));
  nand2 gate1662(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1663(.a(s_159), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1664(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1665(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1666(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate869(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate870(.a(gate162inter0), .b(s_46), .O(gate162inter1));
  and2  gate871(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate872(.a(s_46), .O(gate162inter3));
  inv1  gate873(.a(s_47), .O(gate162inter4));
  nand2 gate874(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate875(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate876(.a(G453), .O(gate162inter7));
  inv1  gate877(.a(G534), .O(gate162inter8));
  nand2 gate878(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate879(.a(s_47), .b(gate162inter3), .O(gate162inter10));
  nor2  gate880(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate881(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate882(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate659(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate660(.a(gate168inter0), .b(s_16), .O(gate168inter1));
  and2  gate661(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate662(.a(s_16), .O(gate168inter3));
  inv1  gate663(.a(s_17), .O(gate168inter4));
  nand2 gate664(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate665(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate666(.a(G471), .O(gate168inter7));
  inv1  gate667(.a(G543), .O(gate168inter8));
  nand2 gate668(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate669(.a(s_17), .b(gate168inter3), .O(gate168inter10));
  nor2  gate670(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate671(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate672(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1709(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1710(.a(gate170inter0), .b(s_166), .O(gate170inter1));
  and2  gate1711(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1712(.a(s_166), .O(gate170inter3));
  inv1  gate1713(.a(s_167), .O(gate170inter4));
  nand2 gate1714(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1715(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1716(.a(G477), .O(gate170inter7));
  inv1  gate1717(.a(G546), .O(gate170inter8));
  nand2 gate1718(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1719(.a(s_167), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1720(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1721(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1722(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1051(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1052(.a(gate171inter0), .b(s_72), .O(gate171inter1));
  and2  gate1053(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1054(.a(s_72), .O(gate171inter3));
  inv1  gate1055(.a(s_73), .O(gate171inter4));
  nand2 gate1056(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1057(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1058(.a(G480), .O(gate171inter7));
  inv1  gate1059(.a(G549), .O(gate171inter8));
  nand2 gate1060(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1061(.a(s_73), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1062(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1063(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1064(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1905(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1906(.a(gate181inter0), .b(s_194), .O(gate181inter1));
  and2  gate1907(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1908(.a(s_194), .O(gate181inter3));
  inv1  gate1909(.a(s_195), .O(gate181inter4));
  nand2 gate1910(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1911(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1912(.a(G510), .O(gate181inter7));
  inv1  gate1913(.a(G564), .O(gate181inter8));
  nand2 gate1914(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1915(.a(s_195), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1916(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1917(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1918(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1401(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1402(.a(gate184inter0), .b(s_122), .O(gate184inter1));
  and2  gate1403(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1404(.a(s_122), .O(gate184inter3));
  inv1  gate1405(.a(s_123), .O(gate184inter4));
  nand2 gate1406(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1407(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1408(.a(G519), .O(gate184inter7));
  inv1  gate1409(.a(G567), .O(gate184inter8));
  nand2 gate1410(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1411(.a(s_123), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1412(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1413(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1414(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1163(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1164(.a(gate193inter0), .b(s_88), .O(gate193inter1));
  and2  gate1165(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1166(.a(s_88), .O(gate193inter3));
  inv1  gate1167(.a(s_89), .O(gate193inter4));
  nand2 gate1168(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1169(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1170(.a(G586), .O(gate193inter7));
  inv1  gate1171(.a(G587), .O(gate193inter8));
  nand2 gate1172(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1173(.a(s_89), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1174(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1175(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1176(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1443(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1444(.a(gate195inter0), .b(s_128), .O(gate195inter1));
  and2  gate1445(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1446(.a(s_128), .O(gate195inter3));
  inv1  gate1447(.a(s_129), .O(gate195inter4));
  nand2 gate1448(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1449(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1450(.a(G590), .O(gate195inter7));
  inv1  gate1451(.a(G591), .O(gate195inter8));
  nand2 gate1452(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1453(.a(s_129), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1454(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1455(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1456(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1191(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1192(.a(gate196inter0), .b(s_92), .O(gate196inter1));
  and2  gate1193(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1194(.a(s_92), .O(gate196inter3));
  inv1  gate1195(.a(s_93), .O(gate196inter4));
  nand2 gate1196(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1197(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1198(.a(G592), .O(gate196inter7));
  inv1  gate1199(.a(G593), .O(gate196inter8));
  nand2 gate1200(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1201(.a(s_93), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1202(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1203(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1204(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1177(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1178(.a(gate199inter0), .b(s_90), .O(gate199inter1));
  and2  gate1179(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1180(.a(s_90), .O(gate199inter3));
  inv1  gate1181(.a(s_91), .O(gate199inter4));
  nand2 gate1182(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1183(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1184(.a(G598), .O(gate199inter7));
  inv1  gate1185(.a(G599), .O(gate199inter8));
  nand2 gate1186(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1187(.a(s_91), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1188(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1189(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1190(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate743(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate744(.a(gate203inter0), .b(s_28), .O(gate203inter1));
  and2  gate745(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate746(.a(s_28), .O(gate203inter3));
  inv1  gate747(.a(s_29), .O(gate203inter4));
  nand2 gate748(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate749(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate750(.a(G602), .O(gate203inter7));
  inv1  gate751(.a(G612), .O(gate203inter8));
  nand2 gate752(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate753(.a(s_29), .b(gate203inter3), .O(gate203inter10));
  nor2  gate754(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate755(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate756(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1807(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1808(.a(gate208inter0), .b(s_180), .O(gate208inter1));
  and2  gate1809(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1810(.a(s_180), .O(gate208inter3));
  inv1  gate1811(.a(s_181), .O(gate208inter4));
  nand2 gate1812(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1813(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1814(.a(G627), .O(gate208inter7));
  inv1  gate1815(.a(G637), .O(gate208inter8));
  nand2 gate1816(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1817(.a(s_181), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1818(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1819(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1820(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1275(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1276(.a(gate210inter0), .b(s_104), .O(gate210inter1));
  and2  gate1277(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1278(.a(s_104), .O(gate210inter3));
  inv1  gate1279(.a(s_105), .O(gate210inter4));
  nand2 gate1280(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1281(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1282(.a(G607), .O(gate210inter7));
  inv1  gate1283(.a(G666), .O(gate210inter8));
  nand2 gate1284(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1285(.a(s_105), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1286(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1287(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1288(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1891(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1892(.a(gate213inter0), .b(s_192), .O(gate213inter1));
  and2  gate1893(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1894(.a(s_192), .O(gate213inter3));
  inv1  gate1895(.a(s_193), .O(gate213inter4));
  nand2 gate1896(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1897(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1898(.a(G602), .O(gate213inter7));
  inv1  gate1899(.a(G672), .O(gate213inter8));
  nand2 gate1900(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1901(.a(s_193), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1902(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1903(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1904(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1303(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1304(.a(gate216inter0), .b(s_108), .O(gate216inter1));
  and2  gate1305(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1306(.a(s_108), .O(gate216inter3));
  inv1  gate1307(.a(s_109), .O(gate216inter4));
  nand2 gate1308(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1309(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1310(.a(G617), .O(gate216inter7));
  inv1  gate1311(.a(G675), .O(gate216inter8));
  nand2 gate1312(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1313(.a(s_109), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1314(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1315(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1316(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1765(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1766(.a(gate221inter0), .b(s_174), .O(gate221inter1));
  and2  gate1767(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1768(.a(s_174), .O(gate221inter3));
  inv1  gate1769(.a(s_175), .O(gate221inter4));
  nand2 gate1770(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1771(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1772(.a(G622), .O(gate221inter7));
  inv1  gate1773(.a(G684), .O(gate221inter8));
  nand2 gate1774(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1775(.a(s_175), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1776(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1777(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1778(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1009(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1010(.a(gate226inter0), .b(s_66), .O(gate226inter1));
  and2  gate1011(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1012(.a(s_66), .O(gate226inter3));
  inv1  gate1013(.a(s_67), .O(gate226inter4));
  nand2 gate1014(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1015(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1016(.a(G692), .O(gate226inter7));
  inv1  gate1017(.a(G693), .O(gate226inter8));
  nand2 gate1018(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1019(.a(s_67), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1020(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1021(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1022(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate841(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate842(.a(gate230inter0), .b(s_42), .O(gate230inter1));
  and2  gate843(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate844(.a(s_42), .O(gate230inter3));
  inv1  gate845(.a(s_43), .O(gate230inter4));
  nand2 gate846(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate847(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate848(.a(G700), .O(gate230inter7));
  inv1  gate849(.a(G701), .O(gate230inter8));
  nand2 gate850(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate851(.a(s_43), .b(gate230inter3), .O(gate230inter10));
  nor2  gate852(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate853(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate854(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate757(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate758(.a(gate245inter0), .b(s_30), .O(gate245inter1));
  and2  gate759(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate760(.a(s_30), .O(gate245inter3));
  inv1  gate761(.a(s_31), .O(gate245inter4));
  nand2 gate762(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate763(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate764(.a(G248), .O(gate245inter7));
  inv1  gate765(.a(G736), .O(gate245inter8));
  nand2 gate766(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate767(.a(s_31), .b(gate245inter3), .O(gate245inter10));
  nor2  gate768(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate769(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate770(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1429(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1430(.a(gate253inter0), .b(s_126), .O(gate253inter1));
  and2  gate1431(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1432(.a(s_126), .O(gate253inter3));
  inv1  gate1433(.a(s_127), .O(gate253inter4));
  nand2 gate1434(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1435(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1436(.a(G260), .O(gate253inter7));
  inv1  gate1437(.a(G748), .O(gate253inter8));
  nand2 gate1438(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1439(.a(s_127), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1440(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1441(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1442(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1919(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1920(.a(gate254inter0), .b(s_196), .O(gate254inter1));
  and2  gate1921(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1922(.a(s_196), .O(gate254inter3));
  inv1  gate1923(.a(s_197), .O(gate254inter4));
  nand2 gate1924(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1925(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1926(.a(G712), .O(gate254inter7));
  inv1  gate1927(.a(G748), .O(gate254inter8));
  nand2 gate1928(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1929(.a(s_197), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1930(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1931(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1932(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1149(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1150(.a(gate260inter0), .b(s_86), .O(gate260inter1));
  and2  gate1151(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1152(.a(s_86), .O(gate260inter3));
  inv1  gate1153(.a(s_87), .O(gate260inter4));
  nand2 gate1154(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1155(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1156(.a(G760), .O(gate260inter7));
  inv1  gate1157(.a(G761), .O(gate260inter8));
  nand2 gate1158(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1159(.a(s_87), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1160(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1161(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1162(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1513(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1514(.a(gate263inter0), .b(s_138), .O(gate263inter1));
  and2  gate1515(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1516(.a(s_138), .O(gate263inter3));
  inv1  gate1517(.a(s_139), .O(gate263inter4));
  nand2 gate1518(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1519(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1520(.a(G766), .O(gate263inter7));
  inv1  gate1521(.a(G767), .O(gate263inter8));
  nand2 gate1522(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1523(.a(s_139), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1524(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1525(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1526(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1849(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1850(.a(gate270inter0), .b(s_186), .O(gate270inter1));
  and2  gate1851(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1852(.a(s_186), .O(gate270inter3));
  inv1  gate1853(.a(s_187), .O(gate270inter4));
  nand2 gate1854(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1855(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1856(.a(G657), .O(gate270inter7));
  inv1  gate1857(.a(G785), .O(gate270inter8));
  nand2 gate1858(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1859(.a(s_187), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1860(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1861(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1862(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate799(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate800(.a(gate272inter0), .b(s_36), .O(gate272inter1));
  and2  gate801(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate802(.a(s_36), .O(gate272inter3));
  inv1  gate803(.a(s_37), .O(gate272inter4));
  nand2 gate804(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate805(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate806(.a(G663), .O(gate272inter7));
  inv1  gate807(.a(G791), .O(gate272inter8));
  nand2 gate808(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate809(.a(s_37), .b(gate272inter3), .O(gate272inter10));
  nor2  gate810(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate811(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate812(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate995(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate996(.a(gate278inter0), .b(s_64), .O(gate278inter1));
  and2  gate997(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate998(.a(s_64), .O(gate278inter3));
  inv1  gate999(.a(s_65), .O(gate278inter4));
  nand2 gate1000(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1001(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1002(.a(G776), .O(gate278inter7));
  inv1  gate1003(.a(G800), .O(gate278inter8));
  nand2 gate1004(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1005(.a(s_65), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1006(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1007(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1008(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1289(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1290(.a(gate287inter0), .b(s_106), .O(gate287inter1));
  and2  gate1291(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1292(.a(s_106), .O(gate287inter3));
  inv1  gate1293(.a(s_107), .O(gate287inter4));
  nand2 gate1294(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1295(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1296(.a(G663), .O(gate287inter7));
  inv1  gate1297(.a(G815), .O(gate287inter8));
  nand2 gate1298(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1299(.a(s_107), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1300(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1301(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1302(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate953(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate954(.a(gate292inter0), .b(s_58), .O(gate292inter1));
  and2  gate955(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate956(.a(s_58), .O(gate292inter3));
  inv1  gate957(.a(s_59), .O(gate292inter4));
  nand2 gate958(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate959(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate960(.a(G824), .O(gate292inter7));
  inv1  gate961(.a(G825), .O(gate292inter8));
  nand2 gate962(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate963(.a(s_59), .b(gate292inter3), .O(gate292inter10));
  nor2  gate964(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate965(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate966(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate925(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate926(.a(gate294inter0), .b(s_54), .O(gate294inter1));
  and2  gate927(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate928(.a(s_54), .O(gate294inter3));
  inv1  gate929(.a(s_55), .O(gate294inter4));
  nand2 gate930(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate931(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate932(.a(G832), .O(gate294inter7));
  inv1  gate933(.a(G833), .O(gate294inter8));
  nand2 gate934(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate935(.a(s_55), .b(gate294inter3), .O(gate294inter10));
  nor2  gate936(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate937(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate938(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate785(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate786(.a(gate398inter0), .b(s_34), .O(gate398inter1));
  and2  gate787(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate788(.a(s_34), .O(gate398inter3));
  inv1  gate789(.a(s_35), .O(gate398inter4));
  nand2 gate790(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate791(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate792(.a(G12), .O(gate398inter7));
  inv1  gate793(.a(G1069), .O(gate398inter8));
  nand2 gate794(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate795(.a(s_35), .b(gate398inter3), .O(gate398inter10));
  nor2  gate796(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate797(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate798(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1261(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1262(.a(gate403inter0), .b(s_102), .O(gate403inter1));
  and2  gate1263(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1264(.a(s_102), .O(gate403inter3));
  inv1  gate1265(.a(s_103), .O(gate403inter4));
  nand2 gate1266(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1267(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1268(.a(G17), .O(gate403inter7));
  inv1  gate1269(.a(G1084), .O(gate403inter8));
  nand2 gate1270(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1271(.a(s_103), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1272(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1273(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1274(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1933(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1934(.a(gate409inter0), .b(s_198), .O(gate409inter1));
  and2  gate1935(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1936(.a(s_198), .O(gate409inter3));
  inv1  gate1937(.a(s_199), .O(gate409inter4));
  nand2 gate1938(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1939(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1940(.a(G23), .O(gate409inter7));
  inv1  gate1941(.a(G1102), .O(gate409inter8));
  nand2 gate1942(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1943(.a(s_199), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1944(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1945(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1946(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1037(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1038(.a(gate410inter0), .b(s_70), .O(gate410inter1));
  and2  gate1039(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1040(.a(s_70), .O(gate410inter3));
  inv1  gate1041(.a(s_71), .O(gate410inter4));
  nand2 gate1042(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1043(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1044(.a(G24), .O(gate410inter7));
  inv1  gate1045(.a(G1105), .O(gate410inter8));
  nand2 gate1046(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1047(.a(s_71), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1048(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1049(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1050(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1541(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1542(.a(gate411inter0), .b(s_142), .O(gate411inter1));
  and2  gate1543(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1544(.a(s_142), .O(gate411inter3));
  inv1  gate1545(.a(s_143), .O(gate411inter4));
  nand2 gate1546(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1547(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1548(.a(G25), .O(gate411inter7));
  inv1  gate1549(.a(G1108), .O(gate411inter8));
  nand2 gate1550(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1551(.a(s_143), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1552(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1553(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1554(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate645(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate646(.a(gate417inter0), .b(s_14), .O(gate417inter1));
  and2  gate647(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate648(.a(s_14), .O(gate417inter3));
  inv1  gate649(.a(s_15), .O(gate417inter4));
  nand2 gate650(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate651(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate652(.a(G31), .O(gate417inter7));
  inv1  gate653(.a(G1126), .O(gate417inter8));
  nand2 gate654(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate655(.a(s_15), .b(gate417inter3), .O(gate417inter10));
  nor2  gate656(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate657(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate658(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate589(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate590(.a(gate420inter0), .b(s_6), .O(gate420inter1));
  and2  gate591(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate592(.a(s_6), .O(gate420inter3));
  inv1  gate593(.a(s_7), .O(gate420inter4));
  nand2 gate594(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate595(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate596(.a(G1036), .O(gate420inter7));
  inv1  gate597(.a(G1132), .O(gate420inter8));
  nand2 gate598(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate599(.a(s_7), .b(gate420inter3), .O(gate420inter10));
  nor2  gate600(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate601(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate602(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate911(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate912(.a(gate424inter0), .b(s_52), .O(gate424inter1));
  and2  gate913(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate914(.a(s_52), .O(gate424inter3));
  inv1  gate915(.a(s_53), .O(gate424inter4));
  nand2 gate916(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate917(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate918(.a(G1042), .O(gate424inter7));
  inv1  gate919(.a(G1138), .O(gate424inter8));
  nand2 gate920(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate921(.a(s_53), .b(gate424inter3), .O(gate424inter10));
  nor2  gate922(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate923(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate924(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate771(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate772(.a(gate428inter0), .b(s_32), .O(gate428inter1));
  and2  gate773(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate774(.a(s_32), .O(gate428inter3));
  inv1  gate775(.a(s_33), .O(gate428inter4));
  nand2 gate776(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate777(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate778(.a(G1048), .O(gate428inter7));
  inv1  gate779(.a(G1144), .O(gate428inter8));
  nand2 gate780(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate781(.a(s_33), .b(gate428inter3), .O(gate428inter10));
  nor2  gate782(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate783(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate784(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1863(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1864(.a(gate429inter0), .b(s_188), .O(gate429inter1));
  and2  gate1865(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1866(.a(s_188), .O(gate429inter3));
  inv1  gate1867(.a(s_189), .O(gate429inter4));
  nand2 gate1868(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1869(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1870(.a(G6), .O(gate429inter7));
  inv1  gate1871(.a(G1147), .O(gate429inter8));
  nand2 gate1872(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1873(.a(s_189), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1874(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1875(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1876(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1877(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1878(.a(gate433inter0), .b(s_190), .O(gate433inter1));
  and2  gate1879(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1880(.a(s_190), .O(gate433inter3));
  inv1  gate1881(.a(s_191), .O(gate433inter4));
  nand2 gate1882(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1883(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1884(.a(G8), .O(gate433inter7));
  inv1  gate1885(.a(G1153), .O(gate433inter8));
  nand2 gate1886(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1887(.a(s_191), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1888(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1889(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1890(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate603(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate604(.a(gate434inter0), .b(s_8), .O(gate434inter1));
  and2  gate605(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate606(.a(s_8), .O(gate434inter3));
  inv1  gate607(.a(s_9), .O(gate434inter4));
  nand2 gate608(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate609(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate610(.a(G1057), .O(gate434inter7));
  inv1  gate611(.a(G1153), .O(gate434inter8));
  nand2 gate612(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate613(.a(s_9), .b(gate434inter3), .O(gate434inter10));
  nor2  gate614(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate615(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate616(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1247(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1248(.a(gate445inter0), .b(s_100), .O(gate445inter1));
  and2  gate1249(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1250(.a(s_100), .O(gate445inter3));
  inv1  gate1251(.a(s_101), .O(gate445inter4));
  nand2 gate1252(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1253(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1254(.a(G14), .O(gate445inter7));
  inv1  gate1255(.a(G1171), .O(gate445inter8));
  nand2 gate1256(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1257(.a(s_101), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1258(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1259(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1260(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate967(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate968(.a(gate446inter0), .b(s_60), .O(gate446inter1));
  and2  gate969(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate970(.a(s_60), .O(gate446inter3));
  inv1  gate971(.a(s_61), .O(gate446inter4));
  nand2 gate972(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate973(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate974(.a(G1075), .O(gate446inter7));
  inv1  gate975(.a(G1171), .O(gate446inter8));
  nand2 gate976(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate977(.a(s_61), .b(gate446inter3), .O(gate446inter10));
  nor2  gate978(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate979(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate980(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1093(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1094(.a(gate450inter0), .b(s_78), .O(gate450inter1));
  and2  gate1095(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1096(.a(s_78), .O(gate450inter3));
  inv1  gate1097(.a(s_79), .O(gate450inter4));
  nand2 gate1098(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1099(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1100(.a(G1081), .O(gate450inter7));
  inv1  gate1101(.a(G1177), .O(gate450inter8));
  nand2 gate1102(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1103(.a(s_79), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1104(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1105(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1106(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1331(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1332(.a(gate457inter0), .b(s_112), .O(gate457inter1));
  and2  gate1333(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1334(.a(s_112), .O(gate457inter3));
  inv1  gate1335(.a(s_113), .O(gate457inter4));
  nand2 gate1336(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1337(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1338(.a(G20), .O(gate457inter7));
  inv1  gate1339(.a(G1189), .O(gate457inter8));
  nand2 gate1340(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1341(.a(s_113), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1342(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1343(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1344(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1135(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1136(.a(gate458inter0), .b(s_84), .O(gate458inter1));
  and2  gate1137(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1138(.a(s_84), .O(gate458inter3));
  inv1  gate1139(.a(s_85), .O(gate458inter4));
  nand2 gate1140(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1141(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1142(.a(G1093), .O(gate458inter7));
  inv1  gate1143(.a(G1189), .O(gate458inter8));
  nand2 gate1144(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1145(.a(s_85), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1146(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1147(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1148(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate561(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate562(.a(gate460inter0), .b(s_2), .O(gate460inter1));
  and2  gate563(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate564(.a(s_2), .O(gate460inter3));
  inv1  gate565(.a(s_3), .O(gate460inter4));
  nand2 gate566(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate567(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate568(.a(G1096), .O(gate460inter7));
  inv1  gate569(.a(G1192), .O(gate460inter8));
  nand2 gate570(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate571(.a(s_3), .b(gate460inter3), .O(gate460inter10));
  nor2  gate572(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate573(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate574(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1485(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1486(.a(gate463inter0), .b(s_134), .O(gate463inter1));
  and2  gate1487(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1488(.a(s_134), .O(gate463inter3));
  inv1  gate1489(.a(s_135), .O(gate463inter4));
  nand2 gate1490(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1491(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1492(.a(G23), .O(gate463inter7));
  inv1  gate1493(.a(G1198), .O(gate463inter8));
  nand2 gate1494(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1495(.a(s_135), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1496(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1497(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1498(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1639(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1640(.a(gate464inter0), .b(s_156), .O(gate464inter1));
  and2  gate1641(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1642(.a(s_156), .O(gate464inter3));
  inv1  gate1643(.a(s_157), .O(gate464inter4));
  nand2 gate1644(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1645(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1646(.a(G1102), .O(gate464inter7));
  inv1  gate1647(.a(G1198), .O(gate464inter8));
  nand2 gate1648(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1649(.a(s_157), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1650(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1651(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1652(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1023(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1024(.a(gate466inter0), .b(s_68), .O(gate466inter1));
  and2  gate1025(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1026(.a(s_68), .O(gate466inter3));
  inv1  gate1027(.a(s_69), .O(gate466inter4));
  nand2 gate1028(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1029(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1030(.a(G1105), .O(gate466inter7));
  inv1  gate1031(.a(G1201), .O(gate466inter8));
  nand2 gate1032(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1033(.a(s_69), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1034(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1035(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1036(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate813(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate814(.a(gate473inter0), .b(s_38), .O(gate473inter1));
  and2  gate815(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate816(.a(s_38), .O(gate473inter3));
  inv1  gate817(.a(s_39), .O(gate473inter4));
  nand2 gate818(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate819(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate820(.a(G28), .O(gate473inter7));
  inv1  gate821(.a(G1213), .O(gate473inter8));
  nand2 gate822(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate823(.a(s_39), .b(gate473inter3), .O(gate473inter10));
  nor2  gate824(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate825(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate826(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1555(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1556(.a(gate476inter0), .b(s_144), .O(gate476inter1));
  and2  gate1557(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1558(.a(s_144), .O(gate476inter3));
  inv1  gate1559(.a(s_145), .O(gate476inter4));
  nand2 gate1560(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1561(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1562(.a(G1120), .O(gate476inter7));
  inv1  gate1563(.a(G1216), .O(gate476inter8));
  nand2 gate1564(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1565(.a(s_145), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1566(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1567(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1568(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1317(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1318(.a(gate479inter0), .b(s_110), .O(gate479inter1));
  and2  gate1319(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1320(.a(s_110), .O(gate479inter3));
  inv1  gate1321(.a(s_111), .O(gate479inter4));
  nand2 gate1322(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1323(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1324(.a(G31), .O(gate479inter7));
  inv1  gate1325(.a(G1222), .O(gate479inter8));
  nand2 gate1326(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1327(.a(s_111), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1328(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1329(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1330(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate687(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate688(.a(gate486inter0), .b(s_20), .O(gate486inter1));
  and2  gate689(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate690(.a(s_20), .O(gate486inter3));
  inv1  gate691(.a(s_21), .O(gate486inter4));
  nand2 gate692(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate693(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate694(.a(G1234), .O(gate486inter7));
  inv1  gate695(.a(G1235), .O(gate486inter8));
  nand2 gate696(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate697(.a(s_21), .b(gate486inter3), .O(gate486inter10));
  nor2  gate698(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate699(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate700(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1751(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1752(.a(gate488inter0), .b(s_172), .O(gate488inter1));
  and2  gate1753(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1754(.a(s_172), .O(gate488inter3));
  inv1  gate1755(.a(s_173), .O(gate488inter4));
  nand2 gate1756(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1757(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1758(.a(G1238), .O(gate488inter7));
  inv1  gate1759(.a(G1239), .O(gate488inter8));
  nand2 gate1760(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1761(.a(s_173), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1762(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1763(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1764(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate715(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate716(.a(gate489inter0), .b(s_24), .O(gate489inter1));
  and2  gate717(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate718(.a(s_24), .O(gate489inter3));
  inv1  gate719(.a(s_25), .O(gate489inter4));
  nand2 gate720(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate721(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate722(.a(G1240), .O(gate489inter7));
  inv1  gate723(.a(G1241), .O(gate489inter8));
  nand2 gate724(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate725(.a(s_25), .b(gate489inter3), .O(gate489inter10));
  nor2  gate726(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate727(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate728(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1667(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1668(.a(gate490inter0), .b(s_160), .O(gate490inter1));
  and2  gate1669(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1670(.a(s_160), .O(gate490inter3));
  inv1  gate1671(.a(s_161), .O(gate490inter4));
  nand2 gate1672(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1673(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1674(.a(G1242), .O(gate490inter7));
  inv1  gate1675(.a(G1243), .O(gate490inter8));
  nand2 gate1676(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1677(.a(s_161), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1678(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1679(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1680(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1681(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1682(.a(gate504inter0), .b(s_162), .O(gate504inter1));
  and2  gate1683(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1684(.a(s_162), .O(gate504inter3));
  inv1  gate1685(.a(s_163), .O(gate504inter4));
  nand2 gate1686(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1687(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1688(.a(G1270), .O(gate504inter7));
  inv1  gate1689(.a(G1271), .O(gate504inter8));
  nand2 gate1690(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1691(.a(s_163), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1692(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1693(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1694(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1695(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1696(.a(gate508inter0), .b(s_164), .O(gate508inter1));
  and2  gate1697(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1698(.a(s_164), .O(gate508inter3));
  inv1  gate1699(.a(s_165), .O(gate508inter4));
  nand2 gate1700(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1701(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1702(.a(G1278), .O(gate508inter7));
  inv1  gate1703(.a(G1279), .O(gate508inter8));
  nand2 gate1704(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1705(.a(s_165), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1706(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1707(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1708(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1205(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1206(.a(gate514inter0), .b(s_94), .O(gate514inter1));
  and2  gate1207(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1208(.a(s_94), .O(gate514inter3));
  inv1  gate1209(.a(s_95), .O(gate514inter4));
  nand2 gate1210(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1211(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1212(.a(G1290), .O(gate514inter7));
  inv1  gate1213(.a(G1291), .O(gate514inter8));
  nand2 gate1214(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1215(.a(s_95), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1216(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1217(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1218(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule