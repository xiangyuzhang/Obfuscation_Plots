module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate7inter0, gate7inter1, gate7inter2, gate7inter3, gate7inter4, gate7inter5, gate7inter6, gate7inter7, gate7inter8, gate7inter9, gate7inter10, gate7inter11, gate7inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );

  xor2  gate1197(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate1198(.a(gate2inter0), .b(s_142), .O(gate2inter1));
  and2  gate1199(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate1200(.a(s_142), .O(gate2inter3));
  inv1  gate1201(.a(s_143), .O(gate2inter4));
  nand2 gate1202(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate1203(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate1204(.a(N9), .O(gate2inter7));
  inv1  gate1205(.a(N13), .O(gate2inter8));
  nand2 gate1206(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate1207(.a(s_143), .b(gate2inter3), .O(gate2inter10));
  nor2  gate1208(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate1209(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate1210(.a(gate2inter12), .b(gate2inter1), .O(N251));

  xor2  gate1141(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate1142(.a(gate3inter0), .b(s_134), .O(gate3inter1));
  and2  gate1143(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate1144(.a(s_134), .O(gate3inter3));
  inv1  gate1145(.a(s_135), .O(gate3inter4));
  nand2 gate1146(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate1147(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate1148(.a(N17), .O(gate3inter7));
  inv1  gate1149(.a(N21), .O(gate3inter8));
  nand2 gate1150(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate1151(.a(s_135), .b(gate3inter3), .O(gate3inter10));
  nor2  gate1152(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate1153(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate1154(.a(gate3inter12), .b(gate3inter1), .O(N252));

  xor2  gate1393(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate1394(.a(gate4inter0), .b(s_170), .O(gate4inter1));
  and2  gate1395(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate1396(.a(s_170), .O(gate4inter3));
  inv1  gate1397(.a(s_171), .O(gate4inter4));
  nand2 gate1398(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate1399(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate1400(.a(N25), .O(gate4inter7));
  inv1  gate1401(.a(N29), .O(gate4inter8));
  nand2 gate1402(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate1403(.a(s_171), .b(gate4inter3), .O(gate4inter10));
  nor2  gate1404(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate1405(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate1406(.a(gate4inter12), .b(gate4inter1), .O(N253));

  xor2  gate945(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate946(.a(gate5inter0), .b(s_106), .O(gate5inter1));
  and2  gate947(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate948(.a(s_106), .O(gate5inter3));
  inv1  gate949(.a(s_107), .O(gate5inter4));
  nand2 gate950(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate951(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate952(.a(N33), .O(gate5inter7));
  inv1  gate953(.a(N37), .O(gate5inter8));
  nand2 gate954(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate955(.a(s_107), .b(gate5inter3), .O(gate5inter10));
  nor2  gate956(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate957(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate958(.a(gate5inter12), .b(gate5inter1), .O(N254));

  xor2  gate805(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate806(.a(gate6inter0), .b(s_86), .O(gate6inter1));
  and2  gate807(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate808(.a(s_86), .O(gate6inter3));
  inv1  gate809(.a(s_87), .O(gate6inter4));
  nand2 gate810(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate811(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate812(.a(N41), .O(gate6inter7));
  inv1  gate813(.a(N45), .O(gate6inter8));
  nand2 gate814(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate815(.a(s_87), .b(gate6inter3), .O(gate6inter10));
  nor2  gate816(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate817(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate818(.a(gate6inter12), .b(gate6inter1), .O(N255));

  xor2  gate721(.a(N53), .b(N49), .O(gate7inter0));
  nand2 gate722(.a(gate7inter0), .b(s_74), .O(gate7inter1));
  and2  gate723(.a(N53), .b(N49), .O(gate7inter2));
  inv1  gate724(.a(s_74), .O(gate7inter3));
  inv1  gate725(.a(s_75), .O(gate7inter4));
  nand2 gate726(.a(gate7inter4), .b(gate7inter3), .O(gate7inter5));
  nor2  gate727(.a(gate7inter5), .b(gate7inter2), .O(gate7inter6));
  inv1  gate728(.a(N49), .O(gate7inter7));
  inv1  gate729(.a(N53), .O(gate7inter8));
  nand2 gate730(.a(gate7inter8), .b(gate7inter7), .O(gate7inter9));
  nand2 gate731(.a(s_75), .b(gate7inter3), .O(gate7inter10));
  nor2  gate732(.a(gate7inter10), .b(gate7inter9), .O(gate7inter11));
  nor2  gate733(.a(gate7inter11), .b(gate7inter6), .O(gate7inter12));
  nand2 gate734(.a(gate7inter12), .b(gate7inter1), .O(N256));

  xor2  gate1379(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate1380(.a(gate8inter0), .b(s_168), .O(gate8inter1));
  and2  gate1381(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate1382(.a(s_168), .O(gate8inter3));
  inv1  gate1383(.a(s_169), .O(gate8inter4));
  nand2 gate1384(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate1385(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate1386(.a(N57), .O(gate8inter7));
  inv1  gate1387(.a(N61), .O(gate8inter8));
  nand2 gate1388(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate1389(.a(s_169), .b(gate8inter3), .O(gate8inter10));
  nor2  gate1390(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate1391(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate1392(.a(gate8inter12), .b(gate8inter1), .O(N257));

  xor2  gate1253(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate1254(.a(gate9inter0), .b(s_150), .O(gate9inter1));
  and2  gate1255(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate1256(.a(s_150), .O(gate9inter3));
  inv1  gate1257(.a(s_151), .O(gate9inter4));
  nand2 gate1258(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1259(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1260(.a(N65), .O(gate9inter7));
  inv1  gate1261(.a(N69), .O(gate9inter8));
  nand2 gate1262(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1263(.a(s_151), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1264(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1265(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1266(.a(gate9inter12), .b(gate9inter1), .O(N258));

  xor2  gate819(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate820(.a(gate10inter0), .b(s_88), .O(gate10inter1));
  and2  gate821(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate822(.a(s_88), .O(gate10inter3));
  inv1  gate823(.a(s_89), .O(gate10inter4));
  nand2 gate824(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate825(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate826(.a(N73), .O(gate10inter7));
  inv1  gate827(.a(N77), .O(gate10inter8));
  nand2 gate828(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate829(.a(s_89), .b(gate10inter3), .O(gate10inter10));
  nor2  gate830(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate831(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate832(.a(gate10inter12), .b(gate10inter1), .O(N259));

  xor2  gate735(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate736(.a(gate11inter0), .b(s_76), .O(gate11inter1));
  and2  gate737(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate738(.a(s_76), .O(gate11inter3));
  inv1  gate739(.a(s_77), .O(gate11inter4));
  nand2 gate740(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate741(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate742(.a(N81), .O(gate11inter7));
  inv1  gate743(.a(N85), .O(gate11inter8));
  nand2 gate744(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate745(.a(s_77), .b(gate11inter3), .O(gate11inter10));
  nor2  gate746(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate747(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate748(.a(gate11inter12), .b(gate11inter1), .O(N260));

  xor2  gate931(.a(N93), .b(N89), .O(gate12inter0));
  nand2 gate932(.a(gate12inter0), .b(s_104), .O(gate12inter1));
  and2  gate933(.a(N93), .b(N89), .O(gate12inter2));
  inv1  gate934(.a(s_104), .O(gate12inter3));
  inv1  gate935(.a(s_105), .O(gate12inter4));
  nand2 gate936(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate937(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate938(.a(N89), .O(gate12inter7));
  inv1  gate939(.a(N93), .O(gate12inter8));
  nand2 gate940(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate941(.a(s_105), .b(gate12inter3), .O(gate12inter10));
  nor2  gate942(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate943(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate944(.a(gate12inter12), .b(gate12inter1), .O(N261));

  xor2  gate483(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate484(.a(gate13inter0), .b(s_40), .O(gate13inter1));
  and2  gate485(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate486(.a(s_40), .O(gate13inter3));
  inv1  gate487(.a(s_41), .O(gate13inter4));
  nand2 gate488(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate489(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate490(.a(N97), .O(gate13inter7));
  inv1  gate491(.a(N101), .O(gate13inter8));
  nand2 gate492(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate493(.a(s_41), .b(gate13inter3), .O(gate13inter10));
  nor2  gate494(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate495(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate496(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );

  xor2  gate1421(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate1422(.a(gate15inter0), .b(s_174), .O(gate15inter1));
  and2  gate1423(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate1424(.a(s_174), .O(gate15inter3));
  inv1  gate1425(.a(s_175), .O(gate15inter4));
  nand2 gate1426(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1427(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1428(.a(N113), .O(gate15inter7));
  inv1  gate1429(.a(N117), .O(gate15inter8));
  nand2 gate1430(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1431(.a(s_175), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1432(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1433(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1434(.a(gate15inter12), .b(gate15inter1), .O(N264));

  xor2  gate665(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate666(.a(gate16inter0), .b(s_66), .O(gate16inter1));
  and2  gate667(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate668(.a(s_66), .O(gate16inter3));
  inv1  gate669(.a(s_67), .O(gate16inter4));
  nand2 gate670(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate671(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate672(.a(N121), .O(gate16inter7));
  inv1  gate673(.a(N125), .O(gate16inter8));
  nand2 gate674(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate675(.a(s_67), .b(gate16inter3), .O(gate16inter10));
  nor2  gate676(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate677(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate678(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate441(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate442(.a(gate25inter0), .b(s_34), .O(gate25inter1));
  and2  gate443(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate444(.a(s_34), .O(gate25inter3));
  inv1  gate445(.a(s_35), .O(gate25inter4));
  nand2 gate446(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate447(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate448(.a(N1), .O(gate25inter7));
  inv1  gate449(.a(N17), .O(gate25inter8));
  nand2 gate450(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate451(.a(s_35), .b(gate25inter3), .O(gate25inter10));
  nor2  gate452(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate453(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate454(.a(gate25inter12), .b(gate25inter1), .O(N274));

  xor2  gate399(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate400(.a(gate26inter0), .b(s_28), .O(gate26inter1));
  and2  gate401(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate402(.a(s_28), .O(gate26inter3));
  inv1  gate403(.a(s_29), .O(gate26inter4));
  nand2 gate404(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate405(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate406(.a(N33), .O(gate26inter7));
  inv1  gate407(.a(N49), .O(gate26inter8));
  nand2 gate408(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate409(.a(s_29), .b(gate26inter3), .O(gate26inter10));
  nor2  gate410(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate411(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate412(.a(gate26inter12), .b(gate26inter1), .O(N275));

  xor2  gate1169(.a(N21), .b(N5), .O(gate27inter0));
  nand2 gate1170(.a(gate27inter0), .b(s_138), .O(gate27inter1));
  and2  gate1171(.a(N21), .b(N5), .O(gate27inter2));
  inv1  gate1172(.a(s_138), .O(gate27inter3));
  inv1  gate1173(.a(s_139), .O(gate27inter4));
  nand2 gate1174(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1175(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1176(.a(N5), .O(gate27inter7));
  inv1  gate1177(.a(N21), .O(gate27inter8));
  nand2 gate1178(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1179(.a(s_139), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1180(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1181(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1182(.a(gate27inter12), .b(gate27inter1), .O(N276));

  xor2  gate791(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate792(.a(gate28inter0), .b(s_84), .O(gate28inter1));
  and2  gate793(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate794(.a(s_84), .O(gate28inter3));
  inv1  gate795(.a(s_85), .O(gate28inter4));
  nand2 gate796(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate797(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate798(.a(N37), .O(gate28inter7));
  inv1  gate799(.a(N53), .O(gate28inter8));
  nand2 gate800(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate801(.a(s_85), .b(gate28inter3), .O(gate28inter10));
  nor2  gate802(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate803(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate804(.a(gate28inter12), .b(gate28inter1), .O(N277));

  xor2  gate763(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate764(.a(gate29inter0), .b(s_80), .O(gate29inter1));
  and2  gate765(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate766(.a(s_80), .O(gate29inter3));
  inv1  gate767(.a(s_81), .O(gate29inter4));
  nand2 gate768(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate769(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate770(.a(N9), .O(gate29inter7));
  inv1  gate771(.a(N25), .O(gate29inter8));
  nand2 gate772(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate773(.a(s_81), .b(gate29inter3), .O(gate29inter10));
  nor2  gate774(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate775(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate776(.a(gate29inter12), .b(gate29inter1), .O(N278));

  xor2  gate987(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate988(.a(gate30inter0), .b(s_112), .O(gate30inter1));
  and2  gate989(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate990(.a(s_112), .O(gate30inter3));
  inv1  gate991(.a(s_113), .O(gate30inter4));
  nand2 gate992(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate993(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate994(.a(N41), .O(gate30inter7));
  inv1  gate995(.a(N57), .O(gate30inter8));
  nand2 gate996(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate997(.a(s_113), .b(gate30inter3), .O(gate30inter10));
  nor2  gate998(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate999(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1000(.a(gate30inter12), .b(gate30inter1), .O(N279));

  xor2  gate539(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate540(.a(gate31inter0), .b(s_48), .O(gate31inter1));
  and2  gate541(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate542(.a(s_48), .O(gate31inter3));
  inv1  gate543(.a(s_49), .O(gate31inter4));
  nand2 gate544(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate545(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate546(.a(N13), .O(gate31inter7));
  inv1  gate547(.a(N29), .O(gate31inter8));
  nand2 gate548(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate549(.a(s_49), .b(gate31inter3), .O(gate31inter10));
  nor2  gate550(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate551(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate552(.a(gate31inter12), .b(gate31inter1), .O(N280));

  xor2  gate245(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate246(.a(gate32inter0), .b(s_6), .O(gate32inter1));
  and2  gate247(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate248(.a(s_6), .O(gate32inter3));
  inv1  gate249(.a(s_7), .O(gate32inter4));
  nand2 gate250(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate251(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate252(.a(N45), .O(gate32inter7));
  inv1  gate253(.a(N61), .O(gate32inter8));
  nand2 gate254(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate255(.a(s_7), .b(gate32inter3), .O(gate32inter10));
  nor2  gate256(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate257(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate258(.a(gate32inter12), .b(gate32inter1), .O(N281));

  xor2  gate511(.a(N81), .b(N65), .O(gate33inter0));
  nand2 gate512(.a(gate33inter0), .b(s_44), .O(gate33inter1));
  and2  gate513(.a(N81), .b(N65), .O(gate33inter2));
  inv1  gate514(.a(s_44), .O(gate33inter3));
  inv1  gate515(.a(s_45), .O(gate33inter4));
  nand2 gate516(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate517(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate518(.a(N65), .O(gate33inter7));
  inv1  gate519(.a(N81), .O(gate33inter8));
  nand2 gate520(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate521(.a(s_45), .b(gate33inter3), .O(gate33inter10));
  nor2  gate522(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate523(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate524(.a(gate33inter12), .b(gate33inter1), .O(N282));

  xor2  gate1029(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate1030(.a(gate34inter0), .b(s_118), .O(gate34inter1));
  and2  gate1031(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate1032(.a(s_118), .O(gate34inter3));
  inv1  gate1033(.a(s_119), .O(gate34inter4));
  nand2 gate1034(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1035(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1036(.a(N97), .O(gate34inter7));
  inv1  gate1037(.a(N113), .O(gate34inter8));
  nand2 gate1038(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1039(.a(s_119), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1040(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1041(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1042(.a(gate34inter12), .b(gate34inter1), .O(N283));

  xor2  gate1071(.a(N85), .b(N69), .O(gate35inter0));
  nand2 gate1072(.a(gate35inter0), .b(s_124), .O(gate35inter1));
  and2  gate1073(.a(N85), .b(N69), .O(gate35inter2));
  inv1  gate1074(.a(s_124), .O(gate35inter3));
  inv1  gate1075(.a(s_125), .O(gate35inter4));
  nand2 gate1076(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1077(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1078(.a(N69), .O(gate35inter7));
  inv1  gate1079(.a(N85), .O(gate35inter8));
  nand2 gate1080(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1081(.a(s_125), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1082(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1083(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1084(.a(gate35inter12), .b(gate35inter1), .O(N284));

  xor2  gate371(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate372(.a(gate36inter0), .b(s_24), .O(gate36inter1));
  and2  gate373(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate374(.a(s_24), .O(gate36inter3));
  inv1  gate375(.a(s_25), .O(gate36inter4));
  nand2 gate376(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate377(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate378(.a(N101), .O(gate36inter7));
  inv1  gate379(.a(N117), .O(gate36inter8));
  nand2 gate380(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate381(.a(s_25), .b(gate36inter3), .O(gate36inter10));
  nor2  gate382(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate383(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate384(.a(gate36inter12), .b(gate36inter1), .O(N285));

  xor2  gate1225(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate1226(.a(gate37inter0), .b(s_146), .O(gate37inter1));
  and2  gate1227(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate1228(.a(s_146), .O(gate37inter3));
  inv1  gate1229(.a(s_147), .O(gate37inter4));
  nand2 gate1230(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1231(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1232(.a(N73), .O(gate37inter7));
  inv1  gate1233(.a(N89), .O(gate37inter8));
  nand2 gate1234(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1235(.a(s_147), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1236(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1237(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1238(.a(gate37inter12), .b(gate37inter1), .O(N286));

  xor2  gate343(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate344(.a(gate38inter0), .b(s_20), .O(gate38inter1));
  and2  gate345(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate346(.a(s_20), .O(gate38inter3));
  inv1  gate347(.a(s_21), .O(gate38inter4));
  nand2 gate348(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate349(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate350(.a(N105), .O(gate38inter7));
  inv1  gate351(.a(N121), .O(gate38inter8));
  nand2 gate352(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate353(.a(s_21), .b(gate38inter3), .O(gate38inter10));
  nor2  gate354(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate355(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate356(.a(gate38inter12), .b(gate38inter1), .O(N287));
xor2 gate39( .a(N77), .b(N93), .O(N288) );

  xor2  gate1435(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate1436(.a(gate40inter0), .b(s_176), .O(gate40inter1));
  and2  gate1437(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate1438(.a(s_176), .O(gate40inter3));
  inv1  gate1439(.a(s_177), .O(gate40inter4));
  nand2 gate1440(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1441(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1442(.a(N109), .O(gate40inter7));
  inv1  gate1443(.a(N125), .O(gate40inter8));
  nand2 gate1444(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1445(.a(s_177), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1446(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1447(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1448(.a(gate40inter12), .b(gate40inter1), .O(N289));

  xor2  gate1001(.a(N251), .b(N250), .O(gate41inter0));
  nand2 gate1002(.a(gate41inter0), .b(s_114), .O(gate41inter1));
  and2  gate1003(.a(N251), .b(N250), .O(gate41inter2));
  inv1  gate1004(.a(s_114), .O(gate41inter3));
  inv1  gate1005(.a(s_115), .O(gate41inter4));
  nand2 gate1006(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1007(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1008(.a(N250), .O(gate41inter7));
  inv1  gate1009(.a(N251), .O(gate41inter8));
  nand2 gate1010(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1011(.a(s_115), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1012(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1013(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1014(.a(gate41inter12), .b(gate41inter1), .O(N290));

  xor2  gate259(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate260(.a(gate42inter0), .b(s_8), .O(gate42inter1));
  and2  gate261(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate262(.a(s_8), .O(gate42inter3));
  inv1  gate263(.a(s_9), .O(gate42inter4));
  nand2 gate264(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate265(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate266(.a(N252), .O(gate42inter7));
  inv1  gate267(.a(N253), .O(gate42inter8));
  nand2 gate268(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate269(.a(s_9), .b(gate42inter3), .O(gate42inter10));
  nor2  gate270(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate271(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate272(.a(gate42inter12), .b(gate42inter1), .O(N293));

  xor2  gate749(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate750(.a(gate43inter0), .b(s_78), .O(gate43inter1));
  and2  gate751(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate752(.a(s_78), .O(gate43inter3));
  inv1  gate753(.a(s_79), .O(gate43inter4));
  nand2 gate754(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate755(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate756(.a(N254), .O(gate43inter7));
  inv1  gate757(.a(N255), .O(gate43inter8));
  nand2 gate758(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate759(.a(s_79), .b(gate43inter3), .O(gate43inter10));
  nor2  gate760(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate761(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate762(.a(gate43inter12), .b(gate43inter1), .O(N296));

  xor2  gate1407(.a(N257), .b(N256), .O(gate44inter0));
  nand2 gate1408(.a(gate44inter0), .b(s_172), .O(gate44inter1));
  and2  gate1409(.a(N257), .b(N256), .O(gate44inter2));
  inv1  gate1410(.a(s_172), .O(gate44inter3));
  inv1  gate1411(.a(s_173), .O(gate44inter4));
  nand2 gate1412(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1413(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1414(.a(N256), .O(gate44inter7));
  inv1  gate1415(.a(N257), .O(gate44inter8));
  nand2 gate1416(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1417(.a(s_173), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1418(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1419(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1420(.a(gate44inter12), .b(gate44inter1), .O(N299));

  xor2  gate567(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate568(.a(gate45inter0), .b(s_52), .O(gate45inter1));
  and2  gate569(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate570(.a(s_52), .O(gate45inter3));
  inv1  gate571(.a(s_53), .O(gate45inter4));
  nand2 gate572(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate573(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate574(.a(N258), .O(gate45inter7));
  inv1  gate575(.a(N259), .O(gate45inter8));
  nand2 gate576(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate577(.a(s_53), .b(gate45inter3), .O(gate45inter10));
  nor2  gate578(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate579(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate580(.a(gate45inter12), .b(gate45inter1), .O(N302));

  xor2  gate1295(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate1296(.a(gate46inter0), .b(s_156), .O(gate46inter1));
  and2  gate1297(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate1298(.a(s_156), .O(gate46inter3));
  inv1  gate1299(.a(s_157), .O(gate46inter4));
  nand2 gate1300(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1301(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1302(.a(N260), .O(gate46inter7));
  inv1  gate1303(.a(N261), .O(gate46inter8));
  nand2 gate1304(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1305(.a(s_157), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1306(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1307(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1308(.a(gate46inter12), .b(gate46inter1), .O(N305));

  xor2  gate623(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate624(.a(gate47inter0), .b(s_60), .O(gate47inter1));
  and2  gate625(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate626(.a(s_60), .O(gate47inter3));
  inv1  gate627(.a(s_61), .O(gate47inter4));
  nand2 gate628(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate629(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate630(.a(N262), .O(gate47inter7));
  inv1  gate631(.a(N263), .O(gate47inter8));
  nand2 gate632(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate633(.a(s_61), .b(gate47inter3), .O(gate47inter10));
  nor2  gate634(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate635(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate636(.a(gate47inter12), .b(gate47inter1), .O(N308));

  xor2  gate1127(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate1128(.a(gate48inter0), .b(s_132), .O(gate48inter1));
  and2  gate1129(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate1130(.a(s_132), .O(gate48inter3));
  inv1  gate1131(.a(s_133), .O(gate48inter4));
  nand2 gate1132(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1133(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1134(.a(N264), .O(gate48inter7));
  inv1  gate1135(.a(N265), .O(gate48inter8));
  nand2 gate1136(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1137(.a(s_133), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1138(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1139(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1140(.a(gate48inter12), .b(gate48inter1), .O(N311));

  xor2  gate1183(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate1184(.a(gate49inter0), .b(s_140), .O(gate49inter1));
  and2  gate1185(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate1186(.a(s_140), .O(gate49inter3));
  inv1  gate1187(.a(s_141), .O(gate49inter4));
  nand2 gate1188(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1189(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1190(.a(N274), .O(gate49inter7));
  inv1  gate1191(.a(N275), .O(gate49inter8));
  nand2 gate1192(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1193(.a(s_141), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1194(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1195(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1196(.a(gate49inter12), .b(gate49inter1), .O(N314));

  xor2  gate595(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate596(.a(gate50inter0), .b(s_56), .O(gate50inter1));
  and2  gate597(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate598(.a(s_56), .O(gate50inter3));
  inv1  gate599(.a(s_57), .O(gate50inter4));
  nand2 gate600(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate601(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate602(.a(N276), .O(gate50inter7));
  inv1  gate603(.a(N277), .O(gate50inter8));
  nand2 gate604(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate605(.a(s_57), .b(gate50inter3), .O(gate50inter10));
  nor2  gate606(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate607(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate608(.a(gate50inter12), .b(gate50inter1), .O(N315));

  xor2  gate903(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate904(.a(gate51inter0), .b(s_100), .O(gate51inter1));
  and2  gate905(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate906(.a(s_100), .O(gate51inter3));
  inv1  gate907(.a(s_101), .O(gate51inter4));
  nand2 gate908(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate909(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate910(.a(N278), .O(gate51inter7));
  inv1  gate911(.a(N279), .O(gate51inter8));
  nand2 gate912(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate913(.a(s_101), .b(gate51inter3), .O(gate51inter10));
  nor2  gate914(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate915(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate916(.a(gate51inter12), .b(gate51inter1), .O(N316));

  xor2  gate581(.a(N281), .b(N280), .O(gate52inter0));
  nand2 gate582(.a(gate52inter0), .b(s_54), .O(gate52inter1));
  and2  gate583(.a(N281), .b(N280), .O(gate52inter2));
  inv1  gate584(.a(s_54), .O(gate52inter3));
  inv1  gate585(.a(s_55), .O(gate52inter4));
  nand2 gate586(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate587(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate588(.a(N280), .O(gate52inter7));
  inv1  gate589(.a(N281), .O(gate52inter8));
  nand2 gate590(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate591(.a(s_55), .b(gate52inter3), .O(gate52inter10));
  nor2  gate592(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate593(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate594(.a(gate52inter12), .b(gate52inter1), .O(N317));

  xor2  gate1449(.a(N283), .b(N282), .O(gate53inter0));
  nand2 gate1450(.a(gate53inter0), .b(s_178), .O(gate53inter1));
  and2  gate1451(.a(N283), .b(N282), .O(gate53inter2));
  inv1  gate1452(.a(s_178), .O(gate53inter3));
  inv1  gate1453(.a(s_179), .O(gate53inter4));
  nand2 gate1454(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1455(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1456(.a(N282), .O(gate53inter7));
  inv1  gate1457(.a(N283), .O(gate53inter8));
  nand2 gate1458(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1459(.a(s_179), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1460(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1461(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1462(.a(gate53inter12), .b(gate53inter1), .O(N318));

  xor2  gate329(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate330(.a(gate54inter0), .b(s_18), .O(gate54inter1));
  and2  gate331(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate332(.a(s_18), .O(gate54inter3));
  inv1  gate333(.a(s_19), .O(gate54inter4));
  nand2 gate334(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate335(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate336(.a(N284), .O(gate54inter7));
  inv1  gate337(.a(N285), .O(gate54inter8));
  nand2 gate338(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate339(.a(s_19), .b(gate54inter3), .O(gate54inter10));
  nor2  gate340(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate341(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate342(.a(gate54inter12), .b(gate54inter1), .O(N319));

  xor2  gate1239(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate1240(.a(gate55inter0), .b(s_148), .O(gate55inter1));
  and2  gate1241(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate1242(.a(s_148), .O(gate55inter3));
  inv1  gate1243(.a(s_149), .O(gate55inter4));
  nand2 gate1244(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1245(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1246(.a(N286), .O(gate55inter7));
  inv1  gate1247(.a(N287), .O(gate55inter8));
  nand2 gate1248(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1249(.a(s_149), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1250(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1251(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1252(.a(gate55inter12), .b(gate55inter1), .O(N320));

  xor2  gate1281(.a(N289), .b(N288), .O(gate56inter0));
  nand2 gate1282(.a(gate56inter0), .b(s_154), .O(gate56inter1));
  and2  gate1283(.a(N289), .b(N288), .O(gate56inter2));
  inv1  gate1284(.a(s_154), .O(gate56inter3));
  inv1  gate1285(.a(s_155), .O(gate56inter4));
  nand2 gate1286(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1287(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1288(.a(N288), .O(gate56inter7));
  inv1  gate1289(.a(N289), .O(gate56inter8));
  nand2 gate1290(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1291(.a(s_155), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1292(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1293(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1294(.a(gate56inter12), .b(gate56inter1), .O(N321));

  xor2  gate553(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate554(.a(gate57inter0), .b(s_50), .O(gate57inter1));
  and2  gate555(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate556(.a(s_50), .O(gate57inter3));
  inv1  gate557(.a(s_51), .O(gate57inter4));
  nand2 gate558(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate559(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate560(.a(N290), .O(gate57inter7));
  inv1  gate561(.a(N293), .O(gate57inter8));
  nand2 gate562(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate563(.a(s_51), .b(gate57inter3), .O(gate57inter10));
  nor2  gate564(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate565(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate566(.a(gate57inter12), .b(gate57inter1), .O(N338));

  xor2  gate1351(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate1352(.a(gate58inter0), .b(s_164), .O(gate58inter1));
  and2  gate1353(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate1354(.a(s_164), .O(gate58inter3));
  inv1  gate1355(.a(s_165), .O(gate58inter4));
  nand2 gate1356(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1357(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1358(.a(N296), .O(gate58inter7));
  inv1  gate1359(.a(N299), .O(gate58inter8));
  nand2 gate1360(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1361(.a(s_165), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1362(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1363(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1364(.a(gate58inter12), .b(gate58inter1), .O(N339));

  xor2  gate217(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate218(.a(gate59inter0), .b(s_2), .O(gate59inter1));
  and2  gate219(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate220(.a(s_2), .O(gate59inter3));
  inv1  gate221(.a(s_3), .O(gate59inter4));
  nand2 gate222(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate223(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate224(.a(N290), .O(gate59inter7));
  inv1  gate225(.a(N296), .O(gate59inter8));
  nand2 gate226(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate227(.a(s_3), .b(gate59inter3), .O(gate59inter10));
  nor2  gate228(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate229(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate230(.a(gate59inter12), .b(gate59inter1), .O(N340));
xor2 gate60( .a(N293), .b(N299), .O(N341) );

  xor2  gate833(.a(N305), .b(N302), .O(gate61inter0));
  nand2 gate834(.a(gate61inter0), .b(s_90), .O(gate61inter1));
  and2  gate835(.a(N305), .b(N302), .O(gate61inter2));
  inv1  gate836(.a(s_90), .O(gate61inter3));
  inv1  gate837(.a(s_91), .O(gate61inter4));
  nand2 gate838(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate839(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate840(.a(N302), .O(gate61inter7));
  inv1  gate841(.a(N305), .O(gate61inter8));
  nand2 gate842(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate843(.a(s_91), .b(gate61inter3), .O(gate61inter10));
  nor2  gate844(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate845(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate846(.a(gate61inter12), .b(gate61inter1), .O(N342));

  xor2  gate203(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate204(.a(gate62inter0), .b(s_0), .O(gate62inter1));
  and2  gate205(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate206(.a(s_0), .O(gate62inter3));
  inv1  gate207(.a(s_1), .O(gate62inter4));
  nand2 gate208(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate209(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate210(.a(N308), .O(gate62inter7));
  inv1  gate211(.a(N311), .O(gate62inter8));
  nand2 gate212(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate213(.a(s_1), .b(gate62inter3), .O(gate62inter10));
  nor2  gate214(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate215(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate216(.a(gate62inter12), .b(gate62inter1), .O(N343));

  xor2  gate1463(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate1464(.a(gate63inter0), .b(s_180), .O(gate63inter1));
  and2  gate1465(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate1466(.a(s_180), .O(gate63inter3));
  inv1  gate1467(.a(s_181), .O(gate63inter4));
  nand2 gate1468(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1469(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1470(.a(N302), .O(gate63inter7));
  inv1  gate1471(.a(N308), .O(gate63inter8));
  nand2 gate1472(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1473(.a(s_181), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1474(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1475(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1476(.a(gate63inter12), .b(gate63inter1), .O(N344));

  xor2  gate455(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate456(.a(gate64inter0), .b(s_36), .O(gate64inter1));
  and2  gate457(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate458(.a(s_36), .O(gate64inter3));
  inv1  gate459(.a(s_37), .O(gate64inter4));
  nand2 gate460(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate461(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate462(.a(N305), .O(gate64inter7));
  inv1  gate463(.a(N311), .O(gate64inter8));
  nand2 gate464(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate465(.a(s_37), .b(gate64inter3), .O(gate64inter10));
  nor2  gate466(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate467(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate468(.a(gate64inter12), .b(gate64inter1), .O(N345));

  xor2  gate1211(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate1212(.a(gate65inter0), .b(s_144), .O(gate65inter1));
  and2  gate1213(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate1214(.a(s_144), .O(gate65inter3));
  inv1  gate1215(.a(s_145), .O(gate65inter4));
  nand2 gate1216(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1217(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1218(.a(N266), .O(gate65inter7));
  inv1  gate1219(.a(N342), .O(gate65inter8));
  nand2 gate1220(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1221(.a(s_145), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1222(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1223(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1224(.a(gate65inter12), .b(gate65inter1), .O(N346));

  xor2  gate231(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate232(.a(gate66inter0), .b(s_4), .O(gate66inter1));
  and2  gate233(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate234(.a(s_4), .O(gate66inter3));
  inv1  gate235(.a(s_5), .O(gate66inter4));
  nand2 gate236(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate237(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate238(.a(N267), .O(gate66inter7));
  inv1  gate239(.a(N343), .O(gate66inter8));
  nand2 gate240(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate241(.a(s_5), .b(gate66inter3), .O(gate66inter10));
  nor2  gate242(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate243(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate244(.a(gate66inter12), .b(gate66inter1), .O(N347));

  xor2  gate287(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate288(.a(gate67inter0), .b(s_12), .O(gate67inter1));
  and2  gate289(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate290(.a(s_12), .O(gate67inter3));
  inv1  gate291(.a(s_13), .O(gate67inter4));
  nand2 gate292(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate293(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate294(.a(N268), .O(gate67inter7));
  inv1  gate295(.a(N344), .O(gate67inter8));
  nand2 gate296(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate297(.a(s_13), .b(gate67inter3), .O(gate67inter10));
  nor2  gate298(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate299(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate300(.a(gate67inter12), .b(gate67inter1), .O(N348));
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate861(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate862(.a(gate70inter0), .b(s_94), .O(gate70inter1));
  and2  gate863(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate864(.a(s_94), .O(gate70inter3));
  inv1  gate865(.a(s_95), .O(gate70inter4));
  nand2 gate866(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate867(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate868(.a(N271), .O(gate70inter7));
  inv1  gate869(.a(N339), .O(gate70inter8));
  nand2 gate870(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate871(.a(s_95), .b(gate70inter3), .O(gate70inter10));
  nor2  gate872(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate873(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate874(.a(gate70inter12), .b(gate70inter1), .O(N351));

  xor2  gate413(.a(N340), .b(N272), .O(gate71inter0));
  nand2 gate414(.a(gate71inter0), .b(s_30), .O(gate71inter1));
  and2  gate415(.a(N340), .b(N272), .O(gate71inter2));
  inv1  gate416(.a(s_30), .O(gate71inter3));
  inv1  gate417(.a(s_31), .O(gate71inter4));
  nand2 gate418(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate419(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate420(.a(N272), .O(gate71inter7));
  inv1  gate421(.a(N340), .O(gate71inter8));
  nand2 gate422(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate423(.a(s_31), .b(gate71inter3), .O(gate71inter10));
  nor2  gate424(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate425(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate426(.a(gate71inter12), .b(gate71inter1), .O(N352));
xor2 gate72( .a(N273), .b(N341), .O(N353) );

  xor2  gate1113(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate1114(.a(gate73inter0), .b(s_130), .O(gate73inter1));
  and2  gate1115(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate1116(.a(s_130), .O(gate73inter3));
  inv1  gate1117(.a(s_131), .O(gate73inter4));
  nand2 gate1118(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1119(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1120(.a(N314), .O(gate73inter7));
  inv1  gate1121(.a(N346), .O(gate73inter8));
  nand2 gate1122(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1123(.a(s_131), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1124(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1125(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1126(.a(gate73inter12), .b(gate73inter1), .O(N354));

  xor2  gate1085(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate1086(.a(gate74inter0), .b(s_126), .O(gate74inter1));
  and2  gate1087(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate1088(.a(s_126), .O(gate74inter3));
  inv1  gate1089(.a(s_127), .O(gate74inter4));
  nand2 gate1090(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1091(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1092(.a(N315), .O(gate74inter7));
  inv1  gate1093(.a(N347), .O(gate74inter8));
  nand2 gate1094(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1095(.a(s_127), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1096(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1097(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1098(.a(gate74inter12), .b(gate74inter1), .O(N367));

  xor2  gate875(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate876(.a(gate75inter0), .b(s_96), .O(gate75inter1));
  and2  gate877(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate878(.a(s_96), .O(gate75inter3));
  inv1  gate879(.a(s_97), .O(gate75inter4));
  nand2 gate880(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate881(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate882(.a(N316), .O(gate75inter7));
  inv1  gate883(.a(N348), .O(gate75inter8));
  nand2 gate884(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate885(.a(s_97), .b(gate75inter3), .O(gate75inter10));
  nor2  gate886(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate887(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate888(.a(gate75inter12), .b(gate75inter1), .O(N380));

  xor2  gate273(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate274(.a(gate76inter0), .b(s_10), .O(gate76inter1));
  and2  gate275(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate276(.a(s_10), .O(gate76inter3));
  inv1  gate277(.a(s_11), .O(gate76inter4));
  nand2 gate278(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate279(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate280(.a(N317), .O(gate76inter7));
  inv1  gate281(.a(N349), .O(gate76inter8));
  nand2 gate282(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate283(.a(s_11), .b(gate76inter3), .O(gate76inter10));
  nor2  gate284(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate285(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate286(.a(gate76inter12), .b(gate76inter1), .O(N393));

  xor2  gate1365(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate1366(.a(gate77inter0), .b(s_166), .O(gate77inter1));
  and2  gate1367(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate1368(.a(s_166), .O(gate77inter3));
  inv1  gate1369(.a(s_167), .O(gate77inter4));
  nand2 gate1370(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1371(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1372(.a(N318), .O(gate77inter7));
  inv1  gate1373(.a(N350), .O(gate77inter8));
  nand2 gate1374(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1375(.a(s_167), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1376(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1377(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1378(.a(gate77inter12), .b(gate77inter1), .O(N406));

  xor2  gate525(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate526(.a(gate78inter0), .b(s_46), .O(gate78inter1));
  and2  gate527(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate528(.a(s_46), .O(gate78inter3));
  inv1  gate529(.a(s_47), .O(gate78inter4));
  nand2 gate530(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate531(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate532(.a(N319), .O(gate78inter7));
  inv1  gate533(.a(N351), .O(gate78inter8));
  nand2 gate534(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate535(.a(s_47), .b(gate78inter3), .O(gate78inter10));
  nor2  gate536(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate537(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate538(.a(gate78inter12), .b(gate78inter1), .O(N419));

  xor2  gate497(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate498(.a(gate79inter0), .b(s_42), .O(gate79inter1));
  and2  gate499(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate500(.a(s_42), .O(gate79inter3));
  inv1  gate501(.a(s_43), .O(gate79inter4));
  nand2 gate502(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate503(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate504(.a(N320), .O(gate79inter7));
  inv1  gate505(.a(N352), .O(gate79inter8));
  nand2 gate506(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate507(.a(s_43), .b(gate79inter3), .O(gate79inter10));
  nor2  gate508(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate509(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate510(.a(gate79inter12), .b(gate79inter1), .O(N432));

  xor2  gate1043(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate1044(.a(gate80inter0), .b(s_120), .O(gate80inter1));
  and2  gate1045(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate1046(.a(s_120), .O(gate80inter3));
  inv1  gate1047(.a(s_121), .O(gate80inter4));
  nand2 gate1048(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1049(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1050(.a(N321), .O(gate80inter7));
  inv1  gate1051(.a(N353), .O(gate80inter8));
  nand2 gate1052(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1053(.a(s_121), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1054(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1055(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1056(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );

  xor2  gate1323(.a(N692), .b(N1), .O(gate171inter0));
  nand2 gate1324(.a(gate171inter0), .b(s_160), .O(gate171inter1));
  and2  gate1325(.a(N692), .b(N1), .O(gate171inter2));
  inv1  gate1326(.a(s_160), .O(gate171inter3));
  inv1  gate1327(.a(s_161), .O(gate171inter4));
  nand2 gate1328(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1329(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1330(.a(N1), .O(gate171inter7));
  inv1  gate1331(.a(N692), .O(gate171inter8));
  nand2 gate1332(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1333(.a(s_161), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1334(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1335(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1336(.a(gate171inter12), .b(gate171inter1), .O(N724));
xor2 gate172( .a(N5), .b(N693), .O(N725) );

  xor2  gate847(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate848(.a(gate173inter0), .b(s_92), .O(gate173inter1));
  and2  gate849(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate850(.a(s_92), .O(gate173inter3));
  inv1  gate851(.a(s_93), .O(gate173inter4));
  nand2 gate852(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate853(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate854(.a(N9), .O(gate173inter7));
  inv1  gate855(.a(N694), .O(gate173inter8));
  nand2 gate856(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate857(.a(s_93), .b(gate173inter3), .O(gate173inter10));
  nor2  gate858(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate859(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate860(.a(gate173inter12), .b(gate173inter1), .O(N726));

  xor2  gate357(.a(N695), .b(N13), .O(gate174inter0));
  nand2 gate358(.a(gate174inter0), .b(s_22), .O(gate174inter1));
  and2  gate359(.a(N695), .b(N13), .O(gate174inter2));
  inv1  gate360(.a(s_22), .O(gate174inter3));
  inv1  gate361(.a(s_23), .O(gate174inter4));
  nand2 gate362(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate363(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate364(.a(N13), .O(gate174inter7));
  inv1  gate365(.a(N695), .O(gate174inter8));
  nand2 gate366(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate367(.a(s_23), .b(gate174inter3), .O(gate174inter10));
  nor2  gate368(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate369(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate370(.a(gate174inter12), .b(gate174inter1), .O(N727));

  xor2  gate1309(.a(N696), .b(N17), .O(gate175inter0));
  nand2 gate1310(.a(gate175inter0), .b(s_158), .O(gate175inter1));
  and2  gate1311(.a(N696), .b(N17), .O(gate175inter2));
  inv1  gate1312(.a(s_158), .O(gate175inter3));
  inv1  gate1313(.a(s_159), .O(gate175inter4));
  nand2 gate1314(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1315(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1316(.a(N17), .O(gate175inter7));
  inv1  gate1317(.a(N696), .O(gate175inter8));
  nand2 gate1318(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1319(.a(s_159), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1320(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1321(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1322(.a(gate175inter12), .b(gate175inter1), .O(N728));

  xor2  gate889(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate890(.a(gate176inter0), .b(s_98), .O(gate176inter1));
  and2  gate891(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate892(.a(s_98), .O(gate176inter3));
  inv1  gate893(.a(s_99), .O(gate176inter4));
  nand2 gate894(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate895(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate896(.a(N21), .O(gate176inter7));
  inv1  gate897(.a(N697), .O(gate176inter8));
  nand2 gate898(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate899(.a(s_99), .b(gate176inter3), .O(gate176inter10));
  nor2  gate900(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate901(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate902(.a(gate176inter12), .b(gate176inter1), .O(N729));

  xor2  gate959(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate960(.a(gate177inter0), .b(s_108), .O(gate177inter1));
  and2  gate961(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate962(.a(s_108), .O(gate177inter3));
  inv1  gate963(.a(s_109), .O(gate177inter4));
  nand2 gate964(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate965(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate966(.a(N25), .O(gate177inter7));
  inv1  gate967(.a(N698), .O(gate177inter8));
  nand2 gate968(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate969(.a(s_109), .b(gate177inter3), .O(gate177inter10));
  nor2  gate970(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate971(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate972(.a(gate177inter12), .b(gate177inter1), .O(N730));

  xor2  gate651(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate652(.a(gate178inter0), .b(s_64), .O(gate178inter1));
  and2  gate653(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate654(.a(s_64), .O(gate178inter3));
  inv1  gate655(.a(s_65), .O(gate178inter4));
  nand2 gate656(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate657(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate658(.a(N29), .O(gate178inter7));
  inv1  gate659(.a(N699), .O(gate178inter8));
  nand2 gate660(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate661(.a(s_65), .b(gate178inter3), .O(gate178inter10));
  nor2  gate662(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate663(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate664(.a(gate178inter12), .b(gate178inter1), .O(N731));

  xor2  gate427(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate428(.a(gate179inter0), .b(s_32), .O(gate179inter1));
  and2  gate429(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate430(.a(s_32), .O(gate179inter3));
  inv1  gate431(.a(s_33), .O(gate179inter4));
  nand2 gate432(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate433(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate434(.a(N33), .O(gate179inter7));
  inv1  gate435(.a(N700), .O(gate179inter8));
  nand2 gate436(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate437(.a(s_33), .b(gate179inter3), .O(gate179inter10));
  nor2  gate438(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate439(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate440(.a(gate179inter12), .b(gate179inter1), .O(N732));

  xor2  gate315(.a(N701), .b(N37), .O(gate180inter0));
  nand2 gate316(.a(gate180inter0), .b(s_16), .O(gate180inter1));
  and2  gate317(.a(N701), .b(N37), .O(gate180inter2));
  inv1  gate318(.a(s_16), .O(gate180inter3));
  inv1  gate319(.a(s_17), .O(gate180inter4));
  nand2 gate320(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate321(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate322(.a(N37), .O(gate180inter7));
  inv1  gate323(.a(N701), .O(gate180inter8));
  nand2 gate324(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate325(.a(s_17), .b(gate180inter3), .O(gate180inter10));
  nor2  gate326(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate327(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate328(.a(gate180inter12), .b(gate180inter1), .O(N733));

  xor2  gate777(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate778(.a(gate181inter0), .b(s_82), .O(gate181inter1));
  and2  gate779(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate780(.a(s_82), .O(gate181inter3));
  inv1  gate781(.a(s_83), .O(gate181inter4));
  nand2 gate782(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate783(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate784(.a(N41), .O(gate181inter7));
  inv1  gate785(.a(N702), .O(gate181inter8));
  nand2 gate786(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate787(.a(s_83), .b(gate181inter3), .O(gate181inter10));
  nor2  gate788(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate789(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate790(.a(gate181inter12), .b(gate181inter1), .O(N734));

  xor2  gate1267(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate1268(.a(gate182inter0), .b(s_152), .O(gate182inter1));
  and2  gate1269(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate1270(.a(s_152), .O(gate182inter3));
  inv1  gate1271(.a(s_153), .O(gate182inter4));
  nand2 gate1272(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1273(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1274(.a(N45), .O(gate182inter7));
  inv1  gate1275(.a(N703), .O(gate182inter8));
  nand2 gate1276(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1277(.a(s_153), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1278(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1279(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1280(.a(gate182inter12), .b(gate182inter1), .O(N735));

  xor2  gate609(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate610(.a(gate183inter0), .b(s_58), .O(gate183inter1));
  and2  gate611(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate612(.a(s_58), .O(gate183inter3));
  inv1  gate613(.a(s_59), .O(gate183inter4));
  nand2 gate614(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate615(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate616(.a(N49), .O(gate183inter7));
  inv1  gate617(.a(N704), .O(gate183inter8));
  nand2 gate618(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate619(.a(s_59), .b(gate183inter3), .O(gate183inter10));
  nor2  gate620(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate621(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate622(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );

  xor2  gate469(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate470(.a(gate185inter0), .b(s_38), .O(gate185inter1));
  and2  gate471(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate472(.a(s_38), .O(gate185inter3));
  inv1  gate473(.a(s_39), .O(gate185inter4));
  nand2 gate474(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate475(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate476(.a(N57), .O(gate185inter7));
  inv1  gate477(.a(N706), .O(gate185inter8));
  nand2 gate478(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate479(.a(s_39), .b(gate185inter3), .O(gate185inter10));
  nor2  gate480(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate481(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate482(.a(gate185inter12), .b(gate185inter1), .O(N738));

  xor2  gate707(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate708(.a(gate186inter0), .b(s_72), .O(gate186inter1));
  and2  gate709(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate710(.a(s_72), .O(gate186inter3));
  inv1  gate711(.a(s_73), .O(gate186inter4));
  nand2 gate712(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate713(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate714(.a(N61), .O(gate186inter7));
  inv1  gate715(.a(N707), .O(gate186inter8));
  nand2 gate716(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate717(.a(s_73), .b(gate186inter3), .O(gate186inter10));
  nor2  gate718(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate719(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate720(.a(gate186inter12), .b(gate186inter1), .O(N739));

  xor2  gate637(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate638(.a(gate187inter0), .b(s_62), .O(gate187inter1));
  and2  gate639(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate640(.a(s_62), .O(gate187inter3));
  inv1  gate641(.a(s_63), .O(gate187inter4));
  nand2 gate642(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate643(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate644(.a(N65), .O(gate187inter7));
  inv1  gate645(.a(N708), .O(gate187inter8));
  nand2 gate646(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate647(.a(s_63), .b(gate187inter3), .O(gate187inter10));
  nor2  gate648(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate649(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate650(.a(gate187inter12), .b(gate187inter1), .O(N740));

  xor2  gate385(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate386(.a(gate188inter0), .b(s_26), .O(gate188inter1));
  and2  gate387(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate388(.a(s_26), .O(gate188inter3));
  inv1  gate389(.a(s_27), .O(gate188inter4));
  nand2 gate390(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate391(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate392(.a(N69), .O(gate188inter7));
  inv1  gate393(.a(N709), .O(gate188inter8));
  nand2 gate394(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate395(.a(s_27), .b(gate188inter3), .O(gate188inter10));
  nor2  gate396(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate397(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate398(.a(gate188inter12), .b(gate188inter1), .O(N741));

  xor2  gate1337(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate1338(.a(gate189inter0), .b(s_162), .O(gate189inter1));
  and2  gate1339(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate1340(.a(s_162), .O(gate189inter3));
  inv1  gate1341(.a(s_163), .O(gate189inter4));
  nand2 gate1342(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1343(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1344(.a(N73), .O(gate189inter7));
  inv1  gate1345(.a(N710), .O(gate189inter8));
  nand2 gate1346(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1347(.a(s_163), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1348(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1349(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1350(.a(gate189inter12), .b(gate189inter1), .O(N742));

  xor2  gate693(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate694(.a(gate190inter0), .b(s_70), .O(gate190inter1));
  and2  gate695(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate696(.a(s_70), .O(gate190inter3));
  inv1  gate697(.a(s_71), .O(gate190inter4));
  nand2 gate698(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate699(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate700(.a(N77), .O(gate190inter7));
  inv1  gate701(.a(N711), .O(gate190inter8));
  nand2 gate702(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate703(.a(s_71), .b(gate190inter3), .O(gate190inter10));
  nor2  gate704(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate705(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate706(.a(gate190inter12), .b(gate190inter1), .O(N743));

  xor2  gate1099(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate1100(.a(gate191inter0), .b(s_128), .O(gate191inter1));
  and2  gate1101(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate1102(.a(s_128), .O(gate191inter3));
  inv1  gate1103(.a(s_129), .O(gate191inter4));
  nand2 gate1104(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1105(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1106(.a(N81), .O(gate191inter7));
  inv1  gate1107(.a(N712), .O(gate191inter8));
  nand2 gate1108(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1109(.a(s_129), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1110(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1111(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1112(.a(gate191inter12), .b(gate191inter1), .O(N744));

  xor2  gate1015(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate1016(.a(gate192inter0), .b(s_116), .O(gate192inter1));
  and2  gate1017(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate1018(.a(s_116), .O(gate192inter3));
  inv1  gate1019(.a(s_117), .O(gate192inter4));
  nand2 gate1020(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1021(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1022(.a(N85), .O(gate192inter7));
  inv1  gate1023(.a(N713), .O(gate192inter8));
  nand2 gate1024(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1025(.a(s_117), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1026(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1027(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1028(.a(gate192inter12), .b(gate192inter1), .O(N745));
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );

  xor2  gate301(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate302(.a(gate196inter0), .b(s_14), .O(gate196inter1));
  and2  gate303(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate304(.a(s_14), .O(gate196inter3));
  inv1  gate305(.a(s_15), .O(gate196inter4));
  nand2 gate306(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate307(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate308(.a(N101), .O(gate196inter7));
  inv1  gate309(.a(N717), .O(gate196inter8));
  nand2 gate310(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate311(.a(s_15), .b(gate196inter3), .O(gate196inter10));
  nor2  gate312(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate313(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate314(.a(gate196inter12), .b(gate196inter1), .O(N749));

  xor2  gate1057(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate1058(.a(gate197inter0), .b(s_122), .O(gate197inter1));
  and2  gate1059(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate1060(.a(s_122), .O(gate197inter3));
  inv1  gate1061(.a(s_123), .O(gate197inter4));
  nand2 gate1062(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1063(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1064(.a(N105), .O(gate197inter7));
  inv1  gate1065(.a(N718), .O(gate197inter8));
  nand2 gate1066(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1067(.a(s_123), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1068(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1069(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1070(.a(gate197inter12), .b(gate197inter1), .O(N750));
xor2 gate198( .a(N109), .b(N719), .O(N751) );

  xor2  gate917(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate918(.a(gate199inter0), .b(s_102), .O(gate199inter1));
  and2  gate919(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate920(.a(s_102), .O(gate199inter3));
  inv1  gate921(.a(s_103), .O(gate199inter4));
  nand2 gate922(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate923(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate924(.a(N113), .O(gate199inter7));
  inv1  gate925(.a(N720), .O(gate199inter8));
  nand2 gate926(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate927(.a(s_103), .b(gate199inter3), .O(gate199inter10));
  nor2  gate928(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate929(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate930(.a(gate199inter12), .b(gate199inter1), .O(N752));

  xor2  gate679(.a(N721), .b(N117), .O(gate200inter0));
  nand2 gate680(.a(gate200inter0), .b(s_68), .O(gate200inter1));
  and2  gate681(.a(N721), .b(N117), .O(gate200inter2));
  inv1  gate682(.a(s_68), .O(gate200inter3));
  inv1  gate683(.a(s_69), .O(gate200inter4));
  nand2 gate684(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate685(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate686(.a(N117), .O(gate200inter7));
  inv1  gate687(.a(N721), .O(gate200inter8));
  nand2 gate688(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate689(.a(s_69), .b(gate200inter3), .O(gate200inter10));
  nor2  gate690(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate691(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate692(.a(gate200inter12), .b(gate200inter1), .O(N753));

  xor2  gate973(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate974(.a(gate201inter0), .b(s_110), .O(gate201inter1));
  and2  gate975(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate976(.a(s_110), .O(gate201inter3));
  inv1  gate977(.a(s_111), .O(gate201inter4));
  nand2 gate978(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate979(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate980(.a(N121), .O(gate201inter7));
  inv1  gate981(.a(N722), .O(gate201inter8));
  nand2 gate982(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate983(.a(s_111), .b(gate201inter3), .O(gate201inter10));
  nor2  gate984(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate985(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate986(.a(gate201inter12), .b(gate201inter1), .O(N754));

  xor2  gate1155(.a(N723), .b(N125), .O(gate202inter0));
  nand2 gate1156(.a(gate202inter0), .b(s_136), .O(gate202inter1));
  and2  gate1157(.a(N723), .b(N125), .O(gate202inter2));
  inv1  gate1158(.a(s_136), .O(gate202inter3));
  inv1  gate1159(.a(s_137), .O(gate202inter4));
  nand2 gate1160(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1161(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1162(.a(N125), .O(gate202inter7));
  inv1  gate1163(.a(N723), .O(gate202inter8));
  nand2 gate1164(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1165(.a(s_137), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1166(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1167(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1168(.a(gate202inter12), .b(gate202inter1), .O(N755));

endmodule