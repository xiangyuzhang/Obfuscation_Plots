module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate385(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate386(.a(gate19inter0), .b(s_32), .O(gate19inter1));
  and2  gate387(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate388(.a(s_32), .O(gate19inter3));
  inv1  gate389(.a(s_33), .O(gate19inter4));
  nand2 gate390(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate391(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate392(.a(N118), .O(gate19inter7));
  inv1  gate393(.a(N4), .O(gate19inter8));
  nand2 gate394(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate395(.a(s_33), .b(gate19inter3), .O(gate19inter10));
  nor2  gate396(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate397(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate398(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate511(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate512(.a(gate20inter0), .b(s_50), .O(gate20inter1));
  and2  gate513(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate514(.a(s_50), .O(gate20inter3));
  inv1  gate515(.a(s_51), .O(gate20inter4));
  nand2 gate516(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate517(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate518(.a(N8), .O(gate20inter7));
  inv1  gate519(.a(N119), .O(gate20inter8));
  nand2 gate520(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate521(.a(s_51), .b(gate20inter3), .O(gate20inter10));
  nor2  gate522(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate523(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate524(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate469(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate470(.a(gate24inter0), .b(s_44), .O(gate24inter1));
  and2  gate471(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate472(.a(s_44), .O(gate24inter3));
  inv1  gate473(.a(s_45), .O(gate24inter4));
  nand2 gate474(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate475(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate476(.a(N130), .O(gate24inter7));
  inv1  gate477(.a(N43), .O(gate24inter8));
  nand2 gate478(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate479(.a(s_45), .b(gate24inter3), .O(gate24inter10));
  nor2  gate480(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate481(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate482(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );

  xor2  gate343(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate344(.a(gate26inter0), .b(s_26), .O(gate26inter1));
  and2  gate345(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate346(.a(s_26), .O(gate26inter3));
  inv1  gate347(.a(s_27), .O(gate26inter4));
  nand2 gate348(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate349(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate350(.a(N138), .O(gate26inter7));
  inv1  gate351(.a(N69), .O(gate26inter8));
  nand2 gate352(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate353(.a(s_27), .b(gate26inter3), .O(gate26inter10));
  nor2  gate354(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate355(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate356(.a(gate26inter12), .b(gate26inter1), .O(N171));
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate609(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate610(.a(gate28inter0), .b(s_64), .O(gate28inter1));
  and2  gate611(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate612(.a(s_64), .O(gate28inter3));
  inv1  gate613(.a(s_65), .O(gate28inter4));
  nand2 gate614(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate615(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate616(.a(N146), .O(gate28inter7));
  inv1  gate617(.a(N95), .O(gate28inter8));
  nand2 gate618(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate619(.a(s_65), .b(gate28inter3), .O(gate28inter10));
  nor2  gate620(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate621(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate622(.a(gate28inter12), .b(gate28inter1), .O(N177));

  xor2  gate413(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate414(.a(gate29inter0), .b(s_36), .O(gate29inter1));
  and2  gate415(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate416(.a(s_36), .O(gate29inter3));
  inv1  gate417(.a(s_37), .O(gate29inter4));
  nand2 gate418(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate419(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate420(.a(N150), .O(gate29inter7));
  inv1  gate421(.a(N108), .O(gate29inter8));
  nand2 gate422(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate423(.a(s_37), .b(gate29inter3), .O(gate29inter10));
  nor2  gate424(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate425(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate426(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );

  xor2  gate567(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate568(.a(gate31inter0), .b(s_58), .O(gate31inter1));
  and2  gate569(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate570(.a(s_58), .O(gate31inter3));
  inv1  gate571(.a(s_59), .O(gate31inter4));
  nand2 gate572(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate573(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate574(.a(N27), .O(gate31inter7));
  inv1  gate575(.a(N123), .O(gate31inter8));
  nand2 gate576(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate577(.a(s_59), .b(gate31inter3), .O(gate31inter10));
  nor2  gate578(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate579(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate580(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );

  xor2  gate231(.a(N127), .b(N40), .O(gate33inter0));
  nand2 gate232(.a(gate33inter0), .b(s_10), .O(gate33inter1));
  and2  gate233(.a(N127), .b(N40), .O(gate33inter2));
  inv1  gate234(.a(s_10), .O(gate33inter3));
  inv1  gate235(.a(s_11), .O(gate33inter4));
  nand2 gate236(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate237(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate238(.a(N40), .O(gate33inter7));
  inv1  gate239(.a(N127), .O(gate33inter8));
  nand2 gate240(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate241(.a(s_11), .b(gate33inter3), .O(gate33inter10));
  nor2  gate242(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate243(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate244(.a(gate33inter12), .b(gate33inter1), .O(N186));

  xor2  gate441(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate442(.a(gate34inter0), .b(s_40), .O(gate34inter1));
  and2  gate443(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate444(.a(s_40), .O(gate34inter3));
  inv1  gate445(.a(s_41), .O(gate34inter4));
  nand2 gate446(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate447(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate448(.a(N47), .O(gate34inter7));
  inv1  gate449(.a(N131), .O(gate34inter8));
  nand2 gate450(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate451(.a(s_41), .b(gate34inter3), .O(gate34inter10));
  nor2  gate452(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate453(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate454(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate427(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate428(.a(gate35inter0), .b(s_38), .O(gate35inter1));
  and2  gate429(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate430(.a(s_38), .O(gate35inter3));
  inv1  gate431(.a(s_39), .O(gate35inter4));
  nand2 gate432(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate433(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate434(.a(N53), .O(gate35inter7));
  inv1  gate435(.a(N131), .O(gate35inter8));
  nand2 gate436(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate437(.a(s_39), .b(gate35inter3), .O(gate35inter10));
  nor2  gate438(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate439(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate440(.a(gate35inter12), .b(gate35inter1), .O(N188));

  xor2  gate217(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate218(.a(gate36inter0), .b(s_8), .O(gate36inter1));
  and2  gate219(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate220(.a(s_8), .O(gate36inter3));
  inv1  gate221(.a(s_9), .O(gate36inter4));
  nand2 gate222(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate223(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate224(.a(N60), .O(gate36inter7));
  inv1  gate225(.a(N135), .O(gate36inter8));
  nand2 gate226(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate227(.a(s_9), .b(gate36inter3), .O(gate36inter10));
  nor2  gate228(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate229(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate230(.a(gate36inter12), .b(gate36inter1), .O(N189));
nor2 gate37( .a(N66), .b(N135), .O(N190) );

  xor2  gate497(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate498(.a(gate38inter0), .b(s_48), .O(gate38inter1));
  and2  gate499(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate500(.a(s_48), .O(gate38inter3));
  inv1  gate501(.a(s_49), .O(gate38inter4));
  nand2 gate502(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate503(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate504(.a(N73), .O(gate38inter7));
  inv1  gate505(.a(N139), .O(gate38inter8));
  nand2 gate506(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate507(.a(s_49), .b(gate38inter3), .O(gate38inter10));
  nor2  gate508(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate509(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate510(.a(gate38inter12), .b(gate38inter1), .O(N191));

  xor2  gate315(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate316(.a(gate39inter0), .b(s_22), .O(gate39inter1));
  and2  gate317(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate318(.a(s_22), .O(gate39inter3));
  inv1  gate319(.a(s_23), .O(gate39inter4));
  nand2 gate320(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate321(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate322(.a(N79), .O(gate39inter7));
  inv1  gate323(.a(N139), .O(gate39inter8));
  nand2 gate324(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate325(.a(s_23), .b(gate39inter3), .O(gate39inter10));
  nor2  gate326(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate327(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate328(.a(gate39inter12), .b(gate39inter1), .O(N192));
nor2 gate40( .a(N86), .b(N143), .O(N193) );

  xor2  gate273(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate274(.a(gate41inter0), .b(s_16), .O(gate41inter1));
  and2  gate275(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate276(.a(s_16), .O(gate41inter3));
  inv1  gate277(.a(s_17), .O(gate41inter4));
  nand2 gate278(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate279(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate280(.a(N92), .O(gate41inter7));
  inv1  gate281(.a(N143), .O(gate41inter8));
  nand2 gate282(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate283(.a(s_17), .b(gate41inter3), .O(gate41inter10));
  nor2  gate284(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate285(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate286(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate203(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate204(.a(gate43inter0), .b(s_6), .O(gate43inter1));
  and2  gate205(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate206(.a(s_6), .O(gate43inter3));
  inv1  gate207(.a(s_7), .O(gate43inter4));
  nand2 gate208(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate209(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate210(.a(N105), .O(gate43inter7));
  inv1  gate211(.a(N147), .O(gate43inter8));
  nand2 gate212(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate213(.a(s_7), .b(gate43inter3), .O(gate43inter10));
  nor2  gate214(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate215(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate216(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate399(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate400(.a(gate50inter0), .b(s_34), .O(gate50inter1));
  and2  gate401(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate402(.a(s_34), .O(gate50inter3));
  inv1  gate403(.a(s_35), .O(gate50inter4));
  nand2 gate404(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate405(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate406(.a(N203), .O(gate50inter7));
  inv1  gate407(.a(N154), .O(gate50inter8));
  nand2 gate408(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate409(.a(s_35), .b(gate50inter3), .O(gate50inter10));
  nor2  gate410(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate411(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate412(.a(gate50inter12), .b(gate50inter1), .O(N224));

  xor2  gate623(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate624(.a(gate51inter0), .b(s_66), .O(gate51inter1));
  and2  gate625(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate626(.a(s_66), .O(gate51inter3));
  inv1  gate627(.a(s_67), .O(gate51inter4));
  nand2 gate628(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate629(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate630(.a(N203), .O(gate51inter7));
  inv1  gate631(.a(N159), .O(gate51inter8));
  nand2 gate632(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate633(.a(s_67), .b(gate51inter3), .O(gate51inter10));
  nor2  gate634(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate635(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate636(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );

  xor2  gate175(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate176(.a(gate54inter0), .b(s_2), .O(gate54inter1));
  and2  gate177(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate178(.a(s_2), .O(gate54inter3));
  inv1  gate179(.a(s_3), .O(gate54inter4));
  nand2 gate180(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate181(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate182(.a(N203), .O(gate54inter7));
  inv1  gate183(.a(N168), .O(gate54inter8));
  nand2 gate184(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate185(.a(s_3), .b(gate54inter3), .O(gate54inter10));
  nor2  gate186(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate187(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate188(.a(gate54inter12), .b(gate54inter1), .O(N236));
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate287(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate288(.a(gate59inter0), .b(s_18), .O(gate59inter1));
  and2  gate289(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate290(.a(s_18), .O(gate59inter3));
  inv1  gate291(.a(s_19), .O(gate59inter4));
  nand2 gate292(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate293(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate294(.a(N203), .O(gate59inter7));
  inv1  gate295(.a(N177), .O(gate59inter8));
  nand2 gate296(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate297(.a(s_19), .b(gate59inter3), .O(gate59inter10));
  nor2  gate298(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate299(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate300(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate259(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate260(.a(gate71inter0), .b(s_14), .O(gate71inter1));
  and2  gate261(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate262(.a(s_14), .O(gate71inter3));
  inv1  gate263(.a(s_15), .O(gate71inter4));
  nand2 gate264(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate265(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate266(.a(N230), .O(gate71inter7));
  inv1  gate267(.a(N185), .O(gate71inter8));
  nand2 gate268(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate269(.a(s_15), .b(gate71inter3), .O(gate71inter10));
  nor2  gate270(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate271(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate272(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate245(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate246(.a(gate73inter0), .b(s_12), .O(gate73inter1));
  and2  gate247(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate248(.a(s_12), .O(gate73inter3));
  inv1  gate249(.a(s_13), .O(gate73inter4));
  nand2 gate250(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate251(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate252(.a(N236), .O(gate73inter7));
  inv1  gate253(.a(N189), .O(gate73inter8));
  nand2 gate254(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate255(.a(s_13), .b(gate73inter3), .O(gate73inter10));
  nor2  gate256(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate257(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate258(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );

  xor2  gate189(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate190(.a(gate81inter0), .b(s_4), .O(gate81inter1));
  and2  gate191(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate192(.a(s_4), .O(gate81inter3));
  inv1  gate193(.a(s_5), .O(gate81inter4));
  nand2 gate194(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate195(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate196(.a(N236), .O(gate81inter7));
  inv1  gate197(.a(N190), .O(gate81inter8));
  nand2 gate198(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate199(.a(s_5), .b(gate81inter3), .O(gate81inter10));
  nor2  gate200(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate201(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate202(.a(gate81inter12), .b(gate81inter1), .O(N291));

  xor2  gate595(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate596(.a(gate82inter0), .b(s_62), .O(gate82inter1));
  and2  gate597(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate598(.a(s_62), .O(gate82inter3));
  inv1  gate599(.a(s_63), .O(gate82inter4));
  nand2 gate600(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate601(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate602(.a(N239), .O(gate82inter7));
  inv1  gate603(.a(N192), .O(gate82inter8));
  nand2 gate604(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate605(.a(s_63), .b(gate82inter3), .O(gate82inter10));
  nor2  gate606(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate607(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate608(.a(gate82inter12), .b(gate82inter1), .O(N292));
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate581(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate582(.a(gate99inter0), .b(s_60), .O(gate99inter1));
  and2  gate583(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate584(.a(s_60), .O(gate99inter3));
  inv1  gate585(.a(s_61), .O(gate99inter4));
  nand2 gate586(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate587(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate588(.a(N309), .O(gate99inter7));
  inv1  gate589(.a(N260), .O(gate99inter8));
  nand2 gate590(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate591(.a(s_61), .b(gate99inter3), .O(gate99inter10));
  nor2  gate592(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate593(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate594(.a(gate99inter12), .b(gate99inter1), .O(N330));

  xor2  gate329(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate330(.a(gate100inter0), .b(s_24), .O(gate100inter1));
  and2  gate331(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate332(.a(s_24), .O(gate100inter3));
  inv1  gate333(.a(s_25), .O(gate100inter4));
  nand2 gate334(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate335(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate336(.a(N309), .O(gate100inter7));
  inv1  gate337(.a(N264), .O(gate100inter8));
  nand2 gate338(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate339(.a(s_25), .b(gate100inter3), .O(gate100inter10));
  nor2  gate340(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate341(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate342(.a(gate100inter12), .b(gate100inter1), .O(N331));
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate539(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate540(.a(gate105inter0), .b(s_54), .O(gate105inter1));
  and2  gate541(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate542(.a(s_54), .O(gate105inter3));
  inv1  gate543(.a(s_55), .O(gate105inter4));
  nand2 gate544(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate545(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate546(.a(N319), .O(gate105inter7));
  inv1  gate547(.a(N21), .O(gate105inter8));
  nand2 gate548(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate549(.a(s_55), .b(gate105inter3), .O(gate105inter10));
  nor2  gate550(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate551(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate552(.a(gate105inter12), .b(gate105inter1), .O(N336));

  xor2  gate455(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate456(.a(gate106inter0), .b(s_42), .O(gate106inter1));
  and2  gate457(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate458(.a(s_42), .O(gate106inter3));
  inv1  gate459(.a(s_43), .O(gate106inter4));
  nand2 gate460(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate461(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate462(.a(N309), .O(gate106inter7));
  inv1  gate463(.a(N276), .O(gate106inter8));
  nand2 gate464(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate465(.a(s_43), .b(gate106inter3), .O(gate106inter10));
  nor2  gate466(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate467(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate468(.a(gate106inter12), .b(gate106inter1), .O(N337));

  xor2  gate371(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate372(.a(gate107inter0), .b(s_30), .O(gate107inter1));
  and2  gate373(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate374(.a(s_30), .O(gate107inter3));
  inv1  gate375(.a(s_31), .O(gate107inter4));
  nand2 gate376(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate377(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate378(.a(N319), .O(gate107inter7));
  inv1  gate379(.a(N34), .O(gate107inter8));
  nand2 gate380(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate381(.a(s_31), .b(gate107inter3), .O(gate107inter10));
  nor2  gate382(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate383(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate384(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate637(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate638(.a(gate111inter0), .b(s_68), .O(gate111inter1));
  and2  gate639(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate640(.a(s_68), .O(gate111inter3));
  inv1  gate641(.a(s_69), .O(gate111inter4));
  nand2 gate642(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate643(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate644(.a(N319), .O(gate111inter7));
  inv1  gate645(.a(N60), .O(gate111inter8));
  nand2 gate646(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate647(.a(s_69), .b(gate111inter3), .O(gate111inter10));
  nor2  gate648(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate649(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate650(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate301(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate302(.a(gate118inter0), .b(s_20), .O(gate118inter1));
  and2  gate303(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate304(.a(s_20), .O(gate118inter3));
  inv1  gate305(.a(s_21), .O(gate118inter4));
  nand2 gate306(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate307(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate308(.a(N331), .O(gate118inter7));
  inv1  gate309(.a(N301), .O(gate118inter8));
  nand2 gate310(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate311(.a(s_21), .b(gate118inter3), .O(gate118inter10));
  nor2  gate312(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate313(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate314(.a(gate118inter12), .b(gate118inter1), .O(N349));

  xor2  gate651(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate652(.a(gate119inter0), .b(s_70), .O(gate119inter1));
  and2  gate653(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate654(.a(s_70), .O(gate119inter3));
  inv1  gate655(.a(s_71), .O(gate119inter4));
  nand2 gate656(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate657(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate658(.a(N332), .O(gate119inter7));
  inv1  gate659(.a(N302), .O(gate119inter8));
  nand2 gate660(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate661(.a(s_71), .b(gate119inter3), .O(gate119inter10));
  nor2  gate662(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate663(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate664(.a(gate119inter12), .b(gate119inter1), .O(N350));
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate483(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate484(.a(gate121inter0), .b(s_46), .O(gate121inter1));
  and2  gate485(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate486(.a(s_46), .O(gate121inter3));
  inv1  gate487(.a(s_47), .O(gate121inter4));
  nand2 gate488(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate489(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate490(.a(N335), .O(gate121inter7));
  inv1  gate491(.a(N304), .O(gate121inter8));
  nand2 gate492(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate493(.a(s_47), .b(gate121inter3), .O(gate121inter10));
  nor2  gate494(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate495(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate496(.a(gate121inter12), .b(gate121inter1), .O(N352));
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate525(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate526(.a(gate132inter0), .b(s_52), .O(gate132inter1));
  and2  gate527(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate528(.a(s_52), .O(gate132inter3));
  inv1  gate529(.a(s_53), .O(gate132inter4));
  nand2 gate530(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate531(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate532(.a(N360), .O(gate132inter7));
  inv1  gate533(.a(N53), .O(gate132inter8));
  nand2 gate534(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate535(.a(s_53), .b(gate132inter3), .O(gate132inter10));
  nor2  gate536(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate537(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate538(.a(gate132inter12), .b(gate132inter1), .O(N374));

  xor2  gate553(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate554(.a(gate133inter0), .b(s_56), .O(gate133inter1));
  and2  gate555(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate556(.a(s_56), .O(gate133inter3));
  inv1  gate557(.a(s_57), .O(gate133inter4));
  nand2 gate558(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate559(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate560(.a(N360), .O(gate133inter7));
  inv1  gate561(.a(N66), .O(gate133inter8));
  nand2 gate562(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate563(.a(s_57), .b(gate133inter3), .O(gate133inter10));
  nor2  gate564(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate565(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate566(.a(gate133inter12), .b(gate133inter1), .O(N375));

  xor2  gate357(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate358(.a(gate134inter0), .b(s_28), .O(gate134inter1));
  and2  gate359(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate360(.a(s_28), .O(gate134inter3));
  inv1  gate361(.a(s_29), .O(gate134inter4));
  nand2 gate362(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate363(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate364(.a(N360), .O(gate134inter7));
  inv1  gate365(.a(N79), .O(gate134inter8));
  nand2 gate366(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate367(.a(s_29), .b(gate134inter3), .O(gate134inter10));
  nor2  gate368(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate369(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate370(.a(gate134inter12), .b(gate134inter1), .O(N376));
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate161(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate162(.a(gate153inter0), .b(s_0), .O(gate153inter1));
  and2  gate163(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate164(.a(s_0), .O(gate153inter3));
  inv1  gate165(.a(s_1), .O(gate153inter4));
  nand2 gate166(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate167(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate168(.a(N415), .O(gate153inter7));
  inv1  gate169(.a(N416), .O(gate153inter8));
  nand2 gate170(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate171(.a(s_1), .b(gate153inter3), .O(gate153inter10));
  nor2  gate172(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate173(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate174(.a(gate153inter12), .b(gate153inter1), .O(N421));
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule