module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1499(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1500(.a(gate9inter0), .b(s_136), .O(gate9inter1));
  and2  gate1501(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1502(.a(s_136), .O(gate9inter3));
  inv1  gate1503(.a(s_137), .O(gate9inter4));
  nand2 gate1504(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1505(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1506(.a(G1), .O(gate9inter7));
  inv1  gate1507(.a(G2), .O(gate9inter8));
  nand2 gate1508(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1509(.a(s_137), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1510(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1511(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1512(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate575(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate576(.a(gate12inter0), .b(s_4), .O(gate12inter1));
  and2  gate577(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate578(.a(s_4), .O(gate12inter3));
  inv1  gate579(.a(s_5), .O(gate12inter4));
  nand2 gate580(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate581(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate582(.a(G7), .O(gate12inter7));
  inv1  gate583(.a(G8), .O(gate12inter8));
  nand2 gate584(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate585(.a(s_5), .b(gate12inter3), .O(gate12inter10));
  nor2  gate586(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate587(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate588(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1737(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1738(.a(gate15inter0), .b(s_170), .O(gate15inter1));
  and2  gate1739(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1740(.a(s_170), .O(gate15inter3));
  inv1  gate1741(.a(s_171), .O(gate15inter4));
  nand2 gate1742(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1743(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1744(.a(G13), .O(gate15inter7));
  inv1  gate1745(.a(G14), .O(gate15inter8));
  nand2 gate1746(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1747(.a(s_171), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1748(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1749(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1750(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1121(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1122(.a(gate16inter0), .b(s_82), .O(gate16inter1));
  and2  gate1123(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1124(.a(s_82), .O(gate16inter3));
  inv1  gate1125(.a(s_83), .O(gate16inter4));
  nand2 gate1126(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1127(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1128(.a(G15), .O(gate16inter7));
  inv1  gate1129(.a(G16), .O(gate16inter8));
  nand2 gate1130(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1131(.a(s_83), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1132(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1133(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1134(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1177(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1178(.a(gate24inter0), .b(s_90), .O(gate24inter1));
  and2  gate1179(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1180(.a(s_90), .O(gate24inter3));
  inv1  gate1181(.a(s_91), .O(gate24inter4));
  nand2 gate1182(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1183(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1184(.a(G31), .O(gate24inter7));
  inv1  gate1185(.a(G32), .O(gate24inter8));
  nand2 gate1186(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1187(.a(s_91), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1188(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1189(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1190(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1261(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1262(.a(gate27inter0), .b(s_102), .O(gate27inter1));
  and2  gate1263(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1264(.a(s_102), .O(gate27inter3));
  inv1  gate1265(.a(s_103), .O(gate27inter4));
  nand2 gate1266(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1267(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1268(.a(G2), .O(gate27inter7));
  inv1  gate1269(.a(G6), .O(gate27inter8));
  nand2 gate1270(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1271(.a(s_103), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1272(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1273(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1274(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1583(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1584(.a(gate28inter0), .b(s_148), .O(gate28inter1));
  and2  gate1585(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1586(.a(s_148), .O(gate28inter3));
  inv1  gate1587(.a(s_149), .O(gate28inter4));
  nand2 gate1588(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1589(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1590(.a(G10), .O(gate28inter7));
  inv1  gate1591(.a(G14), .O(gate28inter8));
  nand2 gate1592(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1593(.a(s_149), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1594(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1595(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1596(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1191(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1192(.a(gate29inter0), .b(s_92), .O(gate29inter1));
  and2  gate1193(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1194(.a(s_92), .O(gate29inter3));
  inv1  gate1195(.a(s_93), .O(gate29inter4));
  nand2 gate1196(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1197(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1198(.a(G3), .O(gate29inter7));
  inv1  gate1199(.a(G7), .O(gate29inter8));
  nand2 gate1200(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1201(.a(s_93), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1202(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1203(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1204(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate911(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate912(.a(gate35inter0), .b(s_52), .O(gate35inter1));
  and2  gate913(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate914(.a(s_52), .O(gate35inter3));
  inv1  gate915(.a(s_53), .O(gate35inter4));
  nand2 gate916(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate917(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate918(.a(G18), .O(gate35inter7));
  inv1  gate919(.a(G22), .O(gate35inter8));
  nand2 gate920(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate921(.a(s_53), .b(gate35inter3), .O(gate35inter10));
  nor2  gate922(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate923(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate924(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1205(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1206(.a(gate39inter0), .b(s_94), .O(gate39inter1));
  and2  gate1207(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1208(.a(s_94), .O(gate39inter3));
  inv1  gate1209(.a(s_95), .O(gate39inter4));
  nand2 gate1210(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1211(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1212(.a(G20), .O(gate39inter7));
  inv1  gate1213(.a(G24), .O(gate39inter8));
  nand2 gate1214(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1215(.a(s_95), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1216(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1217(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1218(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1345(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1346(.a(gate41inter0), .b(s_114), .O(gate41inter1));
  and2  gate1347(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1348(.a(s_114), .O(gate41inter3));
  inv1  gate1349(.a(s_115), .O(gate41inter4));
  nand2 gate1350(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1351(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1352(.a(G1), .O(gate41inter7));
  inv1  gate1353(.a(G266), .O(gate41inter8));
  nand2 gate1354(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1355(.a(s_115), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1356(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1357(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1358(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate981(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate982(.a(gate45inter0), .b(s_62), .O(gate45inter1));
  and2  gate983(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate984(.a(s_62), .O(gate45inter3));
  inv1  gate985(.a(s_63), .O(gate45inter4));
  nand2 gate986(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate987(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate988(.a(G5), .O(gate45inter7));
  inv1  gate989(.a(G272), .O(gate45inter8));
  nand2 gate990(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate991(.a(s_63), .b(gate45inter3), .O(gate45inter10));
  nor2  gate992(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate993(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate994(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1751(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1752(.a(gate46inter0), .b(s_172), .O(gate46inter1));
  and2  gate1753(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1754(.a(s_172), .O(gate46inter3));
  inv1  gate1755(.a(s_173), .O(gate46inter4));
  nand2 gate1756(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1757(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1758(.a(G6), .O(gate46inter7));
  inv1  gate1759(.a(G272), .O(gate46inter8));
  nand2 gate1760(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1761(.a(s_173), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1762(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1763(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1764(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1821(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1822(.a(gate56inter0), .b(s_182), .O(gate56inter1));
  and2  gate1823(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1824(.a(s_182), .O(gate56inter3));
  inv1  gate1825(.a(s_183), .O(gate56inter4));
  nand2 gate1826(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1827(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1828(.a(G16), .O(gate56inter7));
  inv1  gate1829(.a(G287), .O(gate56inter8));
  nand2 gate1830(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1831(.a(s_183), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1832(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1833(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1834(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1415(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1416(.a(gate57inter0), .b(s_124), .O(gate57inter1));
  and2  gate1417(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1418(.a(s_124), .O(gate57inter3));
  inv1  gate1419(.a(s_125), .O(gate57inter4));
  nand2 gate1420(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1421(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1422(.a(G17), .O(gate57inter7));
  inv1  gate1423(.a(G290), .O(gate57inter8));
  nand2 gate1424(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1425(.a(s_125), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1426(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1427(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1428(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1079(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1080(.a(gate60inter0), .b(s_76), .O(gate60inter1));
  and2  gate1081(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1082(.a(s_76), .O(gate60inter3));
  inv1  gate1083(.a(s_77), .O(gate60inter4));
  nand2 gate1084(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1085(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1086(.a(G20), .O(gate60inter7));
  inv1  gate1087(.a(G293), .O(gate60inter8));
  nand2 gate1088(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1089(.a(s_77), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1090(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1091(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1092(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate967(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate968(.a(gate63inter0), .b(s_60), .O(gate63inter1));
  and2  gate969(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate970(.a(s_60), .O(gate63inter3));
  inv1  gate971(.a(s_61), .O(gate63inter4));
  nand2 gate972(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate973(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate974(.a(G23), .O(gate63inter7));
  inv1  gate975(.a(G299), .O(gate63inter8));
  nand2 gate976(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate977(.a(s_61), .b(gate63inter3), .O(gate63inter10));
  nor2  gate978(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate979(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate980(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1527(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1528(.a(gate68inter0), .b(s_140), .O(gate68inter1));
  and2  gate1529(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1530(.a(s_140), .O(gate68inter3));
  inv1  gate1531(.a(s_141), .O(gate68inter4));
  nand2 gate1532(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1533(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1534(.a(G28), .O(gate68inter7));
  inv1  gate1535(.a(G305), .O(gate68inter8));
  nand2 gate1536(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1537(.a(s_141), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1538(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1539(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1540(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate715(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate716(.a(gate70inter0), .b(s_24), .O(gate70inter1));
  and2  gate717(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate718(.a(s_24), .O(gate70inter3));
  inv1  gate719(.a(s_25), .O(gate70inter4));
  nand2 gate720(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate721(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate722(.a(G30), .O(gate70inter7));
  inv1  gate723(.a(G308), .O(gate70inter8));
  nand2 gate724(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate725(.a(s_25), .b(gate70inter3), .O(gate70inter10));
  nor2  gate726(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate727(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate728(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1219(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1220(.a(gate84inter0), .b(s_96), .O(gate84inter1));
  and2  gate1221(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1222(.a(s_96), .O(gate84inter3));
  inv1  gate1223(.a(s_97), .O(gate84inter4));
  nand2 gate1224(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1225(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1226(.a(G15), .O(gate84inter7));
  inv1  gate1227(.a(G329), .O(gate84inter8));
  nand2 gate1228(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1229(.a(s_97), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1230(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1231(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1232(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate939(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate940(.a(gate86inter0), .b(s_56), .O(gate86inter1));
  and2  gate941(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate942(.a(s_56), .O(gate86inter3));
  inv1  gate943(.a(s_57), .O(gate86inter4));
  nand2 gate944(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate945(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate946(.a(G8), .O(gate86inter7));
  inv1  gate947(.a(G332), .O(gate86inter8));
  nand2 gate948(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate949(.a(s_57), .b(gate86inter3), .O(gate86inter10));
  nor2  gate950(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate951(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate952(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1835(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1836(.a(gate87inter0), .b(s_184), .O(gate87inter1));
  and2  gate1837(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1838(.a(s_184), .O(gate87inter3));
  inv1  gate1839(.a(s_185), .O(gate87inter4));
  nand2 gate1840(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1841(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1842(.a(G12), .O(gate87inter7));
  inv1  gate1843(.a(G335), .O(gate87inter8));
  nand2 gate1844(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1845(.a(s_185), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1846(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1847(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1848(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1429(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1430(.a(gate92inter0), .b(s_126), .O(gate92inter1));
  and2  gate1431(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1432(.a(s_126), .O(gate92inter3));
  inv1  gate1433(.a(s_127), .O(gate92inter4));
  nand2 gate1434(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1435(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1436(.a(G29), .O(gate92inter7));
  inv1  gate1437(.a(G341), .O(gate92inter8));
  nand2 gate1438(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1439(.a(s_127), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1440(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1441(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1442(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1555(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1556(.a(gate95inter0), .b(s_144), .O(gate95inter1));
  and2  gate1557(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1558(.a(s_144), .O(gate95inter3));
  inv1  gate1559(.a(s_145), .O(gate95inter4));
  nand2 gate1560(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1561(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1562(.a(G26), .O(gate95inter7));
  inv1  gate1563(.a(G347), .O(gate95inter8));
  nand2 gate1564(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1565(.a(s_145), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1566(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1567(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1568(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1163(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1164(.a(gate98inter0), .b(s_88), .O(gate98inter1));
  and2  gate1165(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1166(.a(s_88), .O(gate98inter3));
  inv1  gate1167(.a(s_89), .O(gate98inter4));
  nand2 gate1168(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1169(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1170(.a(G23), .O(gate98inter7));
  inv1  gate1171(.a(G350), .O(gate98inter8));
  nand2 gate1172(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1173(.a(s_89), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1174(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1175(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1176(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1667(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1668(.a(gate105inter0), .b(s_160), .O(gate105inter1));
  and2  gate1669(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1670(.a(s_160), .O(gate105inter3));
  inv1  gate1671(.a(s_161), .O(gate105inter4));
  nand2 gate1672(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1673(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1674(.a(G362), .O(gate105inter7));
  inv1  gate1675(.a(G363), .O(gate105inter8));
  nand2 gate1676(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1677(.a(s_161), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1678(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1679(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1680(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1779(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1780(.a(gate116inter0), .b(s_176), .O(gate116inter1));
  and2  gate1781(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1782(.a(s_176), .O(gate116inter3));
  inv1  gate1783(.a(s_177), .O(gate116inter4));
  nand2 gate1784(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1785(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1786(.a(G384), .O(gate116inter7));
  inv1  gate1787(.a(G385), .O(gate116inter8));
  nand2 gate1788(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1789(.a(s_177), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1790(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1791(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1792(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate953(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate954(.a(gate119inter0), .b(s_58), .O(gate119inter1));
  and2  gate955(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate956(.a(s_58), .O(gate119inter3));
  inv1  gate957(.a(s_59), .O(gate119inter4));
  nand2 gate958(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate959(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate960(.a(G390), .O(gate119inter7));
  inv1  gate961(.a(G391), .O(gate119inter8));
  nand2 gate962(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate963(.a(s_59), .b(gate119inter3), .O(gate119inter10));
  nor2  gate964(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate965(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate966(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate785(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate786(.a(gate121inter0), .b(s_34), .O(gate121inter1));
  and2  gate787(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate788(.a(s_34), .O(gate121inter3));
  inv1  gate789(.a(s_35), .O(gate121inter4));
  nand2 gate790(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate791(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate792(.a(G394), .O(gate121inter7));
  inv1  gate793(.a(G395), .O(gate121inter8));
  nand2 gate794(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate795(.a(s_35), .b(gate121inter3), .O(gate121inter10));
  nor2  gate796(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate797(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate798(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1709(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1710(.a(gate126inter0), .b(s_166), .O(gate126inter1));
  and2  gate1711(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1712(.a(s_166), .O(gate126inter3));
  inv1  gate1713(.a(s_167), .O(gate126inter4));
  nand2 gate1714(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1715(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1716(.a(G404), .O(gate126inter7));
  inv1  gate1717(.a(G405), .O(gate126inter8));
  nand2 gate1718(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1719(.a(s_167), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1720(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1721(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1722(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate617(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate618(.a(gate133inter0), .b(s_10), .O(gate133inter1));
  and2  gate619(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate620(.a(s_10), .O(gate133inter3));
  inv1  gate621(.a(s_11), .O(gate133inter4));
  nand2 gate622(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate623(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate624(.a(G418), .O(gate133inter7));
  inv1  gate625(.a(G419), .O(gate133inter8));
  nand2 gate626(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate627(.a(s_11), .b(gate133inter3), .O(gate133inter10));
  nor2  gate628(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate629(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate630(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate645(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate646(.a(gate137inter0), .b(s_14), .O(gate137inter1));
  and2  gate647(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate648(.a(s_14), .O(gate137inter3));
  inv1  gate649(.a(s_15), .O(gate137inter4));
  nand2 gate650(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate651(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate652(.a(G426), .O(gate137inter7));
  inv1  gate653(.a(G429), .O(gate137inter8));
  nand2 gate654(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate655(.a(s_15), .b(gate137inter3), .O(gate137inter10));
  nor2  gate656(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate657(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate658(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate561(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate562(.a(gate141inter0), .b(s_2), .O(gate141inter1));
  and2  gate563(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate564(.a(s_2), .O(gate141inter3));
  inv1  gate565(.a(s_3), .O(gate141inter4));
  nand2 gate566(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate567(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate568(.a(G450), .O(gate141inter7));
  inv1  gate569(.a(G453), .O(gate141inter8));
  nand2 gate570(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate571(.a(s_3), .b(gate141inter3), .O(gate141inter10));
  nor2  gate572(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate573(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate574(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1807(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1808(.a(gate144inter0), .b(s_180), .O(gate144inter1));
  and2  gate1809(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1810(.a(s_180), .O(gate144inter3));
  inv1  gate1811(.a(s_181), .O(gate144inter4));
  nand2 gate1812(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1813(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1814(.a(G468), .O(gate144inter7));
  inv1  gate1815(.a(G471), .O(gate144inter8));
  nand2 gate1816(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1817(.a(s_181), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1818(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1819(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1820(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1401(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1402(.a(gate147inter0), .b(s_122), .O(gate147inter1));
  and2  gate1403(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1404(.a(s_122), .O(gate147inter3));
  inv1  gate1405(.a(s_123), .O(gate147inter4));
  nand2 gate1406(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1407(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1408(.a(G486), .O(gate147inter7));
  inv1  gate1409(.a(G489), .O(gate147inter8));
  nand2 gate1410(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1411(.a(s_123), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1412(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1413(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1414(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1443(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1444(.a(gate148inter0), .b(s_128), .O(gate148inter1));
  and2  gate1445(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1446(.a(s_128), .O(gate148inter3));
  inv1  gate1447(.a(s_129), .O(gate148inter4));
  nand2 gate1448(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1449(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1450(.a(G492), .O(gate148inter7));
  inv1  gate1451(.a(G495), .O(gate148inter8));
  nand2 gate1452(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1453(.a(s_129), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1454(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1455(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1456(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1289(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1290(.a(gate151inter0), .b(s_106), .O(gate151inter1));
  and2  gate1291(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1292(.a(s_106), .O(gate151inter3));
  inv1  gate1293(.a(s_107), .O(gate151inter4));
  nand2 gate1294(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1295(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1296(.a(G510), .O(gate151inter7));
  inv1  gate1297(.a(G513), .O(gate151inter8));
  nand2 gate1298(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1299(.a(s_107), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1300(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1301(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1302(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1275(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1276(.a(gate152inter0), .b(s_104), .O(gate152inter1));
  and2  gate1277(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1278(.a(s_104), .O(gate152inter3));
  inv1  gate1279(.a(s_105), .O(gate152inter4));
  nand2 gate1280(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1281(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1282(.a(G516), .O(gate152inter7));
  inv1  gate1283(.a(G519), .O(gate152inter8));
  nand2 gate1284(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1285(.a(s_105), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1286(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1287(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1288(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1765(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1766(.a(gate159inter0), .b(s_174), .O(gate159inter1));
  and2  gate1767(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1768(.a(s_174), .O(gate159inter3));
  inv1  gate1769(.a(s_175), .O(gate159inter4));
  nand2 gate1770(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1771(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1772(.a(G444), .O(gate159inter7));
  inv1  gate1773(.a(G531), .O(gate159inter8));
  nand2 gate1774(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1775(.a(s_175), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1776(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1777(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1778(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1625(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1626(.a(gate160inter0), .b(s_154), .O(gate160inter1));
  and2  gate1627(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1628(.a(s_154), .O(gate160inter3));
  inv1  gate1629(.a(s_155), .O(gate160inter4));
  nand2 gate1630(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1631(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1632(.a(G447), .O(gate160inter7));
  inv1  gate1633(.a(G531), .O(gate160inter8));
  nand2 gate1634(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1635(.a(s_155), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1636(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1637(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1638(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1485(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1486(.a(gate169inter0), .b(s_134), .O(gate169inter1));
  and2  gate1487(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1488(.a(s_134), .O(gate169inter3));
  inv1  gate1489(.a(s_135), .O(gate169inter4));
  nand2 gate1490(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1491(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1492(.a(G474), .O(gate169inter7));
  inv1  gate1493(.a(G546), .O(gate169inter8));
  nand2 gate1494(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1495(.a(s_135), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1496(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1497(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1498(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1009(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1010(.a(gate174inter0), .b(s_66), .O(gate174inter1));
  and2  gate1011(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1012(.a(s_66), .O(gate174inter3));
  inv1  gate1013(.a(s_67), .O(gate174inter4));
  nand2 gate1014(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1015(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1016(.a(G489), .O(gate174inter7));
  inv1  gate1017(.a(G552), .O(gate174inter8));
  nand2 gate1018(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1019(.a(s_67), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1020(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1021(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1022(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1065(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1066(.a(gate176inter0), .b(s_74), .O(gate176inter1));
  and2  gate1067(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1068(.a(s_74), .O(gate176inter3));
  inv1  gate1069(.a(s_75), .O(gate176inter4));
  nand2 gate1070(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1071(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1072(.a(G495), .O(gate176inter7));
  inv1  gate1073(.a(G555), .O(gate176inter8));
  nand2 gate1074(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1075(.a(s_75), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1076(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1077(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1078(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1387(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1388(.a(gate178inter0), .b(s_120), .O(gate178inter1));
  and2  gate1389(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1390(.a(s_120), .O(gate178inter3));
  inv1  gate1391(.a(s_121), .O(gate178inter4));
  nand2 gate1392(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1393(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1394(.a(G501), .O(gate178inter7));
  inv1  gate1395(.a(G558), .O(gate178inter8));
  nand2 gate1396(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1397(.a(s_121), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1398(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1399(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1400(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1947(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1948(.a(gate183inter0), .b(s_200), .O(gate183inter1));
  and2  gate1949(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1950(.a(s_200), .O(gate183inter3));
  inv1  gate1951(.a(s_201), .O(gate183inter4));
  nand2 gate1952(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1953(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1954(.a(G516), .O(gate183inter7));
  inv1  gate1955(.a(G567), .O(gate183inter8));
  nand2 gate1956(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1957(.a(s_201), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1958(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1959(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1960(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate855(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate856(.a(gate184inter0), .b(s_44), .O(gate184inter1));
  and2  gate857(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate858(.a(s_44), .O(gate184inter3));
  inv1  gate859(.a(s_45), .O(gate184inter4));
  nand2 gate860(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate861(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate862(.a(G519), .O(gate184inter7));
  inv1  gate863(.a(G567), .O(gate184inter8));
  nand2 gate864(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate865(.a(s_45), .b(gate184inter3), .O(gate184inter10));
  nor2  gate866(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate867(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate868(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate995(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate996(.a(gate192inter0), .b(s_64), .O(gate192inter1));
  and2  gate997(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate998(.a(s_64), .O(gate192inter3));
  inv1  gate999(.a(s_65), .O(gate192inter4));
  nand2 gate1000(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1001(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1002(.a(G584), .O(gate192inter7));
  inv1  gate1003(.a(G585), .O(gate192inter8));
  nand2 gate1004(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1005(.a(s_65), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1006(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1007(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1008(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1919(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1920(.a(gate194inter0), .b(s_196), .O(gate194inter1));
  and2  gate1921(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1922(.a(s_196), .O(gate194inter3));
  inv1  gate1923(.a(s_197), .O(gate194inter4));
  nand2 gate1924(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1925(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1926(.a(G588), .O(gate194inter7));
  inv1  gate1927(.a(G589), .O(gate194inter8));
  nand2 gate1928(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1929(.a(s_197), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1930(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1931(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1932(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate729(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate730(.a(gate196inter0), .b(s_26), .O(gate196inter1));
  and2  gate731(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate732(.a(s_26), .O(gate196inter3));
  inv1  gate733(.a(s_27), .O(gate196inter4));
  nand2 gate734(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate735(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate736(.a(G592), .O(gate196inter7));
  inv1  gate737(.a(G593), .O(gate196inter8));
  nand2 gate738(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate739(.a(s_27), .b(gate196inter3), .O(gate196inter10));
  nor2  gate740(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate741(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate742(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1863(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1864(.a(gate198inter0), .b(s_188), .O(gate198inter1));
  and2  gate1865(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1866(.a(s_188), .O(gate198inter3));
  inv1  gate1867(.a(s_189), .O(gate198inter4));
  nand2 gate1868(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1869(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1870(.a(G596), .O(gate198inter7));
  inv1  gate1871(.a(G597), .O(gate198inter8));
  nand2 gate1872(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1873(.a(s_189), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1874(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1875(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1876(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1905(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1906(.a(gate201inter0), .b(s_194), .O(gate201inter1));
  and2  gate1907(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1908(.a(s_194), .O(gate201inter3));
  inv1  gate1909(.a(s_195), .O(gate201inter4));
  nand2 gate1910(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1911(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1912(.a(G602), .O(gate201inter7));
  inv1  gate1913(.a(G607), .O(gate201inter8));
  nand2 gate1914(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1915(.a(s_195), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1916(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1917(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1918(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1037(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1038(.a(gate205inter0), .b(s_70), .O(gate205inter1));
  and2  gate1039(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1040(.a(s_70), .O(gate205inter3));
  inv1  gate1041(.a(s_71), .O(gate205inter4));
  nand2 gate1042(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1043(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1044(.a(G622), .O(gate205inter7));
  inv1  gate1045(.a(G627), .O(gate205inter8));
  nand2 gate1046(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1047(.a(s_71), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1048(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1049(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1050(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1597(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1598(.a(gate206inter0), .b(s_150), .O(gate206inter1));
  and2  gate1599(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1600(.a(s_150), .O(gate206inter3));
  inv1  gate1601(.a(s_151), .O(gate206inter4));
  nand2 gate1602(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1603(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1604(.a(G632), .O(gate206inter7));
  inv1  gate1605(.a(G637), .O(gate206inter8));
  nand2 gate1606(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1607(.a(s_151), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1608(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1609(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1610(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate897(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate898(.a(gate209inter0), .b(s_50), .O(gate209inter1));
  and2  gate899(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate900(.a(s_50), .O(gate209inter3));
  inv1  gate901(.a(s_51), .O(gate209inter4));
  nand2 gate902(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate903(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate904(.a(G602), .O(gate209inter7));
  inv1  gate905(.a(G666), .O(gate209inter8));
  nand2 gate906(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate907(.a(s_51), .b(gate209inter3), .O(gate209inter10));
  nor2  gate908(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate909(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate910(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1793(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1794(.a(gate210inter0), .b(s_178), .O(gate210inter1));
  and2  gate1795(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1796(.a(s_178), .O(gate210inter3));
  inv1  gate1797(.a(s_179), .O(gate210inter4));
  nand2 gate1798(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1799(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1800(.a(G607), .O(gate210inter7));
  inv1  gate1801(.a(G666), .O(gate210inter8));
  nand2 gate1802(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1803(.a(s_179), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1804(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1805(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1806(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate701(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate702(.a(gate214inter0), .b(s_22), .O(gate214inter1));
  and2  gate703(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate704(.a(s_22), .O(gate214inter3));
  inv1  gate705(.a(s_23), .O(gate214inter4));
  nand2 gate706(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate707(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate708(.a(G612), .O(gate214inter7));
  inv1  gate709(.a(G672), .O(gate214inter8));
  nand2 gate710(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate711(.a(s_23), .b(gate214inter3), .O(gate214inter10));
  nor2  gate712(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate713(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate714(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate813(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate814(.a(gate215inter0), .b(s_38), .O(gate215inter1));
  and2  gate815(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate816(.a(s_38), .O(gate215inter3));
  inv1  gate817(.a(s_39), .O(gate215inter4));
  nand2 gate818(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate819(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate820(.a(G607), .O(gate215inter7));
  inv1  gate821(.a(G675), .O(gate215inter8));
  nand2 gate822(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate823(.a(s_39), .b(gate215inter3), .O(gate215inter10));
  nor2  gate824(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate825(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate826(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1247(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1248(.a(gate216inter0), .b(s_100), .O(gate216inter1));
  and2  gate1249(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1250(.a(s_100), .O(gate216inter3));
  inv1  gate1251(.a(s_101), .O(gate216inter4));
  nand2 gate1252(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1253(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1254(.a(G617), .O(gate216inter7));
  inv1  gate1255(.a(G675), .O(gate216inter8));
  nand2 gate1256(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1257(.a(s_101), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1258(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1259(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1260(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate883(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate884(.a(gate218inter0), .b(s_48), .O(gate218inter1));
  and2  gate885(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate886(.a(s_48), .O(gate218inter3));
  inv1  gate887(.a(s_49), .O(gate218inter4));
  nand2 gate888(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate889(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate890(.a(G627), .O(gate218inter7));
  inv1  gate891(.a(G678), .O(gate218inter8));
  nand2 gate892(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate893(.a(s_49), .b(gate218inter3), .O(gate218inter10));
  nor2  gate894(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate895(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate896(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1457(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1458(.a(gate219inter0), .b(s_130), .O(gate219inter1));
  and2  gate1459(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1460(.a(s_130), .O(gate219inter3));
  inv1  gate1461(.a(s_131), .O(gate219inter4));
  nand2 gate1462(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1463(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1464(.a(G632), .O(gate219inter7));
  inv1  gate1465(.a(G681), .O(gate219inter8));
  nand2 gate1466(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1467(.a(s_131), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1468(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1469(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1470(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1933(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1934(.a(gate222inter0), .b(s_198), .O(gate222inter1));
  and2  gate1935(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1936(.a(s_198), .O(gate222inter3));
  inv1  gate1937(.a(s_199), .O(gate222inter4));
  nand2 gate1938(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1939(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1940(.a(G632), .O(gate222inter7));
  inv1  gate1941(.a(G684), .O(gate222inter8));
  nand2 gate1942(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1943(.a(s_199), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1944(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1945(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1946(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate869(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate870(.a(gate223inter0), .b(s_46), .O(gate223inter1));
  and2  gate871(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate872(.a(s_46), .O(gate223inter3));
  inv1  gate873(.a(s_47), .O(gate223inter4));
  nand2 gate874(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate875(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate876(.a(G627), .O(gate223inter7));
  inv1  gate877(.a(G687), .O(gate223inter8));
  nand2 gate878(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate879(.a(s_47), .b(gate223inter3), .O(gate223inter10));
  nor2  gate880(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate881(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate882(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1373(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1374(.a(gate236inter0), .b(s_118), .O(gate236inter1));
  and2  gate1375(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1376(.a(s_118), .O(gate236inter3));
  inv1  gate1377(.a(s_119), .O(gate236inter4));
  nand2 gate1378(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1379(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1380(.a(G251), .O(gate236inter7));
  inv1  gate1381(.a(G727), .O(gate236inter8));
  nand2 gate1382(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1383(.a(s_119), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1384(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1385(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1386(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate771(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate772(.a(gate237inter0), .b(s_32), .O(gate237inter1));
  and2  gate773(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate774(.a(s_32), .O(gate237inter3));
  inv1  gate775(.a(s_33), .O(gate237inter4));
  nand2 gate776(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate777(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate778(.a(G254), .O(gate237inter7));
  inv1  gate779(.a(G706), .O(gate237inter8));
  nand2 gate780(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate781(.a(s_33), .b(gate237inter3), .O(gate237inter10));
  nor2  gate782(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate783(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate784(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1681(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1682(.a(gate241inter0), .b(s_162), .O(gate241inter1));
  and2  gate1683(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1684(.a(s_162), .O(gate241inter3));
  inv1  gate1685(.a(s_163), .O(gate241inter4));
  nand2 gate1686(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1687(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1688(.a(G242), .O(gate241inter7));
  inv1  gate1689(.a(G730), .O(gate241inter8));
  nand2 gate1690(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1691(.a(s_163), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1692(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1693(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1694(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1653(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1654(.a(gate244inter0), .b(s_158), .O(gate244inter1));
  and2  gate1655(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1656(.a(s_158), .O(gate244inter3));
  inv1  gate1657(.a(s_159), .O(gate244inter4));
  nand2 gate1658(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1659(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1660(.a(G721), .O(gate244inter7));
  inv1  gate1661(.a(G733), .O(gate244inter8));
  nand2 gate1662(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1663(.a(s_159), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1664(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1665(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1666(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate925(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate926(.a(gate246inter0), .b(s_54), .O(gate246inter1));
  and2  gate927(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate928(.a(s_54), .O(gate246inter3));
  inv1  gate929(.a(s_55), .O(gate246inter4));
  nand2 gate930(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate931(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate932(.a(G724), .O(gate246inter7));
  inv1  gate933(.a(G736), .O(gate246inter8));
  nand2 gate934(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate935(.a(s_55), .b(gate246inter3), .O(gate246inter10));
  nor2  gate936(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate937(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate938(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1513(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1514(.a(gate250inter0), .b(s_138), .O(gate250inter1));
  and2  gate1515(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1516(.a(s_138), .O(gate250inter3));
  inv1  gate1517(.a(s_139), .O(gate250inter4));
  nand2 gate1518(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1519(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1520(.a(G706), .O(gate250inter7));
  inv1  gate1521(.a(G742), .O(gate250inter8));
  nand2 gate1522(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1523(.a(s_139), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1524(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1525(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1526(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1569(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1570(.a(gate268inter0), .b(s_146), .O(gate268inter1));
  and2  gate1571(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1572(.a(s_146), .O(gate268inter3));
  inv1  gate1573(.a(s_147), .O(gate268inter4));
  nand2 gate1574(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1575(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1576(.a(G651), .O(gate268inter7));
  inv1  gate1577(.a(G779), .O(gate268inter8));
  nand2 gate1578(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1579(.a(s_147), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1580(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1581(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1582(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1107(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1108(.a(gate269inter0), .b(s_80), .O(gate269inter1));
  and2  gate1109(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1110(.a(s_80), .O(gate269inter3));
  inv1  gate1111(.a(s_81), .O(gate269inter4));
  nand2 gate1112(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1113(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1114(.a(G654), .O(gate269inter7));
  inv1  gate1115(.a(G782), .O(gate269inter8));
  nand2 gate1116(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1117(.a(s_81), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1118(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1119(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1120(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1023(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1024(.a(gate275inter0), .b(s_68), .O(gate275inter1));
  and2  gate1025(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1026(.a(s_68), .O(gate275inter3));
  inv1  gate1027(.a(s_69), .O(gate275inter4));
  nand2 gate1028(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1029(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1030(.a(G645), .O(gate275inter7));
  inv1  gate1031(.a(G797), .O(gate275inter8));
  nand2 gate1032(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1033(.a(s_69), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1034(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1035(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1036(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate687(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate688(.a(gate276inter0), .b(s_20), .O(gate276inter1));
  and2  gate689(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate690(.a(s_20), .O(gate276inter3));
  inv1  gate691(.a(s_21), .O(gate276inter4));
  nand2 gate692(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate693(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate694(.a(G773), .O(gate276inter7));
  inv1  gate695(.a(G797), .O(gate276inter8));
  nand2 gate696(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate697(.a(s_21), .b(gate276inter3), .O(gate276inter10));
  nor2  gate698(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate699(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate700(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1471(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1472(.a(gate279inter0), .b(s_132), .O(gate279inter1));
  and2  gate1473(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1474(.a(s_132), .O(gate279inter3));
  inv1  gate1475(.a(s_133), .O(gate279inter4));
  nand2 gate1476(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1477(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1478(.a(G651), .O(gate279inter7));
  inv1  gate1479(.a(G803), .O(gate279inter8));
  nand2 gate1480(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1481(.a(s_133), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1482(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1483(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1484(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate631(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate632(.a(gate288inter0), .b(s_12), .O(gate288inter1));
  and2  gate633(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate634(.a(s_12), .O(gate288inter3));
  inv1  gate635(.a(s_13), .O(gate288inter4));
  nand2 gate636(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate637(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate638(.a(G791), .O(gate288inter7));
  inv1  gate639(.a(G815), .O(gate288inter8));
  nand2 gate640(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate641(.a(s_13), .b(gate288inter3), .O(gate288inter10));
  nor2  gate642(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate643(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate644(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate799(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate800(.a(gate294inter0), .b(s_36), .O(gate294inter1));
  and2  gate801(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate802(.a(s_36), .O(gate294inter3));
  inv1  gate803(.a(s_37), .O(gate294inter4));
  nand2 gate804(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate805(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate806(.a(G832), .O(gate294inter7));
  inv1  gate807(.a(G833), .O(gate294inter8));
  nand2 gate808(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate809(.a(s_37), .b(gate294inter3), .O(gate294inter10));
  nor2  gate810(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate811(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate812(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1233(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1234(.a(gate295inter0), .b(s_98), .O(gate295inter1));
  and2  gate1235(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1236(.a(s_98), .O(gate295inter3));
  inv1  gate1237(.a(s_99), .O(gate295inter4));
  nand2 gate1238(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1239(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1240(.a(G830), .O(gate295inter7));
  inv1  gate1241(.a(G831), .O(gate295inter8));
  nand2 gate1242(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1243(.a(s_99), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1244(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1245(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1246(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate841(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate842(.a(gate399inter0), .b(s_42), .O(gate399inter1));
  and2  gate843(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate844(.a(s_42), .O(gate399inter3));
  inv1  gate845(.a(s_43), .O(gate399inter4));
  nand2 gate846(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate847(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate848(.a(G13), .O(gate399inter7));
  inv1  gate849(.a(G1072), .O(gate399inter8));
  nand2 gate850(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate851(.a(s_43), .b(gate399inter3), .O(gate399inter10));
  nor2  gate852(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate853(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate854(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate547(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate548(.a(gate409inter0), .b(s_0), .O(gate409inter1));
  and2  gate549(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate550(.a(s_0), .O(gate409inter3));
  inv1  gate551(.a(s_1), .O(gate409inter4));
  nand2 gate552(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate553(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate554(.a(G23), .O(gate409inter7));
  inv1  gate555(.a(G1102), .O(gate409inter8));
  nand2 gate556(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate557(.a(s_1), .b(gate409inter3), .O(gate409inter10));
  nor2  gate558(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate559(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate560(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1891(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1892(.a(gate417inter0), .b(s_192), .O(gate417inter1));
  and2  gate1893(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1894(.a(s_192), .O(gate417inter3));
  inv1  gate1895(.a(s_193), .O(gate417inter4));
  nand2 gate1896(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1897(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1898(.a(G31), .O(gate417inter7));
  inv1  gate1899(.a(G1126), .O(gate417inter8));
  nand2 gate1900(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1901(.a(s_193), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1902(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1903(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1904(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1877(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1878(.a(gate419inter0), .b(s_190), .O(gate419inter1));
  and2  gate1879(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1880(.a(s_190), .O(gate419inter3));
  inv1  gate1881(.a(s_191), .O(gate419inter4));
  nand2 gate1882(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1883(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1884(.a(G1), .O(gate419inter7));
  inv1  gate1885(.a(G1132), .O(gate419inter8));
  nand2 gate1886(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1887(.a(s_191), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1888(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1889(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1890(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1051(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1052(.a(gate420inter0), .b(s_72), .O(gate420inter1));
  and2  gate1053(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1054(.a(s_72), .O(gate420inter3));
  inv1  gate1055(.a(s_73), .O(gate420inter4));
  nand2 gate1056(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1057(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1058(.a(G1036), .O(gate420inter7));
  inv1  gate1059(.a(G1132), .O(gate420inter8));
  nand2 gate1060(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1061(.a(s_73), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1062(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1063(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1064(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1331(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1332(.a(gate422inter0), .b(s_112), .O(gate422inter1));
  and2  gate1333(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1334(.a(s_112), .O(gate422inter3));
  inv1  gate1335(.a(s_113), .O(gate422inter4));
  nand2 gate1336(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1337(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1338(.a(G1039), .O(gate422inter7));
  inv1  gate1339(.a(G1135), .O(gate422inter8));
  nand2 gate1340(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1341(.a(s_113), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1342(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1343(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1344(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate757(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate758(.a(gate424inter0), .b(s_30), .O(gate424inter1));
  and2  gate759(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate760(.a(s_30), .O(gate424inter3));
  inv1  gate761(.a(s_31), .O(gate424inter4));
  nand2 gate762(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate763(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate764(.a(G1042), .O(gate424inter7));
  inv1  gate765(.a(G1138), .O(gate424inter8));
  nand2 gate766(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate767(.a(s_31), .b(gate424inter3), .O(gate424inter10));
  nor2  gate768(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate769(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate770(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate673(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate674(.a(gate433inter0), .b(s_18), .O(gate433inter1));
  and2  gate675(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate676(.a(s_18), .O(gate433inter3));
  inv1  gate677(.a(s_19), .O(gate433inter4));
  nand2 gate678(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate679(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate680(.a(G8), .O(gate433inter7));
  inv1  gate681(.a(G1153), .O(gate433inter8));
  nand2 gate682(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate683(.a(s_19), .b(gate433inter3), .O(gate433inter10));
  nor2  gate684(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate685(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate686(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1723(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1724(.a(gate450inter0), .b(s_168), .O(gate450inter1));
  and2  gate1725(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1726(.a(s_168), .O(gate450inter3));
  inv1  gate1727(.a(s_169), .O(gate450inter4));
  nand2 gate1728(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1729(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1730(.a(G1081), .O(gate450inter7));
  inv1  gate1731(.a(G1177), .O(gate450inter8));
  nand2 gate1732(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1733(.a(s_169), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1734(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1735(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1736(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate603(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate604(.a(gate451inter0), .b(s_8), .O(gate451inter1));
  and2  gate605(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate606(.a(s_8), .O(gate451inter3));
  inv1  gate607(.a(s_9), .O(gate451inter4));
  nand2 gate608(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate609(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate610(.a(G17), .O(gate451inter7));
  inv1  gate611(.a(G1180), .O(gate451inter8));
  nand2 gate612(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate613(.a(s_9), .b(gate451inter3), .O(gate451inter10));
  nor2  gate614(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate615(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate616(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1639(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1640(.a(gate457inter0), .b(s_156), .O(gate457inter1));
  and2  gate1641(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1642(.a(s_156), .O(gate457inter3));
  inv1  gate1643(.a(s_157), .O(gate457inter4));
  nand2 gate1644(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1645(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1646(.a(G20), .O(gate457inter7));
  inv1  gate1647(.a(G1189), .O(gate457inter8));
  nand2 gate1648(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1649(.a(s_157), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1650(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1651(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1652(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1849(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1850(.a(gate465inter0), .b(s_186), .O(gate465inter1));
  and2  gate1851(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1852(.a(s_186), .O(gate465inter3));
  inv1  gate1853(.a(s_187), .O(gate465inter4));
  nand2 gate1854(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1855(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1856(.a(G24), .O(gate465inter7));
  inv1  gate1857(.a(G1201), .O(gate465inter8));
  nand2 gate1858(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1859(.a(s_187), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1860(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1861(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1862(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1149(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1150(.a(gate466inter0), .b(s_86), .O(gate466inter1));
  and2  gate1151(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1152(.a(s_86), .O(gate466inter3));
  inv1  gate1153(.a(s_87), .O(gate466inter4));
  nand2 gate1154(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1155(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1156(.a(G1105), .O(gate466inter7));
  inv1  gate1157(.a(G1201), .O(gate466inter8));
  nand2 gate1158(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1159(.a(s_87), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1160(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1161(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1162(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1093(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1094(.a(gate469inter0), .b(s_78), .O(gate469inter1));
  and2  gate1095(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1096(.a(s_78), .O(gate469inter3));
  inv1  gate1097(.a(s_79), .O(gate469inter4));
  nand2 gate1098(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1099(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1100(.a(G26), .O(gate469inter7));
  inv1  gate1101(.a(G1207), .O(gate469inter8));
  nand2 gate1102(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1103(.a(s_79), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1104(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1105(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1106(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1303(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1304(.a(gate476inter0), .b(s_108), .O(gate476inter1));
  and2  gate1305(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1306(.a(s_108), .O(gate476inter3));
  inv1  gate1307(.a(s_109), .O(gate476inter4));
  nand2 gate1308(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1309(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1310(.a(G1120), .O(gate476inter7));
  inv1  gate1311(.a(G1216), .O(gate476inter8));
  nand2 gate1312(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1313(.a(s_109), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1314(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1315(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1316(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1317(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1318(.a(gate480inter0), .b(s_110), .O(gate480inter1));
  and2  gate1319(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1320(.a(s_110), .O(gate480inter3));
  inv1  gate1321(.a(s_111), .O(gate480inter4));
  nand2 gate1322(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1323(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1324(.a(G1126), .O(gate480inter7));
  inv1  gate1325(.a(G1222), .O(gate480inter8));
  nand2 gate1326(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1327(.a(s_111), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1328(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1329(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1330(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1359(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1360(.a(gate484inter0), .b(s_116), .O(gate484inter1));
  and2  gate1361(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1362(.a(s_116), .O(gate484inter3));
  inv1  gate1363(.a(s_117), .O(gate484inter4));
  nand2 gate1364(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1365(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1366(.a(G1230), .O(gate484inter7));
  inv1  gate1367(.a(G1231), .O(gate484inter8));
  nand2 gate1368(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1369(.a(s_117), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1370(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1371(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1372(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate743(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate744(.a(gate488inter0), .b(s_28), .O(gate488inter1));
  and2  gate745(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate746(.a(s_28), .O(gate488inter3));
  inv1  gate747(.a(s_29), .O(gate488inter4));
  nand2 gate748(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate749(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate750(.a(G1238), .O(gate488inter7));
  inv1  gate751(.a(G1239), .O(gate488inter8));
  nand2 gate752(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate753(.a(s_29), .b(gate488inter3), .O(gate488inter10));
  nor2  gate754(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate755(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate756(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate659(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate660(.a(gate491inter0), .b(s_16), .O(gate491inter1));
  and2  gate661(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate662(.a(s_16), .O(gate491inter3));
  inv1  gate663(.a(s_17), .O(gate491inter4));
  nand2 gate664(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate665(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate666(.a(G1244), .O(gate491inter7));
  inv1  gate667(.a(G1245), .O(gate491inter8));
  nand2 gate668(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate669(.a(s_17), .b(gate491inter3), .O(gate491inter10));
  nor2  gate670(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate671(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate672(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1135(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1136(.a(gate494inter0), .b(s_84), .O(gate494inter1));
  and2  gate1137(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1138(.a(s_84), .O(gate494inter3));
  inv1  gate1139(.a(s_85), .O(gate494inter4));
  nand2 gate1140(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1141(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1142(.a(G1250), .O(gate494inter7));
  inv1  gate1143(.a(G1251), .O(gate494inter8));
  nand2 gate1144(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1145(.a(s_85), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1146(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1147(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1148(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate589(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate590(.a(gate496inter0), .b(s_6), .O(gate496inter1));
  and2  gate591(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate592(.a(s_6), .O(gate496inter3));
  inv1  gate593(.a(s_7), .O(gate496inter4));
  nand2 gate594(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate595(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate596(.a(G1254), .O(gate496inter7));
  inv1  gate597(.a(G1255), .O(gate496inter8));
  nand2 gate598(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate599(.a(s_7), .b(gate496inter3), .O(gate496inter10));
  nor2  gate600(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate601(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate602(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1541(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1542(.a(gate499inter0), .b(s_142), .O(gate499inter1));
  and2  gate1543(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1544(.a(s_142), .O(gate499inter3));
  inv1  gate1545(.a(s_143), .O(gate499inter4));
  nand2 gate1546(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1547(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1548(.a(G1260), .O(gate499inter7));
  inv1  gate1549(.a(G1261), .O(gate499inter8));
  nand2 gate1550(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1551(.a(s_143), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1552(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1553(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1554(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1695(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1696(.a(gate501inter0), .b(s_164), .O(gate501inter1));
  and2  gate1697(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1698(.a(s_164), .O(gate501inter3));
  inv1  gate1699(.a(s_165), .O(gate501inter4));
  nand2 gate1700(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1701(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1702(.a(G1264), .O(gate501inter7));
  inv1  gate1703(.a(G1265), .O(gate501inter8));
  nand2 gate1704(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1705(.a(s_165), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1706(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1707(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1708(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate827(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate828(.a(gate504inter0), .b(s_40), .O(gate504inter1));
  and2  gate829(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate830(.a(s_40), .O(gate504inter3));
  inv1  gate831(.a(s_41), .O(gate504inter4));
  nand2 gate832(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate833(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate834(.a(G1270), .O(gate504inter7));
  inv1  gate835(.a(G1271), .O(gate504inter8));
  nand2 gate836(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate837(.a(s_41), .b(gate504inter3), .O(gate504inter10));
  nor2  gate838(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate839(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate840(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1611(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1612(.a(gate508inter0), .b(s_152), .O(gate508inter1));
  and2  gate1613(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1614(.a(s_152), .O(gate508inter3));
  inv1  gate1615(.a(s_153), .O(gate508inter4));
  nand2 gate1616(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1617(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1618(.a(G1278), .O(gate508inter7));
  inv1  gate1619(.a(G1279), .O(gate508inter8));
  nand2 gate1620(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1621(.a(s_153), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1622(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1623(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1624(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule