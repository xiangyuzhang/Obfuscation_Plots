module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate413(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate414(.a(gate6inter0), .b(s_30), .O(gate6inter1));
  and2  gate415(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate416(.a(s_30), .O(gate6inter3));
  inv1  gate417(.a(s_31), .O(gate6inter4));
  nand2 gate418(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate419(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate420(.a(N41), .O(gate6inter7));
  inv1  gate421(.a(N45), .O(gate6inter8));
  nand2 gate422(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate423(.a(s_31), .b(gate6inter3), .O(gate6inter10));
  nor2  gate424(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate425(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate426(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate287(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate288(.a(gate8inter0), .b(s_12), .O(gate8inter1));
  and2  gate289(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate290(.a(s_12), .O(gate8inter3));
  inv1  gate291(.a(s_13), .O(gate8inter4));
  nand2 gate292(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate293(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate294(.a(N57), .O(gate8inter7));
  inv1  gate295(.a(N61), .O(gate8inter8));
  nand2 gate296(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate297(.a(s_13), .b(gate8inter3), .O(gate8inter10));
  nor2  gate298(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate299(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate300(.a(gate8inter12), .b(gate8inter1), .O(N257));
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );

  xor2  gate329(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate330(.a(gate15inter0), .b(s_18), .O(gate15inter1));
  and2  gate331(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate332(.a(s_18), .O(gate15inter3));
  inv1  gate333(.a(s_19), .O(gate15inter4));
  nand2 gate334(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate335(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate336(.a(N113), .O(gate15inter7));
  inv1  gate337(.a(N117), .O(gate15inter8));
  nand2 gate338(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate339(.a(s_19), .b(gate15inter3), .O(gate15inter10));
  nor2  gate340(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate341(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate342(.a(gate15inter12), .b(gate15inter1), .O(N264));
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );

  xor2  gate259(.a(N251), .b(N250), .O(gate41inter0));
  nand2 gate260(.a(gate41inter0), .b(s_8), .O(gate41inter1));
  and2  gate261(.a(N251), .b(N250), .O(gate41inter2));
  inv1  gate262(.a(s_8), .O(gate41inter3));
  inv1  gate263(.a(s_9), .O(gate41inter4));
  nand2 gate264(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate265(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate266(.a(N250), .O(gate41inter7));
  inv1  gate267(.a(N251), .O(gate41inter8));
  nand2 gate268(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate269(.a(s_9), .b(gate41inter3), .O(gate41inter10));
  nor2  gate270(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate271(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate272(.a(gate41inter12), .b(gate41inter1), .O(N290));
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );

  xor2  gate203(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate204(.a(gate48inter0), .b(s_0), .O(gate48inter1));
  and2  gate205(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate206(.a(s_0), .O(gate48inter3));
  inv1  gate207(.a(s_1), .O(gate48inter4));
  nand2 gate208(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate209(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate210(.a(N264), .O(gate48inter7));
  inv1  gate211(.a(N265), .O(gate48inter8));
  nand2 gate212(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate213(.a(s_1), .b(gate48inter3), .O(gate48inter10));
  nor2  gate214(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate215(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate216(.a(gate48inter12), .b(gate48inter1), .O(N311));
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );

  xor2  gate217(.a(N311), .b(N305), .O(gate64inter0));
  nand2 gate218(.a(gate64inter0), .b(s_2), .O(gate64inter1));
  and2  gate219(.a(N311), .b(N305), .O(gate64inter2));
  inv1  gate220(.a(s_2), .O(gate64inter3));
  inv1  gate221(.a(s_3), .O(gate64inter4));
  nand2 gate222(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate223(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate224(.a(N305), .O(gate64inter7));
  inv1  gate225(.a(N311), .O(gate64inter8));
  nand2 gate226(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate227(.a(s_3), .b(gate64inter3), .O(gate64inter10));
  nor2  gate228(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate229(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate230(.a(gate64inter12), .b(gate64inter1), .O(N345));
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate357(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate358(.a(gate172inter0), .b(s_22), .O(gate172inter1));
  and2  gate359(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate360(.a(s_22), .O(gate172inter3));
  inv1  gate361(.a(s_23), .O(gate172inter4));
  nand2 gate362(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate363(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate364(.a(N5), .O(gate172inter7));
  inv1  gate365(.a(N693), .O(gate172inter8));
  nand2 gate366(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate367(.a(s_23), .b(gate172inter3), .O(gate172inter10));
  nor2  gate368(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate369(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate370(.a(gate172inter12), .b(gate172inter1), .O(N725));

  xor2  gate273(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate274(.a(gate173inter0), .b(s_10), .O(gate173inter1));
  and2  gate275(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate276(.a(s_10), .O(gate173inter3));
  inv1  gate277(.a(s_11), .O(gate173inter4));
  nand2 gate278(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate279(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate280(.a(N9), .O(gate173inter7));
  inv1  gate281(.a(N694), .O(gate173inter8));
  nand2 gate282(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate283(.a(s_11), .b(gate173inter3), .O(gate173inter10));
  nor2  gate284(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate285(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate286(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate343(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate344(.a(gate176inter0), .b(s_20), .O(gate176inter1));
  and2  gate345(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate346(.a(s_20), .O(gate176inter3));
  inv1  gate347(.a(s_21), .O(gate176inter4));
  nand2 gate348(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate349(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate350(.a(N21), .O(gate176inter7));
  inv1  gate351(.a(N697), .O(gate176inter8));
  nand2 gate352(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate353(.a(s_21), .b(gate176inter3), .O(gate176inter10));
  nor2  gate354(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate355(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate356(.a(gate176inter12), .b(gate176inter1), .O(N729));
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );

  xor2  gate245(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate246(.a(gate181inter0), .b(s_6), .O(gate181inter1));
  and2  gate247(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate248(.a(s_6), .O(gate181inter3));
  inv1  gate249(.a(s_7), .O(gate181inter4));
  nand2 gate250(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate251(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate252(.a(N41), .O(gate181inter7));
  inv1  gate253(.a(N702), .O(gate181inter8));
  nand2 gate254(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate255(.a(s_7), .b(gate181inter3), .O(gate181inter10));
  nor2  gate256(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate257(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate258(.a(gate181inter12), .b(gate181inter1), .O(N734));
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );

  xor2  gate315(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate316(.a(gate189inter0), .b(s_16), .O(gate189inter1));
  and2  gate317(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate318(.a(s_16), .O(gate189inter3));
  inv1  gate319(.a(s_17), .O(gate189inter4));
  nand2 gate320(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate321(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate322(.a(N73), .O(gate189inter7));
  inv1  gate323(.a(N710), .O(gate189inter8));
  nand2 gate324(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate325(.a(s_17), .b(gate189inter3), .O(gate189inter10));
  nor2  gate326(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate327(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate328(.a(gate189inter12), .b(gate189inter1), .O(N742));
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );

  xor2  gate301(.a(N714), .b(N89), .O(gate193inter0));
  nand2 gate302(.a(gate193inter0), .b(s_14), .O(gate193inter1));
  and2  gate303(.a(N714), .b(N89), .O(gate193inter2));
  inv1  gate304(.a(s_14), .O(gate193inter3));
  inv1  gate305(.a(s_15), .O(gate193inter4));
  nand2 gate306(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate307(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate308(.a(N89), .O(gate193inter7));
  inv1  gate309(.a(N714), .O(gate193inter8));
  nand2 gate310(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate311(.a(s_15), .b(gate193inter3), .O(gate193inter10));
  nor2  gate312(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate313(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate314(.a(gate193inter12), .b(gate193inter1), .O(N746));

  xor2  gate385(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate386(.a(gate194inter0), .b(s_26), .O(gate194inter1));
  and2  gate387(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate388(.a(s_26), .O(gate194inter3));
  inv1  gate389(.a(s_27), .O(gate194inter4));
  nand2 gate390(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate391(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate392(.a(N93), .O(gate194inter7));
  inv1  gate393(.a(N715), .O(gate194inter8));
  nand2 gate394(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate395(.a(s_27), .b(gate194inter3), .O(gate194inter10));
  nor2  gate396(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate397(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate398(.a(gate194inter12), .b(gate194inter1), .O(N747));

  xor2  gate371(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate372(.a(gate195inter0), .b(s_24), .O(gate195inter1));
  and2  gate373(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate374(.a(s_24), .O(gate195inter3));
  inv1  gate375(.a(s_25), .O(gate195inter4));
  nand2 gate376(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate377(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate378(.a(N97), .O(gate195inter7));
  inv1  gate379(.a(N716), .O(gate195inter8));
  nand2 gate380(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate381(.a(s_25), .b(gate195inter3), .O(gate195inter10));
  nor2  gate382(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate383(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate384(.a(gate195inter12), .b(gate195inter1), .O(N748));
xor2 gate196( .a(N101), .b(N717), .O(N749) );

  xor2  gate231(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate232(.a(gate197inter0), .b(s_4), .O(gate197inter1));
  and2  gate233(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate234(.a(s_4), .O(gate197inter3));
  inv1  gate235(.a(s_5), .O(gate197inter4));
  nand2 gate236(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate237(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate238(.a(N105), .O(gate197inter7));
  inv1  gate239(.a(N718), .O(gate197inter8));
  nand2 gate240(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate241(.a(s_5), .b(gate197inter3), .O(gate197inter10));
  nor2  gate242(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate243(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate244(.a(gate197inter12), .b(gate197inter1), .O(N750));

  xor2  gate399(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate400(.a(gate198inter0), .b(s_28), .O(gate198inter1));
  and2  gate401(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate402(.a(s_28), .O(gate198inter3));
  inv1  gate403(.a(s_29), .O(gate198inter4));
  nand2 gate404(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate405(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate406(.a(N109), .O(gate198inter7));
  inv1  gate407(.a(N719), .O(gate198inter8));
  nand2 gate408(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate409(.a(s_29), .b(gate198inter3), .O(gate198inter10));
  nor2  gate410(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate411(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate412(.a(gate198inter12), .b(gate198inter1), .O(N751));
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule