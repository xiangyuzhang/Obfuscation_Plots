module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1891(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1892(.a(gate12inter0), .b(s_192), .O(gate12inter1));
  and2  gate1893(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1894(.a(s_192), .O(gate12inter3));
  inv1  gate1895(.a(s_193), .O(gate12inter4));
  nand2 gate1896(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1897(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1898(.a(G7), .O(gate12inter7));
  inv1  gate1899(.a(G8), .O(gate12inter8));
  nand2 gate1900(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1901(.a(s_193), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1902(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1903(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1904(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1625(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1626(.a(gate16inter0), .b(s_154), .O(gate16inter1));
  and2  gate1627(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1628(.a(s_154), .O(gate16inter3));
  inv1  gate1629(.a(s_155), .O(gate16inter4));
  nand2 gate1630(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1631(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1632(.a(G15), .O(gate16inter7));
  inv1  gate1633(.a(G16), .O(gate16inter8));
  nand2 gate1634(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1635(.a(s_155), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1636(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1637(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1638(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1779(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1780(.a(gate18inter0), .b(s_176), .O(gate18inter1));
  and2  gate1781(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1782(.a(s_176), .O(gate18inter3));
  inv1  gate1783(.a(s_177), .O(gate18inter4));
  nand2 gate1784(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1785(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1786(.a(G19), .O(gate18inter7));
  inv1  gate1787(.a(G20), .O(gate18inter8));
  nand2 gate1788(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1789(.a(s_177), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1790(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1791(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1792(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1387(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1388(.a(gate20inter0), .b(s_120), .O(gate20inter1));
  and2  gate1389(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1390(.a(s_120), .O(gate20inter3));
  inv1  gate1391(.a(s_121), .O(gate20inter4));
  nand2 gate1392(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1393(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1394(.a(G23), .O(gate20inter7));
  inv1  gate1395(.a(G24), .O(gate20inter8));
  nand2 gate1396(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1397(.a(s_121), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1398(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1399(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1400(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate603(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate604(.a(gate22inter0), .b(s_8), .O(gate22inter1));
  and2  gate605(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate606(.a(s_8), .O(gate22inter3));
  inv1  gate607(.a(s_9), .O(gate22inter4));
  nand2 gate608(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate609(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate610(.a(G27), .O(gate22inter7));
  inv1  gate611(.a(G28), .O(gate22inter8));
  nand2 gate612(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate613(.a(s_9), .b(gate22inter3), .O(gate22inter10));
  nor2  gate614(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate615(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate616(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1835(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1836(.a(gate23inter0), .b(s_184), .O(gate23inter1));
  and2  gate1837(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1838(.a(s_184), .O(gate23inter3));
  inv1  gate1839(.a(s_185), .O(gate23inter4));
  nand2 gate1840(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1841(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1842(.a(G29), .O(gate23inter7));
  inv1  gate1843(.a(G30), .O(gate23inter8));
  nand2 gate1844(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1845(.a(s_185), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1846(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1847(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1848(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate687(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate688(.a(gate28inter0), .b(s_20), .O(gate28inter1));
  and2  gate689(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate690(.a(s_20), .O(gate28inter3));
  inv1  gate691(.a(s_21), .O(gate28inter4));
  nand2 gate692(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate693(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate694(.a(G10), .O(gate28inter7));
  inv1  gate695(.a(G14), .O(gate28inter8));
  nand2 gate696(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate697(.a(s_21), .b(gate28inter3), .O(gate28inter10));
  nor2  gate698(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate699(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate700(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1275(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1276(.a(gate29inter0), .b(s_104), .O(gate29inter1));
  and2  gate1277(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1278(.a(s_104), .O(gate29inter3));
  inv1  gate1279(.a(s_105), .O(gate29inter4));
  nand2 gate1280(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1281(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1282(.a(G3), .O(gate29inter7));
  inv1  gate1283(.a(G7), .O(gate29inter8));
  nand2 gate1284(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1285(.a(s_105), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1286(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1287(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1288(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate981(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate982(.a(gate32inter0), .b(s_62), .O(gate32inter1));
  and2  gate983(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate984(.a(s_62), .O(gate32inter3));
  inv1  gate985(.a(s_63), .O(gate32inter4));
  nand2 gate986(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate987(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate988(.a(G12), .O(gate32inter7));
  inv1  gate989(.a(G16), .O(gate32inter8));
  nand2 gate990(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate991(.a(s_63), .b(gate32inter3), .O(gate32inter10));
  nor2  gate992(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate993(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate994(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1121(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1122(.a(gate34inter0), .b(s_82), .O(gate34inter1));
  and2  gate1123(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1124(.a(s_82), .O(gate34inter3));
  inv1  gate1125(.a(s_83), .O(gate34inter4));
  nand2 gate1126(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1127(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1128(.a(G25), .O(gate34inter7));
  inv1  gate1129(.a(G29), .O(gate34inter8));
  nand2 gate1130(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1131(.a(s_83), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1132(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1133(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1134(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1247(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1248(.a(gate35inter0), .b(s_100), .O(gate35inter1));
  and2  gate1249(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1250(.a(s_100), .O(gate35inter3));
  inv1  gate1251(.a(s_101), .O(gate35inter4));
  nand2 gate1252(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1253(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1254(.a(G18), .O(gate35inter7));
  inv1  gate1255(.a(G22), .O(gate35inter8));
  nand2 gate1256(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1257(.a(s_101), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1258(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1259(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1260(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1415(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1416(.a(gate43inter0), .b(s_124), .O(gate43inter1));
  and2  gate1417(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1418(.a(s_124), .O(gate43inter3));
  inv1  gate1419(.a(s_125), .O(gate43inter4));
  nand2 gate1420(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1421(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1422(.a(G3), .O(gate43inter7));
  inv1  gate1423(.a(G269), .O(gate43inter8));
  nand2 gate1424(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1425(.a(s_125), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1426(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1427(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1428(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1709(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1710(.a(gate46inter0), .b(s_166), .O(gate46inter1));
  and2  gate1711(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1712(.a(s_166), .O(gate46inter3));
  inv1  gate1713(.a(s_167), .O(gate46inter4));
  nand2 gate1714(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1715(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1716(.a(G6), .O(gate46inter7));
  inv1  gate1717(.a(G272), .O(gate46inter8));
  nand2 gate1718(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1719(.a(s_167), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1720(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1721(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1722(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate855(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate856(.a(gate48inter0), .b(s_44), .O(gate48inter1));
  and2  gate857(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate858(.a(s_44), .O(gate48inter3));
  inv1  gate859(.a(s_45), .O(gate48inter4));
  nand2 gate860(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate861(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate862(.a(G8), .O(gate48inter7));
  inv1  gate863(.a(G275), .O(gate48inter8));
  nand2 gate864(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate865(.a(s_45), .b(gate48inter3), .O(gate48inter10));
  nor2  gate866(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate867(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate868(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1667(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1668(.a(gate49inter0), .b(s_160), .O(gate49inter1));
  and2  gate1669(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1670(.a(s_160), .O(gate49inter3));
  inv1  gate1671(.a(s_161), .O(gate49inter4));
  nand2 gate1672(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1673(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1674(.a(G9), .O(gate49inter7));
  inv1  gate1675(.a(G278), .O(gate49inter8));
  nand2 gate1676(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1677(.a(s_161), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1678(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1679(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1680(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1079(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1080(.a(gate55inter0), .b(s_76), .O(gate55inter1));
  and2  gate1081(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1082(.a(s_76), .O(gate55inter3));
  inv1  gate1083(.a(s_77), .O(gate55inter4));
  nand2 gate1084(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1085(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1086(.a(G15), .O(gate55inter7));
  inv1  gate1087(.a(G287), .O(gate55inter8));
  nand2 gate1088(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1089(.a(s_77), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1090(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1091(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1092(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate757(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate758(.a(gate58inter0), .b(s_30), .O(gate58inter1));
  and2  gate759(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate760(.a(s_30), .O(gate58inter3));
  inv1  gate761(.a(s_31), .O(gate58inter4));
  nand2 gate762(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate763(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate764(.a(G18), .O(gate58inter7));
  inv1  gate765(.a(G290), .O(gate58inter8));
  nand2 gate766(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate767(.a(s_31), .b(gate58inter3), .O(gate58inter10));
  nor2  gate768(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate769(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate770(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate1163(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1164(.a(gate59inter0), .b(s_88), .O(gate59inter1));
  and2  gate1165(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1166(.a(s_88), .O(gate59inter3));
  inv1  gate1167(.a(s_89), .O(gate59inter4));
  nand2 gate1168(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1169(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1170(.a(G19), .O(gate59inter7));
  inv1  gate1171(.a(G293), .O(gate59inter8));
  nand2 gate1172(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1173(.a(s_89), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1174(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1175(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1176(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate967(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate968(.a(gate62inter0), .b(s_60), .O(gate62inter1));
  and2  gate969(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate970(.a(s_60), .O(gate62inter3));
  inv1  gate971(.a(s_61), .O(gate62inter4));
  nand2 gate972(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate973(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate974(.a(G22), .O(gate62inter7));
  inv1  gate975(.a(G296), .O(gate62inter8));
  nand2 gate976(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate977(.a(s_61), .b(gate62inter3), .O(gate62inter10));
  nor2  gate978(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate979(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate980(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate561(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate562(.a(gate63inter0), .b(s_2), .O(gate63inter1));
  and2  gate563(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate564(.a(s_2), .O(gate63inter3));
  inv1  gate565(.a(s_3), .O(gate63inter4));
  nand2 gate566(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate567(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate568(.a(G23), .O(gate63inter7));
  inv1  gate569(.a(G299), .O(gate63inter8));
  nand2 gate570(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate571(.a(s_3), .b(gate63inter3), .O(gate63inter10));
  nor2  gate572(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate573(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate574(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1611(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1612(.a(gate64inter0), .b(s_152), .O(gate64inter1));
  and2  gate1613(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1614(.a(s_152), .O(gate64inter3));
  inv1  gate1615(.a(s_153), .O(gate64inter4));
  nand2 gate1616(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1617(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1618(.a(G24), .O(gate64inter7));
  inv1  gate1619(.a(G299), .O(gate64inter8));
  nand2 gate1620(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1621(.a(s_153), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1622(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1623(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1624(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate897(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate898(.a(gate71inter0), .b(s_50), .O(gate71inter1));
  and2  gate899(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate900(.a(s_50), .O(gate71inter3));
  inv1  gate901(.a(s_51), .O(gate71inter4));
  nand2 gate902(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate903(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate904(.a(G31), .O(gate71inter7));
  inv1  gate905(.a(G311), .O(gate71inter8));
  nand2 gate906(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate907(.a(s_51), .b(gate71inter3), .O(gate71inter10));
  nor2  gate908(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate909(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate910(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1401(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1402(.a(gate73inter0), .b(s_122), .O(gate73inter1));
  and2  gate1403(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1404(.a(s_122), .O(gate73inter3));
  inv1  gate1405(.a(s_123), .O(gate73inter4));
  nand2 gate1406(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1407(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1408(.a(G1), .O(gate73inter7));
  inv1  gate1409(.a(G314), .O(gate73inter8));
  nand2 gate1410(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1411(.a(s_123), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1412(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1413(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1414(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate911(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate912(.a(gate79inter0), .b(s_52), .O(gate79inter1));
  and2  gate913(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate914(.a(s_52), .O(gate79inter3));
  inv1  gate915(.a(s_53), .O(gate79inter4));
  nand2 gate916(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate917(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate918(.a(G10), .O(gate79inter7));
  inv1  gate919(.a(G323), .O(gate79inter8));
  nand2 gate920(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate921(.a(s_53), .b(gate79inter3), .O(gate79inter10));
  nor2  gate922(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate923(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate924(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1149(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1150(.a(gate89inter0), .b(s_86), .O(gate89inter1));
  and2  gate1151(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1152(.a(s_86), .O(gate89inter3));
  inv1  gate1153(.a(s_87), .O(gate89inter4));
  nand2 gate1154(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1155(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1156(.a(G17), .O(gate89inter7));
  inv1  gate1157(.a(G338), .O(gate89inter8));
  nand2 gate1158(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1159(.a(s_87), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1160(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1161(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1162(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate939(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate940(.a(gate98inter0), .b(s_56), .O(gate98inter1));
  and2  gate941(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate942(.a(s_56), .O(gate98inter3));
  inv1  gate943(.a(s_57), .O(gate98inter4));
  nand2 gate944(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate945(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate946(.a(G23), .O(gate98inter7));
  inv1  gate947(.a(G350), .O(gate98inter8));
  nand2 gate948(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate949(.a(s_57), .b(gate98inter3), .O(gate98inter10));
  nor2  gate950(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate951(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate952(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1443(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1444(.a(gate104inter0), .b(s_128), .O(gate104inter1));
  and2  gate1445(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1446(.a(s_128), .O(gate104inter3));
  inv1  gate1447(.a(s_129), .O(gate104inter4));
  nand2 gate1448(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1449(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1450(.a(G32), .O(gate104inter7));
  inv1  gate1451(.a(G359), .O(gate104inter8));
  nand2 gate1452(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1453(.a(s_129), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1454(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1455(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1456(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1905(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1906(.a(gate108inter0), .b(s_194), .O(gate108inter1));
  and2  gate1907(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1908(.a(s_194), .O(gate108inter3));
  inv1  gate1909(.a(s_195), .O(gate108inter4));
  nand2 gate1910(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1911(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1912(.a(G368), .O(gate108inter7));
  inv1  gate1913(.a(G369), .O(gate108inter8));
  nand2 gate1914(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1915(.a(s_195), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1916(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1917(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1918(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1331(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1332(.a(gate112inter0), .b(s_112), .O(gate112inter1));
  and2  gate1333(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1334(.a(s_112), .O(gate112inter3));
  inv1  gate1335(.a(s_113), .O(gate112inter4));
  nand2 gate1336(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1337(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1338(.a(G376), .O(gate112inter7));
  inv1  gate1339(.a(G377), .O(gate112inter8));
  nand2 gate1340(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1341(.a(s_113), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1342(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1343(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1344(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate659(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate660(.a(gate116inter0), .b(s_16), .O(gate116inter1));
  and2  gate661(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate662(.a(s_16), .O(gate116inter3));
  inv1  gate663(.a(s_17), .O(gate116inter4));
  nand2 gate664(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate665(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate666(.a(G384), .O(gate116inter7));
  inv1  gate667(.a(G385), .O(gate116inter8));
  nand2 gate668(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate669(.a(s_17), .b(gate116inter3), .O(gate116inter10));
  nor2  gate670(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate671(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate672(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate841(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate842(.a(gate122inter0), .b(s_42), .O(gate122inter1));
  and2  gate843(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate844(.a(s_42), .O(gate122inter3));
  inv1  gate845(.a(s_43), .O(gate122inter4));
  nand2 gate846(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate847(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate848(.a(G396), .O(gate122inter7));
  inv1  gate849(.a(G397), .O(gate122inter8));
  nand2 gate850(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate851(.a(s_43), .b(gate122inter3), .O(gate122inter10));
  nor2  gate852(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate853(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate854(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1009(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1010(.a(gate125inter0), .b(s_66), .O(gate125inter1));
  and2  gate1011(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1012(.a(s_66), .O(gate125inter3));
  inv1  gate1013(.a(s_67), .O(gate125inter4));
  nand2 gate1014(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1015(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1016(.a(G402), .O(gate125inter7));
  inv1  gate1017(.a(G403), .O(gate125inter8));
  nand2 gate1018(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1019(.a(s_67), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1020(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1021(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1022(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1107(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1108(.a(gate127inter0), .b(s_80), .O(gate127inter1));
  and2  gate1109(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1110(.a(s_80), .O(gate127inter3));
  inv1  gate1111(.a(s_81), .O(gate127inter4));
  nand2 gate1112(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1113(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1114(.a(G406), .O(gate127inter7));
  inv1  gate1115(.a(G407), .O(gate127inter8));
  nand2 gate1116(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1117(.a(s_81), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1118(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1119(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1120(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1499(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1500(.a(gate132inter0), .b(s_136), .O(gate132inter1));
  and2  gate1501(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1502(.a(s_136), .O(gate132inter3));
  inv1  gate1503(.a(s_137), .O(gate132inter4));
  nand2 gate1504(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1505(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1506(.a(G416), .O(gate132inter7));
  inv1  gate1507(.a(G417), .O(gate132inter8));
  nand2 gate1508(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1509(.a(s_137), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1510(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1511(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1512(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1807(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1808(.a(gate133inter0), .b(s_180), .O(gate133inter1));
  and2  gate1809(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1810(.a(s_180), .O(gate133inter3));
  inv1  gate1811(.a(s_181), .O(gate133inter4));
  nand2 gate1812(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1813(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1814(.a(G418), .O(gate133inter7));
  inv1  gate1815(.a(G419), .O(gate133inter8));
  nand2 gate1816(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1817(.a(s_181), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1818(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1819(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1820(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1751(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1752(.a(gate137inter0), .b(s_172), .O(gate137inter1));
  and2  gate1753(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1754(.a(s_172), .O(gate137inter3));
  inv1  gate1755(.a(s_173), .O(gate137inter4));
  nand2 gate1756(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1757(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1758(.a(G426), .O(gate137inter7));
  inv1  gate1759(.a(G429), .O(gate137inter8));
  nand2 gate1760(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1761(.a(s_173), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1762(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1763(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1764(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate785(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate786(.a(gate142inter0), .b(s_34), .O(gate142inter1));
  and2  gate787(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate788(.a(s_34), .O(gate142inter3));
  inv1  gate789(.a(s_35), .O(gate142inter4));
  nand2 gate790(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate791(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate792(.a(G456), .O(gate142inter7));
  inv1  gate793(.a(G459), .O(gate142inter8));
  nand2 gate794(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate795(.a(s_35), .b(gate142inter3), .O(gate142inter10));
  nor2  gate796(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate797(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate798(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1513(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1514(.a(gate147inter0), .b(s_138), .O(gate147inter1));
  and2  gate1515(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1516(.a(s_138), .O(gate147inter3));
  inv1  gate1517(.a(s_139), .O(gate147inter4));
  nand2 gate1518(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1519(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1520(.a(G486), .O(gate147inter7));
  inv1  gate1521(.a(G489), .O(gate147inter8));
  nand2 gate1522(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1523(.a(s_139), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1524(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1525(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1526(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1037(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1038(.a(gate148inter0), .b(s_70), .O(gate148inter1));
  and2  gate1039(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1040(.a(s_70), .O(gate148inter3));
  inv1  gate1041(.a(s_71), .O(gate148inter4));
  nand2 gate1042(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1043(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1044(.a(G492), .O(gate148inter7));
  inv1  gate1045(.a(G495), .O(gate148inter8));
  nand2 gate1046(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1047(.a(s_71), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1048(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1049(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1050(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1289(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1290(.a(gate150inter0), .b(s_106), .O(gate150inter1));
  and2  gate1291(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1292(.a(s_106), .O(gate150inter3));
  inv1  gate1293(.a(s_107), .O(gate150inter4));
  nand2 gate1294(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1295(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1296(.a(G504), .O(gate150inter7));
  inv1  gate1297(.a(G507), .O(gate150inter8));
  nand2 gate1298(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1299(.a(s_107), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1300(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1301(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1302(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate701(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate702(.a(gate151inter0), .b(s_22), .O(gate151inter1));
  and2  gate703(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate704(.a(s_22), .O(gate151inter3));
  inv1  gate705(.a(s_23), .O(gate151inter4));
  nand2 gate706(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate707(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate708(.a(G510), .O(gate151inter7));
  inv1  gate709(.a(G513), .O(gate151inter8));
  nand2 gate710(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate711(.a(s_23), .b(gate151inter3), .O(gate151inter10));
  nor2  gate712(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate713(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate714(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1527(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1528(.a(gate159inter0), .b(s_140), .O(gate159inter1));
  and2  gate1529(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1530(.a(s_140), .O(gate159inter3));
  inv1  gate1531(.a(s_141), .O(gate159inter4));
  nand2 gate1532(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1533(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1534(.a(G444), .O(gate159inter7));
  inv1  gate1535(.a(G531), .O(gate159inter8));
  nand2 gate1536(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1537(.a(s_141), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1538(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1539(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1540(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1471(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1472(.a(gate161inter0), .b(s_132), .O(gate161inter1));
  and2  gate1473(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1474(.a(s_132), .O(gate161inter3));
  inv1  gate1475(.a(s_133), .O(gate161inter4));
  nand2 gate1476(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1477(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1478(.a(G450), .O(gate161inter7));
  inv1  gate1479(.a(G534), .O(gate161inter8));
  nand2 gate1480(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1481(.a(s_133), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1482(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1483(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1484(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1639(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1640(.a(gate166inter0), .b(s_156), .O(gate166inter1));
  and2  gate1641(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1642(.a(s_156), .O(gate166inter3));
  inv1  gate1643(.a(s_157), .O(gate166inter4));
  nand2 gate1644(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1645(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1646(.a(G465), .O(gate166inter7));
  inv1  gate1647(.a(G540), .O(gate166inter8));
  nand2 gate1648(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1649(.a(s_157), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1650(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1651(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1652(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1177(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1178(.a(gate167inter0), .b(s_90), .O(gate167inter1));
  and2  gate1179(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1180(.a(s_90), .O(gate167inter3));
  inv1  gate1181(.a(s_91), .O(gate167inter4));
  nand2 gate1182(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1183(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1184(.a(G468), .O(gate167inter7));
  inv1  gate1185(.a(G543), .O(gate167inter8));
  nand2 gate1186(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1187(.a(s_91), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1188(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1189(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1190(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1023(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1024(.a(gate178inter0), .b(s_68), .O(gate178inter1));
  and2  gate1025(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1026(.a(s_68), .O(gate178inter3));
  inv1  gate1027(.a(s_69), .O(gate178inter4));
  nand2 gate1028(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1029(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1030(.a(G501), .O(gate178inter7));
  inv1  gate1031(.a(G558), .O(gate178inter8));
  nand2 gate1032(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1033(.a(s_69), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1034(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1035(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1036(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate589(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate590(.a(gate182inter0), .b(s_6), .O(gate182inter1));
  and2  gate591(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate592(.a(s_6), .O(gate182inter3));
  inv1  gate593(.a(s_7), .O(gate182inter4));
  nand2 gate594(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate595(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate596(.a(G513), .O(gate182inter7));
  inv1  gate597(.a(G564), .O(gate182inter8));
  nand2 gate598(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate599(.a(s_7), .b(gate182inter3), .O(gate182inter10));
  nor2  gate600(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate601(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate602(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1793(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1794(.a(gate185inter0), .b(s_178), .O(gate185inter1));
  and2  gate1795(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1796(.a(s_178), .O(gate185inter3));
  inv1  gate1797(.a(s_179), .O(gate185inter4));
  nand2 gate1798(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1799(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1800(.a(G570), .O(gate185inter7));
  inv1  gate1801(.a(G571), .O(gate185inter8));
  nand2 gate1802(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1803(.a(s_179), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1804(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1805(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1806(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1723(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1724(.a(gate191inter0), .b(s_168), .O(gate191inter1));
  and2  gate1725(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1726(.a(s_168), .O(gate191inter3));
  inv1  gate1727(.a(s_169), .O(gate191inter4));
  nand2 gate1728(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1729(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1730(.a(G582), .O(gate191inter7));
  inv1  gate1731(.a(G583), .O(gate191inter8));
  nand2 gate1732(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1733(.a(s_169), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1734(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1735(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1736(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate645(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate646(.a(gate195inter0), .b(s_14), .O(gate195inter1));
  and2  gate647(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate648(.a(s_14), .O(gate195inter3));
  inv1  gate649(.a(s_15), .O(gate195inter4));
  nand2 gate650(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate651(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate652(.a(G590), .O(gate195inter7));
  inv1  gate653(.a(G591), .O(gate195inter8));
  nand2 gate654(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate655(.a(s_15), .b(gate195inter3), .O(gate195inter10));
  nor2  gate656(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate657(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate658(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate673(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate674(.a(gate205inter0), .b(s_18), .O(gate205inter1));
  and2  gate675(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate676(.a(s_18), .O(gate205inter3));
  inv1  gate677(.a(s_19), .O(gate205inter4));
  nand2 gate678(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate679(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate680(.a(G622), .O(gate205inter7));
  inv1  gate681(.a(G627), .O(gate205inter8));
  nand2 gate682(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate683(.a(s_19), .b(gate205inter3), .O(gate205inter10));
  nor2  gate684(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate685(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate686(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1373(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1374(.a(gate207inter0), .b(s_118), .O(gate207inter1));
  and2  gate1375(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1376(.a(s_118), .O(gate207inter3));
  inv1  gate1377(.a(s_119), .O(gate207inter4));
  nand2 gate1378(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1379(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1380(.a(G622), .O(gate207inter7));
  inv1  gate1381(.a(G632), .O(gate207inter8));
  nand2 gate1382(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1383(.a(s_119), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1384(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1385(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1386(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1681(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1682(.a(gate208inter0), .b(s_162), .O(gate208inter1));
  and2  gate1683(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1684(.a(s_162), .O(gate208inter3));
  inv1  gate1685(.a(s_163), .O(gate208inter4));
  nand2 gate1686(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1687(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1688(.a(G627), .O(gate208inter7));
  inv1  gate1689(.a(G637), .O(gate208inter8));
  nand2 gate1690(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1691(.a(s_163), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1692(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1693(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1694(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1695(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1696(.a(gate209inter0), .b(s_164), .O(gate209inter1));
  and2  gate1697(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1698(.a(s_164), .O(gate209inter3));
  inv1  gate1699(.a(s_165), .O(gate209inter4));
  nand2 gate1700(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1701(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1702(.a(G602), .O(gate209inter7));
  inv1  gate1703(.a(G666), .O(gate209inter8));
  nand2 gate1704(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1705(.a(s_165), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1706(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1707(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1708(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1947(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1948(.a(gate210inter0), .b(s_200), .O(gate210inter1));
  and2  gate1949(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1950(.a(s_200), .O(gate210inter3));
  inv1  gate1951(.a(s_201), .O(gate210inter4));
  nand2 gate1952(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1953(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1954(.a(G607), .O(gate210inter7));
  inv1  gate1955(.a(G666), .O(gate210inter8));
  nand2 gate1956(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1957(.a(s_201), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1958(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1959(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1960(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate953(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate954(.a(gate216inter0), .b(s_58), .O(gate216inter1));
  and2  gate955(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate956(.a(s_58), .O(gate216inter3));
  inv1  gate957(.a(s_59), .O(gate216inter4));
  nand2 gate958(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate959(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate960(.a(G617), .O(gate216inter7));
  inv1  gate961(.a(G675), .O(gate216inter8));
  nand2 gate962(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate963(.a(s_59), .b(gate216inter3), .O(gate216inter10));
  nor2  gate964(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate965(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate966(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1821(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1822(.a(gate228inter0), .b(s_182), .O(gate228inter1));
  and2  gate1823(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1824(.a(s_182), .O(gate228inter3));
  inv1  gate1825(.a(s_183), .O(gate228inter4));
  nand2 gate1826(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1827(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1828(.a(G696), .O(gate228inter7));
  inv1  gate1829(.a(G697), .O(gate228inter8));
  nand2 gate1830(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1831(.a(s_183), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1832(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1833(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1834(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1359(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1360(.a(gate229inter0), .b(s_116), .O(gate229inter1));
  and2  gate1361(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1362(.a(s_116), .O(gate229inter3));
  inv1  gate1363(.a(s_117), .O(gate229inter4));
  nand2 gate1364(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1365(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1366(.a(G698), .O(gate229inter7));
  inv1  gate1367(.a(G699), .O(gate229inter8));
  nand2 gate1368(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1369(.a(s_117), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1370(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1371(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1372(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate883(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate884(.a(gate232inter0), .b(s_48), .O(gate232inter1));
  and2  gate885(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate886(.a(s_48), .O(gate232inter3));
  inv1  gate887(.a(s_49), .O(gate232inter4));
  nand2 gate888(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate889(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate890(.a(G704), .O(gate232inter7));
  inv1  gate891(.a(G705), .O(gate232inter8));
  nand2 gate892(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate893(.a(s_49), .b(gate232inter3), .O(gate232inter10));
  nor2  gate894(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate895(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate896(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate547(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate548(.a(gate233inter0), .b(s_0), .O(gate233inter1));
  and2  gate549(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate550(.a(s_0), .O(gate233inter3));
  inv1  gate551(.a(s_1), .O(gate233inter4));
  nand2 gate552(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate553(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate554(.a(G242), .O(gate233inter7));
  inv1  gate555(.a(G718), .O(gate233inter8));
  nand2 gate556(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate557(.a(s_1), .b(gate233inter3), .O(gate233inter10));
  nor2  gate558(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate559(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate560(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate925(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate926(.a(gate234inter0), .b(s_54), .O(gate234inter1));
  and2  gate927(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate928(.a(s_54), .O(gate234inter3));
  inv1  gate929(.a(s_55), .O(gate234inter4));
  nand2 gate930(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate931(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate932(.a(G245), .O(gate234inter7));
  inv1  gate933(.a(G721), .O(gate234inter8));
  nand2 gate934(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate935(.a(s_55), .b(gate234inter3), .O(gate234inter10));
  nor2  gate936(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate937(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate938(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1653(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1654(.a(gate235inter0), .b(s_158), .O(gate235inter1));
  and2  gate1655(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1656(.a(s_158), .O(gate235inter3));
  inv1  gate1657(.a(s_159), .O(gate235inter4));
  nand2 gate1658(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1659(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1660(.a(G248), .O(gate235inter7));
  inv1  gate1661(.a(G724), .O(gate235inter8));
  nand2 gate1662(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1663(.a(s_159), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1664(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1665(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1666(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1919(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1920(.a(gate237inter0), .b(s_196), .O(gate237inter1));
  and2  gate1921(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1922(.a(s_196), .O(gate237inter3));
  inv1  gate1923(.a(s_197), .O(gate237inter4));
  nand2 gate1924(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1925(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1926(.a(G254), .O(gate237inter7));
  inv1  gate1927(.a(G706), .O(gate237inter8));
  nand2 gate1928(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1929(.a(s_197), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1930(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1931(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1932(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1457(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1458(.a(gate238inter0), .b(s_130), .O(gate238inter1));
  and2  gate1459(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1460(.a(s_130), .O(gate238inter3));
  inv1  gate1461(.a(s_131), .O(gate238inter4));
  nand2 gate1462(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1463(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1464(.a(G257), .O(gate238inter7));
  inv1  gate1465(.a(G709), .O(gate238inter8));
  nand2 gate1466(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1467(.a(s_131), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1468(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1469(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1470(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate799(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate800(.a(gate244inter0), .b(s_36), .O(gate244inter1));
  and2  gate801(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate802(.a(s_36), .O(gate244inter3));
  inv1  gate803(.a(s_37), .O(gate244inter4));
  nand2 gate804(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate805(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate806(.a(G721), .O(gate244inter7));
  inv1  gate807(.a(G733), .O(gate244inter8));
  nand2 gate808(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate809(.a(s_37), .b(gate244inter3), .O(gate244inter10));
  nor2  gate810(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate811(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate812(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate995(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate996(.a(gate246inter0), .b(s_64), .O(gate246inter1));
  and2  gate997(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate998(.a(s_64), .O(gate246inter3));
  inv1  gate999(.a(s_65), .O(gate246inter4));
  nand2 gate1000(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1001(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1002(.a(G724), .O(gate246inter7));
  inv1  gate1003(.a(G736), .O(gate246inter8));
  nand2 gate1004(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1005(.a(s_65), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1006(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1007(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1008(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1555(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1556(.a(gate248inter0), .b(s_144), .O(gate248inter1));
  and2  gate1557(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1558(.a(s_144), .O(gate248inter3));
  inv1  gate1559(.a(s_145), .O(gate248inter4));
  nand2 gate1560(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1561(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1562(.a(G727), .O(gate248inter7));
  inv1  gate1563(.a(G739), .O(gate248inter8));
  nand2 gate1564(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1565(.a(s_145), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1566(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1567(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1568(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1219(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1220(.a(gate250inter0), .b(s_96), .O(gate250inter1));
  and2  gate1221(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1222(.a(s_96), .O(gate250inter3));
  inv1  gate1223(.a(s_97), .O(gate250inter4));
  nand2 gate1224(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1225(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1226(.a(G706), .O(gate250inter7));
  inv1  gate1227(.a(G742), .O(gate250inter8));
  nand2 gate1228(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1229(.a(s_97), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1230(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1231(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1232(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate813(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate814(.a(gate251inter0), .b(s_38), .O(gate251inter1));
  and2  gate815(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate816(.a(s_38), .O(gate251inter3));
  inv1  gate817(.a(s_39), .O(gate251inter4));
  nand2 gate818(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate819(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate820(.a(G257), .O(gate251inter7));
  inv1  gate821(.a(G745), .O(gate251inter8));
  nand2 gate822(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate823(.a(s_39), .b(gate251inter3), .O(gate251inter10));
  nor2  gate824(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate825(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate826(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1849(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1850(.a(gate254inter0), .b(s_186), .O(gate254inter1));
  and2  gate1851(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1852(.a(s_186), .O(gate254inter3));
  inv1  gate1853(.a(s_187), .O(gate254inter4));
  nand2 gate1854(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1855(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1856(.a(G712), .O(gate254inter7));
  inv1  gate1857(.a(G748), .O(gate254inter8));
  nand2 gate1858(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1859(.a(s_187), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1860(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1861(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1862(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1205(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1206(.a(gate261inter0), .b(s_94), .O(gate261inter1));
  and2  gate1207(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1208(.a(s_94), .O(gate261inter3));
  inv1  gate1209(.a(s_95), .O(gate261inter4));
  nand2 gate1210(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1211(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1212(.a(G762), .O(gate261inter7));
  inv1  gate1213(.a(G763), .O(gate261inter8));
  nand2 gate1214(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1215(.a(s_95), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1216(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1217(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1218(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1261(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1262(.a(gate267inter0), .b(s_102), .O(gate267inter1));
  and2  gate1263(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1264(.a(s_102), .O(gate267inter3));
  inv1  gate1265(.a(s_103), .O(gate267inter4));
  nand2 gate1266(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1267(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1268(.a(G648), .O(gate267inter7));
  inv1  gate1269(.a(G776), .O(gate267inter8));
  nand2 gate1270(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1271(.a(s_103), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1272(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1273(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1274(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1583(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1584(.a(gate269inter0), .b(s_148), .O(gate269inter1));
  and2  gate1585(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1586(.a(s_148), .O(gate269inter3));
  inv1  gate1587(.a(s_149), .O(gate269inter4));
  nand2 gate1588(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1589(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1590(.a(G654), .O(gate269inter7));
  inv1  gate1591(.a(G782), .O(gate269inter8));
  nand2 gate1592(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1593(.a(s_149), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1594(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1595(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1596(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate617(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate618(.a(gate273inter0), .b(s_10), .O(gate273inter1));
  and2  gate619(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate620(.a(s_10), .O(gate273inter3));
  inv1  gate621(.a(s_11), .O(gate273inter4));
  nand2 gate622(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate623(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate624(.a(G642), .O(gate273inter7));
  inv1  gate625(.a(G794), .O(gate273inter8));
  nand2 gate626(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate627(.a(s_11), .b(gate273inter3), .O(gate273inter10));
  nor2  gate628(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate629(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate630(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1863(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1864(.a(gate278inter0), .b(s_188), .O(gate278inter1));
  and2  gate1865(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1866(.a(s_188), .O(gate278inter3));
  inv1  gate1867(.a(s_189), .O(gate278inter4));
  nand2 gate1868(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1869(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1870(.a(G776), .O(gate278inter7));
  inv1  gate1871(.a(G800), .O(gate278inter8));
  nand2 gate1872(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1873(.a(s_189), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1874(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1875(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1876(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1569(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1570(.a(gate280inter0), .b(s_146), .O(gate280inter1));
  and2  gate1571(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1572(.a(s_146), .O(gate280inter3));
  inv1  gate1573(.a(s_147), .O(gate280inter4));
  nand2 gate1574(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1575(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1576(.a(G779), .O(gate280inter7));
  inv1  gate1577(.a(G803), .O(gate280inter8));
  nand2 gate1578(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1579(.a(s_147), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1580(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1581(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1582(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1093(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1094(.a(gate284inter0), .b(s_78), .O(gate284inter1));
  and2  gate1095(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1096(.a(s_78), .O(gate284inter3));
  inv1  gate1097(.a(s_79), .O(gate284inter4));
  nand2 gate1098(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1099(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1100(.a(G785), .O(gate284inter7));
  inv1  gate1101(.a(G809), .O(gate284inter8));
  nand2 gate1102(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1103(.a(s_79), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1104(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1105(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1106(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate827(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate828(.a(gate285inter0), .b(s_40), .O(gate285inter1));
  and2  gate829(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate830(.a(s_40), .O(gate285inter3));
  inv1  gate831(.a(s_41), .O(gate285inter4));
  nand2 gate832(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate833(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate834(.a(G660), .O(gate285inter7));
  inv1  gate835(.a(G812), .O(gate285inter8));
  nand2 gate836(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate837(.a(s_41), .b(gate285inter3), .O(gate285inter10));
  nor2  gate838(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate839(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate840(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1485(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1486(.a(gate288inter0), .b(s_134), .O(gate288inter1));
  and2  gate1487(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1488(.a(s_134), .O(gate288inter3));
  inv1  gate1489(.a(s_135), .O(gate288inter4));
  nand2 gate1490(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1491(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1492(.a(G791), .O(gate288inter7));
  inv1  gate1493(.a(G815), .O(gate288inter8));
  nand2 gate1494(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1495(.a(s_135), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1496(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1497(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1498(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate715(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate716(.a(gate290inter0), .b(s_24), .O(gate290inter1));
  and2  gate717(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate718(.a(s_24), .O(gate290inter3));
  inv1  gate719(.a(s_25), .O(gate290inter4));
  nand2 gate720(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate721(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate722(.a(G820), .O(gate290inter7));
  inv1  gate723(.a(G821), .O(gate290inter8));
  nand2 gate724(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate725(.a(s_25), .b(gate290inter3), .O(gate290inter10));
  nor2  gate726(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate727(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate728(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate631(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate632(.a(gate391inter0), .b(s_12), .O(gate391inter1));
  and2  gate633(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate634(.a(s_12), .O(gate391inter3));
  inv1  gate635(.a(s_13), .O(gate391inter4));
  nand2 gate636(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate637(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate638(.a(G5), .O(gate391inter7));
  inv1  gate639(.a(G1048), .O(gate391inter8));
  nand2 gate640(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate641(.a(s_13), .b(gate391inter3), .O(gate391inter10));
  nor2  gate642(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate643(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate644(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1065(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1066(.a(gate393inter0), .b(s_74), .O(gate393inter1));
  and2  gate1067(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1068(.a(s_74), .O(gate393inter3));
  inv1  gate1069(.a(s_75), .O(gate393inter4));
  nand2 gate1070(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1071(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1072(.a(G7), .O(gate393inter7));
  inv1  gate1073(.a(G1054), .O(gate393inter8));
  nand2 gate1074(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1075(.a(s_75), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1076(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1077(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1078(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1541(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1542(.a(gate407inter0), .b(s_142), .O(gate407inter1));
  and2  gate1543(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1544(.a(s_142), .O(gate407inter3));
  inv1  gate1545(.a(s_143), .O(gate407inter4));
  nand2 gate1546(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1547(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1548(.a(G21), .O(gate407inter7));
  inv1  gate1549(.a(G1096), .O(gate407inter8));
  nand2 gate1550(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1551(.a(s_143), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1552(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1553(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1554(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate575(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate576(.a(gate420inter0), .b(s_4), .O(gate420inter1));
  and2  gate577(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate578(.a(s_4), .O(gate420inter3));
  inv1  gate579(.a(s_5), .O(gate420inter4));
  nand2 gate580(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate581(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate582(.a(G1036), .O(gate420inter7));
  inv1  gate583(.a(G1132), .O(gate420inter8));
  nand2 gate584(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate585(.a(s_5), .b(gate420inter3), .O(gate420inter10));
  nor2  gate586(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate587(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate588(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1737(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1738(.a(gate426inter0), .b(s_170), .O(gate426inter1));
  and2  gate1739(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1740(.a(s_170), .O(gate426inter3));
  inv1  gate1741(.a(s_171), .O(gate426inter4));
  nand2 gate1742(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1743(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1744(.a(G1045), .O(gate426inter7));
  inv1  gate1745(.a(G1141), .O(gate426inter8));
  nand2 gate1746(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1747(.a(s_171), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1748(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1749(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1750(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1191(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1192(.a(gate432inter0), .b(s_92), .O(gate432inter1));
  and2  gate1193(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1194(.a(s_92), .O(gate432inter3));
  inv1  gate1195(.a(s_93), .O(gate432inter4));
  nand2 gate1196(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1197(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1198(.a(G1054), .O(gate432inter7));
  inv1  gate1199(.a(G1150), .O(gate432inter8));
  nand2 gate1200(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1201(.a(s_93), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1202(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1203(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1204(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1135(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1136(.a(gate434inter0), .b(s_84), .O(gate434inter1));
  and2  gate1137(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1138(.a(s_84), .O(gate434inter3));
  inv1  gate1139(.a(s_85), .O(gate434inter4));
  nand2 gate1140(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1141(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1142(.a(G1057), .O(gate434inter7));
  inv1  gate1143(.a(G1153), .O(gate434inter8));
  nand2 gate1144(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1145(.a(s_85), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1146(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1147(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1148(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1317(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1318(.a(gate439inter0), .b(s_110), .O(gate439inter1));
  and2  gate1319(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1320(.a(s_110), .O(gate439inter3));
  inv1  gate1321(.a(s_111), .O(gate439inter4));
  nand2 gate1322(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1323(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1324(.a(G11), .O(gate439inter7));
  inv1  gate1325(.a(G1162), .O(gate439inter8));
  nand2 gate1326(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1327(.a(s_111), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1328(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1329(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1330(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1765(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1766(.a(gate449inter0), .b(s_174), .O(gate449inter1));
  and2  gate1767(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1768(.a(s_174), .O(gate449inter3));
  inv1  gate1769(.a(s_175), .O(gate449inter4));
  nand2 gate1770(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1771(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1772(.a(G16), .O(gate449inter7));
  inv1  gate1773(.a(G1177), .O(gate449inter8));
  nand2 gate1774(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1775(.a(s_175), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1776(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1777(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1778(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate771(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate772(.a(gate450inter0), .b(s_32), .O(gate450inter1));
  and2  gate773(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate774(.a(s_32), .O(gate450inter3));
  inv1  gate775(.a(s_33), .O(gate450inter4));
  nand2 gate776(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate777(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate778(.a(G1081), .O(gate450inter7));
  inv1  gate779(.a(G1177), .O(gate450inter8));
  nand2 gate780(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate781(.a(s_33), .b(gate450inter3), .O(gate450inter10));
  nor2  gate782(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate783(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate784(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1933(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1934(.a(gate453inter0), .b(s_198), .O(gate453inter1));
  and2  gate1935(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1936(.a(s_198), .O(gate453inter3));
  inv1  gate1937(.a(s_199), .O(gate453inter4));
  nand2 gate1938(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1939(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1940(.a(G18), .O(gate453inter7));
  inv1  gate1941(.a(G1183), .O(gate453inter8));
  nand2 gate1942(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1943(.a(s_199), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1944(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1945(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1946(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1303(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1304(.a(gate459inter0), .b(s_108), .O(gate459inter1));
  and2  gate1305(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1306(.a(s_108), .O(gate459inter3));
  inv1  gate1307(.a(s_109), .O(gate459inter4));
  nand2 gate1308(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1309(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1310(.a(G21), .O(gate459inter7));
  inv1  gate1311(.a(G1192), .O(gate459inter8));
  nand2 gate1312(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1313(.a(s_109), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1314(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1315(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1316(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1345(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1346(.a(gate461inter0), .b(s_114), .O(gate461inter1));
  and2  gate1347(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1348(.a(s_114), .O(gate461inter3));
  inv1  gate1349(.a(s_115), .O(gate461inter4));
  nand2 gate1350(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1351(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1352(.a(G22), .O(gate461inter7));
  inv1  gate1353(.a(G1195), .O(gate461inter8));
  nand2 gate1354(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1355(.a(s_115), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1356(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1357(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1358(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate729(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate730(.a(gate473inter0), .b(s_26), .O(gate473inter1));
  and2  gate731(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate732(.a(s_26), .O(gate473inter3));
  inv1  gate733(.a(s_27), .O(gate473inter4));
  nand2 gate734(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate735(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate736(.a(G28), .O(gate473inter7));
  inv1  gate737(.a(G1213), .O(gate473inter8));
  nand2 gate738(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate739(.a(s_27), .b(gate473inter3), .O(gate473inter10));
  nor2  gate740(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate741(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate742(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1877(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1878(.a(gate478inter0), .b(s_190), .O(gate478inter1));
  and2  gate1879(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1880(.a(s_190), .O(gate478inter3));
  inv1  gate1881(.a(s_191), .O(gate478inter4));
  nand2 gate1882(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1883(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1884(.a(G1123), .O(gate478inter7));
  inv1  gate1885(.a(G1219), .O(gate478inter8));
  nand2 gate1886(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1887(.a(s_191), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1888(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1889(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1890(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1429(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1430(.a(gate485inter0), .b(s_126), .O(gate485inter1));
  and2  gate1431(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1432(.a(s_126), .O(gate485inter3));
  inv1  gate1433(.a(s_127), .O(gate485inter4));
  nand2 gate1434(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1435(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1436(.a(G1232), .O(gate485inter7));
  inv1  gate1437(.a(G1233), .O(gate485inter8));
  nand2 gate1438(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1439(.a(s_127), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1440(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1441(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1442(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1233(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1234(.a(gate488inter0), .b(s_98), .O(gate488inter1));
  and2  gate1235(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1236(.a(s_98), .O(gate488inter3));
  inv1  gate1237(.a(s_99), .O(gate488inter4));
  nand2 gate1238(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1239(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1240(.a(G1238), .O(gate488inter7));
  inv1  gate1241(.a(G1239), .O(gate488inter8));
  nand2 gate1242(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1243(.a(s_99), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1244(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1245(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1246(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1597(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1598(.a(gate490inter0), .b(s_150), .O(gate490inter1));
  and2  gate1599(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1600(.a(s_150), .O(gate490inter3));
  inv1  gate1601(.a(s_151), .O(gate490inter4));
  nand2 gate1602(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1603(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1604(.a(G1242), .O(gate490inter7));
  inv1  gate1605(.a(G1243), .O(gate490inter8));
  nand2 gate1606(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1607(.a(s_151), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1608(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1609(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1610(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate869(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate870(.a(gate500inter0), .b(s_46), .O(gate500inter1));
  and2  gate871(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate872(.a(s_46), .O(gate500inter3));
  inv1  gate873(.a(s_47), .O(gate500inter4));
  nand2 gate874(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate875(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate876(.a(G1262), .O(gate500inter7));
  inv1  gate877(.a(G1263), .O(gate500inter8));
  nand2 gate878(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate879(.a(s_47), .b(gate500inter3), .O(gate500inter10));
  nor2  gate880(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate881(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate882(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate743(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate744(.a(gate502inter0), .b(s_28), .O(gate502inter1));
  and2  gate745(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate746(.a(s_28), .O(gate502inter3));
  inv1  gate747(.a(s_29), .O(gate502inter4));
  nand2 gate748(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate749(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate750(.a(G1266), .O(gate502inter7));
  inv1  gate751(.a(G1267), .O(gate502inter8));
  nand2 gate752(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate753(.a(s_29), .b(gate502inter3), .O(gate502inter10));
  nor2  gate754(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate755(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate756(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1051(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1052(.a(gate508inter0), .b(s_72), .O(gate508inter1));
  and2  gate1053(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1054(.a(s_72), .O(gate508inter3));
  inv1  gate1055(.a(s_73), .O(gate508inter4));
  nand2 gate1056(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1057(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1058(.a(G1278), .O(gate508inter7));
  inv1  gate1059(.a(G1279), .O(gate508inter8));
  nand2 gate1060(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1061(.a(s_73), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1062(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1063(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1064(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule