module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1527(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1528(.a(gate12inter0), .b(s_140), .O(gate12inter1));
  and2  gate1529(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1530(.a(s_140), .O(gate12inter3));
  inv1  gate1531(.a(s_141), .O(gate12inter4));
  nand2 gate1532(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1533(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1534(.a(G7), .O(gate12inter7));
  inv1  gate1535(.a(G8), .O(gate12inter8));
  nand2 gate1536(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1537(.a(s_141), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1538(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1539(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1540(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1961(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1962(.a(gate21inter0), .b(s_202), .O(gate21inter1));
  and2  gate1963(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1964(.a(s_202), .O(gate21inter3));
  inv1  gate1965(.a(s_203), .O(gate21inter4));
  nand2 gate1966(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1967(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1968(.a(G25), .O(gate21inter7));
  inv1  gate1969(.a(G26), .O(gate21inter8));
  nand2 gate1970(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1971(.a(s_203), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1972(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1973(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1974(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1723(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1724(.a(gate22inter0), .b(s_168), .O(gate22inter1));
  and2  gate1725(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1726(.a(s_168), .O(gate22inter3));
  inv1  gate1727(.a(s_169), .O(gate22inter4));
  nand2 gate1728(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1729(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1730(.a(G27), .O(gate22inter7));
  inv1  gate1731(.a(G28), .O(gate22inter8));
  nand2 gate1732(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1733(.a(s_169), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1734(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1735(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1736(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1569(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1570(.a(gate24inter0), .b(s_146), .O(gate24inter1));
  and2  gate1571(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1572(.a(s_146), .O(gate24inter3));
  inv1  gate1573(.a(s_147), .O(gate24inter4));
  nand2 gate1574(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1575(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1576(.a(G31), .O(gate24inter7));
  inv1  gate1577(.a(G32), .O(gate24inter8));
  nand2 gate1578(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1579(.a(s_147), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1580(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1581(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1582(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate561(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate562(.a(gate27inter0), .b(s_2), .O(gate27inter1));
  and2  gate563(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate564(.a(s_2), .O(gate27inter3));
  inv1  gate565(.a(s_3), .O(gate27inter4));
  nand2 gate566(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate567(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate568(.a(G2), .O(gate27inter7));
  inv1  gate569(.a(G6), .O(gate27inter8));
  nand2 gate570(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate571(.a(s_3), .b(gate27inter3), .O(gate27inter10));
  nor2  gate572(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate573(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate574(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1303(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1304(.a(gate28inter0), .b(s_108), .O(gate28inter1));
  and2  gate1305(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1306(.a(s_108), .O(gate28inter3));
  inv1  gate1307(.a(s_109), .O(gate28inter4));
  nand2 gate1308(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1309(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1310(.a(G10), .O(gate28inter7));
  inv1  gate1311(.a(G14), .O(gate28inter8));
  nand2 gate1312(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1313(.a(s_109), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1314(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1315(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1316(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1611(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1612(.a(gate34inter0), .b(s_152), .O(gate34inter1));
  and2  gate1613(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1614(.a(s_152), .O(gate34inter3));
  inv1  gate1615(.a(s_153), .O(gate34inter4));
  nand2 gate1616(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1617(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1618(.a(G25), .O(gate34inter7));
  inv1  gate1619(.a(G29), .O(gate34inter8));
  nand2 gate1620(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1621(.a(s_153), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1622(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1623(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1624(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1429(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1430(.a(gate36inter0), .b(s_126), .O(gate36inter1));
  and2  gate1431(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1432(.a(s_126), .O(gate36inter3));
  inv1  gate1433(.a(s_127), .O(gate36inter4));
  nand2 gate1434(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1435(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1436(.a(G26), .O(gate36inter7));
  inv1  gate1437(.a(G30), .O(gate36inter8));
  nand2 gate1438(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1439(.a(s_127), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1440(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1441(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1442(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1709(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1710(.a(gate42inter0), .b(s_166), .O(gate42inter1));
  and2  gate1711(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1712(.a(s_166), .O(gate42inter3));
  inv1  gate1713(.a(s_167), .O(gate42inter4));
  nand2 gate1714(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1715(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1716(.a(G2), .O(gate42inter7));
  inv1  gate1717(.a(G266), .O(gate42inter8));
  nand2 gate1718(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1719(.a(s_167), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1720(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1721(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1722(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1681(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1682(.a(gate44inter0), .b(s_162), .O(gate44inter1));
  and2  gate1683(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1684(.a(s_162), .O(gate44inter3));
  inv1  gate1685(.a(s_163), .O(gate44inter4));
  nand2 gate1686(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1687(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1688(.a(G4), .O(gate44inter7));
  inv1  gate1689(.a(G269), .O(gate44inter8));
  nand2 gate1690(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1691(.a(s_163), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1692(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1693(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1694(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2143(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2144(.a(gate45inter0), .b(s_228), .O(gate45inter1));
  and2  gate2145(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2146(.a(s_228), .O(gate45inter3));
  inv1  gate2147(.a(s_229), .O(gate45inter4));
  nand2 gate2148(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2149(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2150(.a(G5), .O(gate45inter7));
  inv1  gate2151(.a(G272), .O(gate45inter8));
  nand2 gate2152(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2153(.a(s_229), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2154(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2155(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2156(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2437(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2438(.a(gate49inter0), .b(s_270), .O(gate49inter1));
  and2  gate2439(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2440(.a(s_270), .O(gate49inter3));
  inv1  gate2441(.a(s_271), .O(gate49inter4));
  nand2 gate2442(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2443(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2444(.a(G9), .O(gate49inter7));
  inv1  gate2445(.a(G278), .O(gate49inter8));
  nand2 gate2446(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2447(.a(s_271), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2448(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2449(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2450(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1163(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1164(.a(gate51inter0), .b(s_88), .O(gate51inter1));
  and2  gate1165(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1166(.a(s_88), .O(gate51inter3));
  inv1  gate1167(.a(s_89), .O(gate51inter4));
  nand2 gate1168(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1169(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1170(.a(G11), .O(gate51inter7));
  inv1  gate1171(.a(G281), .O(gate51inter8));
  nand2 gate1172(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1173(.a(s_89), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1174(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1175(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1176(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1751(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1752(.a(gate52inter0), .b(s_172), .O(gate52inter1));
  and2  gate1753(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1754(.a(s_172), .O(gate52inter3));
  inv1  gate1755(.a(s_173), .O(gate52inter4));
  nand2 gate1756(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1757(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1758(.a(G12), .O(gate52inter7));
  inv1  gate1759(.a(G281), .O(gate52inter8));
  nand2 gate1760(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1761(.a(s_173), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1762(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1763(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1764(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1219(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1220(.a(gate56inter0), .b(s_96), .O(gate56inter1));
  and2  gate1221(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1222(.a(s_96), .O(gate56inter3));
  inv1  gate1223(.a(s_97), .O(gate56inter4));
  nand2 gate1224(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1225(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1226(.a(G16), .O(gate56inter7));
  inv1  gate1227(.a(G287), .O(gate56inter8));
  nand2 gate1228(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1229(.a(s_97), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1230(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1231(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1232(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2241(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2242(.a(gate58inter0), .b(s_242), .O(gate58inter1));
  and2  gate2243(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2244(.a(s_242), .O(gate58inter3));
  inv1  gate2245(.a(s_243), .O(gate58inter4));
  nand2 gate2246(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2247(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2248(.a(G18), .O(gate58inter7));
  inv1  gate2249(.a(G290), .O(gate58inter8));
  nand2 gate2250(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2251(.a(s_243), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2252(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2253(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2254(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate575(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate576(.a(gate59inter0), .b(s_4), .O(gate59inter1));
  and2  gate577(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate578(.a(s_4), .O(gate59inter3));
  inv1  gate579(.a(s_5), .O(gate59inter4));
  nand2 gate580(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate581(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate582(.a(G19), .O(gate59inter7));
  inv1  gate583(.a(G293), .O(gate59inter8));
  nand2 gate584(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate585(.a(s_5), .b(gate59inter3), .O(gate59inter10));
  nor2  gate586(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate587(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate588(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2017(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2018(.a(gate61inter0), .b(s_210), .O(gate61inter1));
  and2  gate2019(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2020(.a(s_210), .O(gate61inter3));
  inv1  gate2021(.a(s_211), .O(gate61inter4));
  nand2 gate2022(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2023(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2024(.a(G21), .O(gate61inter7));
  inv1  gate2025(.a(G296), .O(gate61inter8));
  nand2 gate2026(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2027(.a(s_211), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2028(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2029(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2030(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate2423(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2424(.a(gate62inter0), .b(s_268), .O(gate62inter1));
  and2  gate2425(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2426(.a(s_268), .O(gate62inter3));
  inv1  gate2427(.a(s_269), .O(gate62inter4));
  nand2 gate2428(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2429(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2430(.a(G22), .O(gate62inter7));
  inv1  gate2431(.a(G296), .O(gate62inter8));
  nand2 gate2432(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2433(.a(s_269), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2434(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2435(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2436(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1247(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1248(.a(gate63inter0), .b(s_100), .O(gate63inter1));
  and2  gate1249(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1250(.a(s_100), .O(gate63inter3));
  inv1  gate1251(.a(s_101), .O(gate63inter4));
  nand2 gate1252(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1253(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1254(.a(G23), .O(gate63inter7));
  inv1  gate1255(.a(G299), .O(gate63inter8));
  nand2 gate1256(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1257(.a(s_101), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1258(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1259(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1260(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1457(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1458(.a(gate65inter0), .b(s_130), .O(gate65inter1));
  and2  gate1459(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1460(.a(s_130), .O(gate65inter3));
  inv1  gate1461(.a(s_131), .O(gate65inter4));
  nand2 gate1462(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1463(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1464(.a(G25), .O(gate65inter7));
  inv1  gate1465(.a(G302), .O(gate65inter8));
  nand2 gate1466(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1467(.a(s_131), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1468(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1469(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1470(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1289(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1290(.a(gate67inter0), .b(s_106), .O(gate67inter1));
  and2  gate1291(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1292(.a(s_106), .O(gate67inter3));
  inv1  gate1293(.a(s_107), .O(gate67inter4));
  nand2 gate1294(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1295(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1296(.a(G27), .O(gate67inter7));
  inv1  gate1297(.a(G305), .O(gate67inter8));
  nand2 gate1298(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1299(.a(s_107), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1300(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1301(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1302(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2213(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2214(.a(gate70inter0), .b(s_238), .O(gate70inter1));
  and2  gate2215(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2216(.a(s_238), .O(gate70inter3));
  inv1  gate2217(.a(s_239), .O(gate70inter4));
  nand2 gate2218(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2219(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2220(.a(G30), .O(gate70inter7));
  inv1  gate2221(.a(G308), .O(gate70inter8));
  nand2 gate2222(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2223(.a(s_239), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2224(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2225(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2226(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1975(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1976(.a(gate72inter0), .b(s_204), .O(gate72inter1));
  and2  gate1977(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1978(.a(s_204), .O(gate72inter3));
  inv1  gate1979(.a(s_205), .O(gate72inter4));
  nand2 gate1980(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1981(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1982(.a(G32), .O(gate72inter7));
  inv1  gate1983(.a(G311), .O(gate72inter8));
  nand2 gate1984(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1985(.a(s_205), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1986(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1987(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1988(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2101(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2102(.a(gate74inter0), .b(s_222), .O(gate74inter1));
  and2  gate2103(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2104(.a(s_222), .O(gate74inter3));
  inv1  gate2105(.a(s_223), .O(gate74inter4));
  nand2 gate2106(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2107(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2108(.a(G5), .O(gate74inter7));
  inv1  gate2109(.a(G314), .O(gate74inter8));
  nand2 gate2110(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2111(.a(s_223), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2112(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2113(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2114(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate813(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate814(.a(gate78inter0), .b(s_38), .O(gate78inter1));
  and2  gate815(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate816(.a(s_38), .O(gate78inter3));
  inv1  gate817(.a(s_39), .O(gate78inter4));
  nand2 gate818(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate819(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate820(.a(G6), .O(gate78inter7));
  inv1  gate821(.a(G320), .O(gate78inter8));
  nand2 gate822(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate823(.a(s_39), .b(gate78inter3), .O(gate78inter10));
  nor2  gate824(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate825(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate826(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2381(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2382(.a(gate79inter0), .b(s_262), .O(gate79inter1));
  and2  gate2383(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2384(.a(s_262), .O(gate79inter3));
  inv1  gate2385(.a(s_263), .O(gate79inter4));
  nand2 gate2386(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2387(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2388(.a(G10), .O(gate79inter7));
  inv1  gate2389(.a(G323), .O(gate79inter8));
  nand2 gate2390(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2391(.a(s_263), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2392(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2393(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2394(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2297(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2298(.a(gate82inter0), .b(s_250), .O(gate82inter1));
  and2  gate2299(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2300(.a(s_250), .O(gate82inter3));
  inv1  gate2301(.a(s_251), .O(gate82inter4));
  nand2 gate2302(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2303(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2304(.a(G7), .O(gate82inter7));
  inv1  gate2305(.a(G326), .O(gate82inter8));
  nand2 gate2306(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2307(.a(s_251), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2308(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2309(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2310(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2255(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2256(.a(gate86inter0), .b(s_244), .O(gate86inter1));
  and2  gate2257(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2258(.a(s_244), .O(gate86inter3));
  inv1  gate2259(.a(s_245), .O(gate86inter4));
  nand2 gate2260(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2261(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2262(.a(G8), .O(gate86inter7));
  inv1  gate2263(.a(G332), .O(gate86inter8));
  nand2 gate2264(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2265(.a(s_245), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2266(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2267(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2268(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2325(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2326(.a(gate91inter0), .b(s_254), .O(gate91inter1));
  and2  gate2327(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2328(.a(s_254), .O(gate91inter3));
  inv1  gate2329(.a(s_255), .O(gate91inter4));
  nand2 gate2330(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2331(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2332(.a(G25), .O(gate91inter7));
  inv1  gate2333(.a(G341), .O(gate91inter8));
  nand2 gate2334(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2335(.a(s_255), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2336(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2337(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2338(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2115(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2116(.a(gate95inter0), .b(s_224), .O(gate95inter1));
  and2  gate2117(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2118(.a(s_224), .O(gate95inter3));
  inv1  gate2119(.a(s_225), .O(gate95inter4));
  nand2 gate2120(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2121(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2122(.a(G26), .O(gate95inter7));
  inv1  gate2123(.a(G347), .O(gate95inter8));
  nand2 gate2124(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2125(.a(s_225), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2126(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2127(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2128(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1597(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1598(.a(gate99inter0), .b(s_150), .O(gate99inter1));
  and2  gate1599(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1600(.a(s_150), .O(gate99inter3));
  inv1  gate1601(.a(s_151), .O(gate99inter4));
  nand2 gate1602(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1603(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1604(.a(G27), .O(gate99inter7));
  inv1  gate1605(.a(G353), .O(gate99inter8));
  nand2 gate1606(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1607(.a(s_151), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1608(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1609(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1610(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate617(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate618(.a(gate107inter0), .b(s_10), .O(gate107inter1));
  and2  gate619(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate620(.a(s_10), .O(gate107inter3));
  inv1  gate621(.a(s_11), .O(gate107inter4));
  nand2 gate622(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate623(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate624(.a(G366), .O(gate107inter7));
  inv1  gate625(.a(G367), .O(gate107inter8));
  nand2 gate626(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate627(.a(s_11), .b(gate107inter3), .O(gate107inter10));
  nor2  gate628(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate629(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate630(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate2045(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate2046(.a(gate110inter0), .b(s_214), .O(gate110inter1));
  and2  gate2047(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate2048(.a(s_214), .O(gate110inter3));
  inv1  gate2049(.a(s_215), .O(gate110inter4));
  nand2 gate2050(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate2051(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate2052(.a(G372), .O(gate110inter7));
  inv1  gate2053(.a(G373), .O(gate110inter8));
  nand2 gate2054(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate2055(.a(s_215), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2056(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2057(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2058(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate939(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate940(.a(gate113inter0), .b(s_56), .O(gate113inter1));
  and2  gate941(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate942(.a(s_56), .O(gate113inter3));
  inv1  gate943(.a(s_57), .O(gate113inter4));
  nand2 gate944(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate945(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate946(.a(G378), .O(gate113inter7));
  inv1  gate947(.a(G379), .O(gate113inter8));
  nand2 gate948(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate949(.a(s_57), .b(gate113inter3), .O(gate113inter10));
  nor2  gate950(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate951(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate952(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate1695(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1696(.a(gate114inter0), .b(s_164), .O(gate114inter1));
  and2  gate1697(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1698(.a(s_164), .O(gate114inter3));
  inv1  gate1699(.a(s_165), .O(gate114inter4));
  nand2 gate1700(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1701(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1702(.a(G380), .O(gate114inter7));
  inv1  gate1703(.a(G381), .O(gate114inter8));
  nand2 gate1704(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1705(.a(s_165), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1706(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1707(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1708(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate2339(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate2340(.a(gate120inter0), .b(s_256), .O(gate120inter1));
  and2  gate2341(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate2342(.a(s_256), .O(gate120inter3));
  inv1  gate2343(.a(s_257), .O(gate120inter4));
  nand2 gate2344(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate2345(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate2346(.a(G392), .O(gate120inter7));
  inv1  gate2347(.a(G393), .O(gate120inter8));
  nand2 gate2348(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate2349(.a(s_257), .b(gate120inter3), .O(gate120inter10));
  nor2  gate2350(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate2351(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate2352(.a(gate120inter12), .b(gate120inter1), .O(G471));

  xor2  gate967(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate968(.a(gate121inter0), .b(s_60), .O(gate121inter1));
  and2  gate969(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate970(.a(s_60), .O(gate121inter3));
  inv1  gate971(.a(s_61), .O(gate121inter4));
  nand2 gate972(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate973(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate974(.a(G394), .O(gate121inter7));
  inv1  gate975(.a(G395), .O(gate121inter8));
  nand2 gate976(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate977(.a(s_61), .b(gate121inter3), .O(gate121inter10));
  nor2  gate978(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate979(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate980(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate897(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate898(.a(gate126inter0), .b(s_50), .O(gate126inter1));
  and2  gate899(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate900(.a(s_50), .O(gate126inter3));
  inv1  gate901(.a(s_51), .O(gate126inter4));
  nand2 gate902(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate903(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate904(.a(G404), .O(gate126inter7));
  inv1  gate905(.a(G405), .O(gate126inter8));
  nand2 gate906(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate907(.a(s_51), .b(gate126inter3), .O(gate126inter10));
  nor2  gate908(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate909(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate910(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate2353(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2354(.a(gate130inter0), .b(s_258), .O(gate130inter1));
  and2  gate2355(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2356(.a(s_258), .O(gate130inter3));
  inv1  gate2357(.a(s_259), .O(gate130inter4));
  nand2 gate2358(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2359(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2360(.a(G412), .O(gate130inter7));
  inv1  gate2361(.a(G413), .O(gate130inter8));
  nand2 gate2362(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2363(.a(s_259), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2364(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2365(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2366(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1793(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1794(.a(gate132inter0), .b(s_178), .O(gate132inter1));
  and2  gate1795(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1796(.a(s_178), .O(gate132inter3));
  inv1  gate1797(.a(s_179), .O(gate132inter4));
  nand2 gate1798(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1799(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1800(.a(G416), .O(gate132inter7));
  inv1  gate1801(.a(G417), .O(gate132inter8));
  nand2 gate1802(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1803(.a(s_179), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1804(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1805(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1806(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1261(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1262(.a(gate135inter0), .b(s_102), .O(gate135inter1));
  and2  gate1263(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1264(.a(s_102), .O(gate135inter3));
  inv1  gate1265(.a(s_103), .O(gate135inter4));
  nand2 gate1266(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1267(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1268(.a(G422), .O(gate135inter7));
  inv1  gate1269(.a(G423), .O(gate135inter8));
  nand2 gate1270(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1271(.a(s_103), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1272(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1273(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1274(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2367(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2368(.a(gate137inter0), .b(s_260), .O(gate137inter1));
  and2  gate2369(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2370(.a(s_260), .O(gate137inter3));
  inv1  gate2371(.a(s_261), .O(gate137inter4));
  nand2 gate2372(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2373(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2374(.a(G426), .O(gate137inter7));
  inv1  gate2375(.a(G429), .O(gate137inter8));
  nand2 gate2376(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2377(.a(s_261), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2378(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2379(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2380(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate827(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate828(.a(gate138inter0), .b(s_40), .O(gate138inter1));
  and2  gate829(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate830(.a(s_40), .O(gate138inter3));
  inv1  gate831(.a(s_41), .O(gate138inter4));
  nand2 gate832(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate833(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate834(.a(G432), .O(gate138inter7));
  inv1  gate835(.a(G435), .O(gate138inter8));
  nand2 gate836(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate837(.a(s_41), .b(gate138inter3), .O(gate138inter10));
  nor2  gate838(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate839(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate840(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1121(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1122(.a(gate144inter0), .b(s_82), .O(gate144inter1));
  and2  gate1123(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1124(.a(s_82), .O(gate144inter3));
  inv1  gate1125(.a(s_83), .O(gate144inter4));
  nand2 gate1126(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1127(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1128(.a(G468), .O(gate144inter7));
  inv1  gate1129(.a(G471), .O(gate144inter8));
  nand2 gate1130(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1131(.a(s_83), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1132(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1133(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1134(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1583(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1584(.a(gate145inter0), .b(s_148), .O(gate145inter1));
  and2  gate1585(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1586(.a(s_148), .O(gate145inter3));
  inv1  gate1587(.a(s_149), .O(gate145inter4));
  nand2 gate1588(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1589(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1590(.a(G474), .O(gate145inter7));
  inv1  gate1591(.a(G477), .O(gate145inter8));
  nand2 gate1592(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1593(.a(s_149), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1594(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1595(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1596(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate869(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate870(.a(gate147inter0), .b(s_46), .O(gate147inter1));
  and2  gate871(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate872(.a(s_46), .O(gate147inter3));
  inv1  gate873(.a(s_47), .O(gate147inter4));
  nand2 gate874(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate875(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate876(.a(G486), .O(gate147inter7));
  inv1  gate877(.a(G489), .O(gate147inter8));
  nand2 gate878(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate879(.a(s_47), .b(gate147inter3), .O(gate147inter10));
  nor2  gate880(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate881(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate882(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate911(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate912(.a(gate153inter0), .b(s_52), .O(gate153inter1));
  and2  gate913(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate914(.a(s_52), .O(gate153inter3));
  inv1  gate915(.a(s_53), .O(gate153inter4));
  nand2 gate916(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate917(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate918(.a(G426), .O(gate153inter7));
  inv1  gate919(.a(G522), .O(gate153inter8));
  nand2 gate920(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate921(.a(s_53), .b(gate153inter3), .O(gate153inter10));
  nor2  gate922(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate923(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate924(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1107(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1108(.a(gate154inter0), .b(s_80), .O(gate154inter1));
  and2  gate1109(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1110(.a(s_80), .O(gate154inter3));
  inv1  gate1111(.a(s_81), .O(gate154inter4));
  nand2 gate1112(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1113(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1114(.a(G429), .O(gate154inter7));
  inv1  gate1115(.a(G522), .O(gate154inter8));
  nand2 gate1116(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1117(.a(s_81), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1118(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1119(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1120(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1051(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1052(.a(gate165inter0), .b(s_72), .O(gate165inter1));
  and2  gate1053(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1054(.a(s_72), .O(gate165inter3));
  inv1  gate1055(.a(s_73), .O(gate165inter4));
  nand2 gate1056(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1057(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1058(.a(G462), .O(gate165inter7));
  inv1  gate1059(.a(G540), .O(gate165inter8));
  nand2 gate1060(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1061(.a(s_73), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1062(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1063(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1064(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1555(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1556(.a(gate167inter0), .b(s_144), .O(gate167inter1));
  and2  gate1557(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1558(.a(s_144), .O(gate167inter3));
  inv1  gate1559(.a(s_145), .O(gate167inter4));
  nand2 gate1560(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1561(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1562(.a(G468), .O(gate167inter7));
  inv1  gate1563(.a(G543), .O(gate167inter8));
  nand2 gate1564(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1565(.a(s_145), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1566(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1567(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1568(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1779(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1780(.a(gate168inter0), .b(s_176), .O(gate168inter1));
  and2  gate1781(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1782(.a(s_176), .O(gate168inter3));
  inv1  gate1783(.a(s_177), .O(gate168inter4));
  nand2 gate1784(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1785(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1786(.a(G471), .O(gate168inter7));
  inv1  gate1787(.a(G543), .O(gate168inter8));
  nand2 gate1788(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1789(.a(s_177), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1790(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1791(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1792(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1275(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1276(.a(gate170inter0), .b(s_104), .O(gate170inter1));
  and2  gate1277(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1278(.a(s_104), .O(gate170inter3));
  inv1  gate1279(.a(s_105), .O(gate170inter4));
  nand2 gate1280(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1281(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1282(.a(G477), .O(gate170inter7));
  inv1  gate1283(.a(G546), .O(gate170inter8));
  nand2 gate1284(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1285(.a(s_105), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1286(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1287(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1288(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2269(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2270(.a(gate172inter0), .b(s_246), .O(gate172inter1));
  and2  gate2271(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2272(.a(s_246), .O(gate172inter3));
  inv1  gate2273(.a(s_247), .O(gate172inter4));
  nand2 gate2274(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2275(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2276(.a(G483), .O(gate172inter7));
  inv1  gate2277(.a(G549), .O(gate172inter8));
  nand2 gate2278(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2279(.a(s_247), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2280(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2281(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2282(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2171(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2172(.a(gate173inter0), .b(s_232), .O(gate173inter1));
  and2  gate2173(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2174(.a(s_232), .O(gate173inter3));
  inv1  gate2175(.a(s_233), .O(gate173inter4));
  nand2 gate2176(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2177(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2178(.a(G486), .O(gate173inter7));
  inv1  gate2179(.a(G552), .O(gate173inter8));
  nand2 gate2180(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2181(.a(s_233), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2182(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2183(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2184(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1947(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1948(.a(gate174inter0), .b(s_200), .O(gate174inter1));
  and2  gate1949(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1950(.a(s_200), .O(gate174inter3));
  inv1  gate1951(.a(s_201), .O(gate174inter4));
  nand2 gate1952(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1953(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1954(.a(G489), .O(gate174inter7));
  inv1  gate1955(.a(G552), .O(gate174inter8));
  nand2 gate1956(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1957(.a(s_201), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1958(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1959(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1960(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate701(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate702(.a(gate177inter0), .b(s_22), .O(gate177inter1));
  and2  gate703(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate704(.a(s_22), .O(gate177inter3));
  inv1  gate705(.a(s_23), .O(gate177inter4));
  nand2 gate706(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate707(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate708(.a(G498), .O(gate177inter7));
  inv1  gate709(.a(G558), .O(gate177inter8));
  nand2 gate710(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate711(.a(s_23), .b(gate177inter3), .O(gate177inter10));
  nor2  gate712(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate713(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate714(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2283(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2284(.a(gate185inter0), .b(s_248), .O(gate185inter1));
  and2  gate2285(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2286(.a(s_248), .O(gate185inter3));
  inv1  gate2287(.a(s_249), .O(gate185inter4));
  nand2 gate2288(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2289(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2290(.a(G570), .O(gate185inter7));
  inv1  gate2291(.a(G571), .O(gate185inter8));
  nand2 gate2292(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2293(.a(s_249), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2294(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2295(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2296(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1037(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1038(.a(gate186inter0), .b(s_70), .O(gate186inter1));
  and2  gate1039(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1040(.a(s_70), .O(gate186inter3));
  inv1  gate1041(.a(s_71), .O(gate186inter4));
  nand2 gate1042(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1043(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1044(.a(G572), .O(gate186inter7));
  inv1  gate1045(.a(G573), .O(gate186inter8));
  nand2 gate1046(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1047(.a(s_71), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1048(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1049(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1050(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1177(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1178(.a(gate192inter0), .b(s_90), .O(gate192inter1));
  and2  gate1179(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1180(.a(s_90), .O(gate192inter3));
  inv1  gate1181(.a(s_91), .O(gate192inter4));
  nand2 gate1182(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1183(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1184(.a(G584), .O(gate192inter7));
  inv1  gate1185(.a(G585), .O(gate192inter8));
  nand2 gate1186(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1187(.a(s_91), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1188(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1189(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1190(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1807(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1808(.a(gate193inter0), .b(s_180), .O(gate193inter1));
  and2  gate1809(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1810(.a(s_180), .O(gate193inter3));
  inv1  gate1811(.a(s_181), .O(gate193inter4));
  nand2 gate1812(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1813(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1814(.a(G586), .O(gate193inter7));
  inv1  gate1815(.a(G587), .O(gate193inter8));
  nand2 gate1816(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1817(.a(s_181), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1818(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1819(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1820(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate2129(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2130(.a(gate194inter0), .b(s_226), .O(gate194inter1));
  and2  gate2131(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2132(.a(s_226), .O(gate194inter3));
  inv1  gate2133(.a(s_227), .O(gate194inter4));
  nand2 gate2134(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2135(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2136(.a(G588), .O(gate194inter7));
  inv1  gate2137(.a(G589), .O(gate194inter8));
  nand2 gate2138(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2139(.a(s_227), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2140(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2141(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2142(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2311(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2312(.a(gate195inter0), .b(s_252), .O(gate195inter1));
  and2  gate2313(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2314(.a(s_252), .O(gate195inter3));
  inv1  gate2315(.a(s_253), .O(gate195inter4));
  nand2 gate2316(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2317(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2318(.a(G590), .O(gate195inter7));
  inv1  gate2319(.a(G591), .O(gate195inter8));
  nand2 gate2320(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2321(.a(s_253), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2322(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2323(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2324(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate785(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate786(.a(gate197inter0), .b(s_34), .O(gate197inter1));
  and2  gate787(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate788(.a(s_34), .O(gate197inter3));
  inv1  gate789(.a(s_35), .O(gate197inter4));
  nand2 gate790(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate791(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate792(.a(G594), .O(gate197inter7));
  inv1  gate793(.a(G595), .O(gate197inter8));
  nand2 gate794(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate795(.a(s_35), .b(gate197inter3), .O(gate197inter10));
  nor2  gate796(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate797(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate798(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1499(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1500(.a(gate201inter0), .b(s_136), .O(gate201inter1));
  and2  gate1501(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1502(.a(s_136), .O(gate201inter3));
  inv1  gate1503(.a(s_137), .O(gate201inter4));
  nand2 gate1504(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1505(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1506(.a(G602), .O(gate201inter7));
  inv1  gate1507(.a(G607), .O(gate201inter8));
  nand2 gate1508(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1509(.a(s_137), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1510(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1511(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1512(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1891(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1892(.a(gate205inter0), .b(s_192), .O(gate205inter1));
  and2  gate1893(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1894(.a(s_192), .O(gate205inter3));
  inv1  gate1895(.a(s_193), .O(gate205inter4));
  nand2 gate1896(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1897(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1898(.a(G622), .O(gate205inter7));
  inv1  gate1899(.a(G627), .O(gate205inter8));
  nand2 gate1900(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1901(.a(s_193), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1902(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1903(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1904(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1849(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1850(.a(gate206inter0), .b(s_186), .O(gate206inter1));
  and2  gate1851(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1852(.a(s_186), .O(gate206inter3));
  inv1  gate1853(.a(s_187), .O(gate206inter4));
  nand2 gate1854(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1855(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1856(.a(G632), .O(gate206inter7));
  inv1  gate1857(.a(G637), .O(gate206inter8));
  nand2 gate1858(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1859(.a(s_187), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1860(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1861(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1862(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate925(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate926(.a(gate209inter0), .b(s_54), .O(gate209inter1));
  and2  gate927(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate928(.a(s_54), .O(gate209inter3));
  inv1  gate929(.a(s_55), .O(gate209inter4));
  nand2 gate930(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate931(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate932(.a(G602), .O(gate209inter7));
  inv1  gate933(.a(G666), .O(gate209inter8));
  nand2 gate934(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate935(.a(s_55), .b(gate209inter3), .O(gate209inter10));
  nor2  gate936(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate937(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate938(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1401(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1402(.a(gate211inter0), .b(s_122), .O(gate211inter1));
  and2  gate1403(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1404(.a(s_122), .O(gate211inter3));
  inv1  gate1405(.a(s_123), .O(gate211inter4));
  nand2 gate1406(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1407(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1408(.a(G612), .O(gate211inter7));
  inv1  gate1409(.a(G669), .O(gate211inter8));
  nand2 gate1410(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1411(.a(s_123), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1412(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1413(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1414(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate631(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate632(.a(gate218inter0), .b(s_12), .O(gate218inter1));
  and2  gate633(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate634(.a(s_12), .O(gate218inter3));
  inv1  gate635(.a(s_13), .O(gate218inter4));
  nand2 gate636(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate637(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate638(.a(G627), .O(gate218inter7));
  inv1  gate639(.a(G678), .O(gate218inter8));
  nand2 gate640(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate641(.a(s_13), .b(gate218inter3), .O(gate218inter10));
  nor2  gate642(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate643(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate644(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate2395(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate2396(.a(gate219inter0), .b(s_264), .O(gate219inter1));
  and2  gate2397(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate2398(.a(s_264), .O(gate219inter3));
  inv1  gate2399(.a(s_265), .O(gate219inter4));
  nand2 gate2400(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate2401(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate2402(.a(G632), .O(gate219inter7));
  inv1  gate2403(.a(G681), .O(gate219inter8));
  nand2 gate2404(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate2405(.a(s_265), .b(gate219inter3), .O(gate219inter10));
  nor2  gate2406(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate2407(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate2408(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1009(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1010(.a(gate222inter0), .b(s_66), .O(gate222inter1));
  and2  gate1011(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1012(.a(s_66), .O(gate222inter3));
  inv1  gate1013(.a(s_67), .O(gate222inter4));
  nand2 gate1014(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1015(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1016(.a(G632), .O(gate222inter7));
  inv1  gate1017(.a(G684), .O(gate222inter8));
  nand2 gate1018(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1019(.a(s_67), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1020(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1021(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1022(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1989(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1990(.a(gate227inter0), .b(s_206), .O(gate227inter1));
  and2  gate1991(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1992(.a(s_206), .O(gate227inter3));
  inv1  gate1993(.a(s_207), .O(gate227inter4));
  nand2 gate1994(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1995(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1996(.a(G694), .O(gate227inter7));
  inv1  gate1997(.a(G695), .O(gate227inter8));
  nand2 gate1998(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1999(.a(s_207), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2000(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2001(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2002(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1625(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1626(.a(gate231inter0), .b(s_154), .O(gate231inter1));
  and2  gate1627(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1628(.a(s_154), .O(gate231inter3));
  inv1  gate1629(.a(s_155), .O(gate231inter4));
  nand2 gate1630(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1631(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1632(.a(G702), .O(gate231inter7));
  inv1  gate1633(.a(G703), .O(gate231inter8));
  nand2 gate1634(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1635(.a(s_155), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1636(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1637(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1638(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2059(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2060(.a(gate233inter0), .b(s_216), .O(gate233inter1));
  and2  gate2061(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2062(.a(s_216), .O(gate233inter3));
  inv1  gate2063(.a(s_217), .O(gate233inter4));
  nand2 gate2064(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2065(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2066(.a(G242), .O(gate233inter7));
  inv1  gate2067(.a(G718), .O(gate233inter8));
  nand2 gate2068(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2069(.a(s_217), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2070(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2071(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2072(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1373(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1374(.a(gate242inter0), .b(s_118), .O(gate242inter1));
  and2  gate1375(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1376(.a(s_118), .O(gate242inter3));
  inv1  gate1377(.a(s_119), .O(gate242inter4));
  nand2 gate1378(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1379(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1380(.a(G718), .O(gate242inter7));
  inv1  gate1381(.a(G730), .O(gate242inter8));
  nand2 gate1382(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1383(.a(s_119), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1384(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1385(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1386(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate799(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate800(.a(gate245inter0), .b(s_36), .O(gate245inter1));
  and2  gate801(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate802(.a(s_36), .O(gate245inter3));
  inv1  gate803(.a(s_37), .O(gate245inter4));
  nand2 gate804(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate805(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate806(.a(G248), .O(gate245inter7));
  inv1  gate807(.a(G736), .O(gate245inter8));
  nand2 gate808(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate809(.a(s_37), .b(gate245inter3), .O(gate245inter10));
  nor2  gate810(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate811(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate812(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1317(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1318(.a(gate247inter0), .b(s_110), .O(gate247inter1));
  and2  gate1319(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1320(.a(s_110), .O(gate247inter3));
  inv1  gate1321(.a(s_111), .O(gate247inter4));
  nand2 gate1322(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1323(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1324(.a(G251), .O(gate247inter7));
  inv1  gate1325(.a(G739), .O(gate247inter8));
  nand2 gate1326(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1327(.a(s_111), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1328(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1329(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1330(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1359(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1360(.a(gate250inter0), .b(s_116), .O(gate250inter1));
  and2  gate1361(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1362(.a(s_116), .O(gate250inter3));
  inv1  gate1363(.a(s_117), .O(gate250inter4));
  nand2 gate1364(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1365(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1366(.a(G706), .O(gate250inter7));
  inv1  gate1367(.a(G742), .O(gate250inter8));
  nand2 gate1368(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1369(.a(s_117), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1370(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1371(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1372(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate603(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate604(.a(gate255inter0), .b(s_8), .O(gate255inter1));
  and2  gate605(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate606(.a(s_8), .O(gate255inter3));
  inv1  gate607(.a(s_9), .O(gate255inter4));
  nand2 gate608(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate609(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate610(.a(G263), .O(gate255inter7));
  inv1  gate611(.a(G751), .O(gate255inter8));
  nand2 gate612(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate613(.a(s_9), .b(gate255inter3), .O(gate255inter10));
  nor2  gate614(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate615(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate616(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1149(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1150(.a(gate256inter0), .b(s_86), .O(gate256inter1));
  and2  gate1151(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1152(.a(s_86), .O(gate256inter3));
  inv1  gate1153(.a(s_87), .O(gate256inter4));
  nand2 gate1154(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1155(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1156(.a(G715), .O(gate256inter7));
  inv1  gate1157(.a(G751), .O(gate256inter8));
  nand2 gate1158(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1159(.a(s_87), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1160(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1161(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1162(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1485(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1486(.a(gate259inter0), .b(s_134), .O(gate259inter1));
  and2  gate1487(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1488(.a(s_134), .O(gate259inter3));
  inv1  gate1489(.a(s_135), .O(gate259inter4));
  nand2 gate1490(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1491(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1492(.a(G758), .O(gate259inter7));
  inv1  gate1493(.a(G759), .O(gate259inter8));
  nand2 gate1494(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1495(.a(s_135), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1496(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1497(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1498(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2003(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2004(.a(gate261inter0), .b(s_208), .O(gate261inter1));
  and2  gate2005(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2006(.a(s_208), .O(gate261inter3));
  inv1  gate2007(.a(s_209), .O(gate261inter4));
  nand2 gate2008(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2009(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2010(.a(G762), .O(gate261inter7));
  inv1  gate2011(.a(G763), .O(gate261inter8));
  nand2 gate2012(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2013(.a(s_209), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2014(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2015(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2016(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1443(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1444(.a(gate262inter0), .b(s_128), .O(gate262inter1));
  and2  gate1445(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1446(.a(s_128), .O(gate262inter3));
  inv1  gate1447(.a(s_129), .O(gate262inter4));
  nand2 gate1448(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1449(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1450(.a(G764), .O(gate262inter7));
  inv1  gate1451(.a(G765), .O(gate262inter8));
  nand2 gate1452(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1453(.a(s_129), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1454(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1455(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1456(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2185(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2186(.a(gate263inter0), .b(s_234), .O(gate263inter1));
  and2  gate2187(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2188(.a(s_234), .O(gate263inter3));
  inv1  gate2189(.a(s_235), .O(gate263inter4));
  nand2 gate2190(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2191(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2192(.a(G766), .O(gate263inter7));
  inv1  gate2193(.a(G767), .O(gate263inter8));
  nand2 gate2194(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2195(.a(s_235), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2196(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2197(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2198(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2199(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2200(.a(gate265inter0), .b(s_236), .O(gate265inter1));
  and2  gate2201(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2202(.a(s_236), .O(gate265inter3));
  inv1  gate2203(.a(s_237), .O(gate265inter4));
  nand2 gate2204(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2205(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2206(.a(G642), .O(gate265inter7));
  inv1  gate2207(.a(G770), .O(gate265inter8));
  nand2 gate2208(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2209(.a(s_237), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2210(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2211(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2212(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1205(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1206(.a(gate266inter0), .b(s_94), .O(gate266inter1));
  and2  gate1207(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1208(.a(s_94), .O(gate266inter3));
  inv1  gate1209(.a(s_95), .O(gate266inter4));
  nand2 gate1210(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1211(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1212(.a(G645), .O(gate266inter7));
  inv1  gate1213(.a(G773), .O(gate266inter8));
  nand2 gate1214(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1215(.a(s_95), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1216(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1217(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1218(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate995(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate996(.a(gate268inter0), .b(s_64), .O(gate268inter1));
  and2  gate997(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate998(.a(s_64), .O(gate268inter3));
  inv1  gate999(.a(s_65), .O(gate268inter4));
  nand2 gate1000(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1001(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1002(.a(G651), .O(gate268inter7));
  inv1  gate1003(.a(G779), .O(gate268inter8));
  nand2 gate1004(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1005(.a(s_65), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1006(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1007(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1008(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1877(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1878(.a(gate273inter0), .b(s_190), .O(gate273inter1));
  and2  gate1879(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1880(.a(s_190), .O(gate273inter3));
  inv1  gate1881(.a(s_191), .O(gate273inter4));
  nand2 gate1882(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1883(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1884(.a(G642), .O(gate273inter7));
  inv1  gate1885(.a(G794), .O(gate273inter8));
  nand2 gate1886(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1887(.a(s_191), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1888(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1889(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1890(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate673(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate674(.a(gate274inter0), .b(s_18), .O(gate274inter1));
  and2  gate675(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate676(.a(s_18), .O(gate274inter3));
  inv1  gate677(.a(s_19), .O(gate274inter4));
  nand2 gate678(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate679(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate680(.a(G770), .O(gate274inter7));
  inv1  gate681(.a(G794), .O(gate274inter8));
  nand2 gate682(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate683(.a(s_19), .b(gate274inter3), .O(gate274inter10));
  nor2  gate684(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate685(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate686(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1863(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1864(.a(gate275inter0), .b(s_188), .O(gate275inter1));
  and2  gate1865(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1866(.a(s_188), .O(gate275inter3));
  inv1  gate1867(.a(s_189), .O(gate275inter4));
  nand2 gate1868(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1869(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1870(.a(G645), .O(gate275inter7));
  inv1  gate1871(.a(G797), .O(gate275inter8));
  nand2 gate1872(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1873(.a(s_189), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1874(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1875(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1876(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate953(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate954(.a(gate278inter0), .b(s_58), .O(gate278inter1));
  and2  gate955(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate956(.a(s_58), .O(gate278inter3));
  inv1  gate957(.a(s_59), .O(gate278inter4));
  nand2 gate958(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate959(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate960(.a(G776), .O(gate278inter7));
  inv1  gate961(.a(G800), .O(gate278inter8));
  nand2 gate962(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate963(.a(s_59), .b(gate278inter3), .O(gate278inter10));
  nor2  gate964(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate965(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate966(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate589(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate590(.a(gate284inter0), .b(s_6), .O(gate284inter1));
  and2  gate591(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate592(.a(s_6), .O(gate284inter3));
  inv1  gate593(.a(s_7), .O(gate284inter4));
  nand2 gate594(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate595(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate596(.a(G785), .O(gate284inter7));
  inv1  gate597(.a(G809), .O(gate284inter8));
  nand2 gate598(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate599(.a(s_7), .b(gate284inter3), .O(gate284inter10));
  nor2  gate600(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate601(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate602(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1415(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1416(.a(gate286inter0), .b(s_124), .O(gate286inter1));
  and2  gate1417(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1418(.a(s_124), .O(gate286inter3));
  inv1  gate1419(.a(s_125), .O(gate286inter4));
  nand2 gate1420(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1421(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1422(.a(G788), .O(gate286inter7));
  inv1  gate1423(.a(G812), .O(gate286inter8));
  nand2 gate1424(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1425(.a(s_125), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1426(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1427(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1428(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1513(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1514(.a(gate287inter0), .b(s_138), .O(gate287inter1));
  and2  gate1515(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1516(.a(s_138), .O(gate287inter3));
  inv1  gate1517(.a(s_139), .O(gate287inter4));
  nand2 gate1518(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1519(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1520(.a(G663), .O(gate287inter7));
  inv1  gate1521(.a(G815), .O(gate287inter8));
  nand2 gate1522(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1523(.a(s_139), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1524(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1525(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1526(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1233(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1234(.a(gate289inter0), .b(s_98), .O(gate289inter1));
  and2  gate1235(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1236(.a(s_98), .O(gate289inter3));
  inv1  gate1237(.a(s_99), .O(gate289inter4));
  nand2 gate1238(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1239(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1240(.a(G818), .O(gate289inter7));
  inv1  gate1241(.a(G819), .O(gate289inter8));
  nand2 gate1242(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1243(.a(s_99), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1244(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1245(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1246(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1135(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1136(.a(gate290inter0), .b(s_84), .O(gate290inter1));
  and2  gate1137(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1138(.a(s_84), .O(gate290inter3));
  inv1  gate1139(.a(s_85), .O(gate290inter4));
  nand2 gate1140(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1141(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1142(.a(G820), .O(gate290inter7));
  inv1  gate1143(.a(G821), .O(gate290inter8));
  nand2 gate1144(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1145(.a(s_85), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1146(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1147(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1148(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1667(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1668(.a(gate293inter0), .b(s_160), .O(gate293inter1));
  and2  gate1669(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1670(.a(s_160), .O(gate293inter3));
  inv1  gate1671(.a(s_161), .O(gate293inter4));
  nand2 gate1672(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1673(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1674(.a(G828), .O(gate293inter7));
  inv1  gate1675(.a(G829), .O(gate293inter8));
  nand2 gate1676(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1677(.a(s_161), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1678(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1679(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1680(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate547(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate548(.a(gate389inter0), .b(s_0), .O(gate389inter1));
  and2  gate549(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate550(.a(s_0), .O(gate389inter3));
  inv1  gate551(.a(s_1), .O(gate389inter4));
  nand2 gate552(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate553(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate554(.a(G3), .O(gate389inter7));
  inv1  gate555(.a(G1042), .O(gate389inter8));
  nand2 gate556(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate557(.a(s_1), .b(gate389inter3), .O(gate389inter10));
  nor2  gate558(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate559(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate560(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1919(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1920(.a(gate390inter0), .b(s_196), .O(gate390inter1));
  and2  gate1921(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1922(.a(s_196), .O(gate390inter3));
  inv1  gate1923(.a(s_197), .O(gate390inter4));
  nand2 gate1924(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1925(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1926(.a(G4), .O(gate390inter7));
  inv1  gate1927(.a(G1045), .O(gate390inter8));
  nand2 gate1928(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1929(.a(s_197), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1930(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1931(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1932(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1905(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1906(.a(gate391inter0), .b(s_194), .O(gate391inter1));
  and2  gate1907(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1908(.a(s_194), .O(gate391inter3));
  inv1  gate1909(.a(s_195), .O(gate391inter4));
  nand2 gate1910(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1911(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1912(.a(G5), .O(gate391inter7));
  inv1  gate1913(.a(G1048), .O(gate391inter8));
  nand2 gate1914(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1915(.a(s_195), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1916(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1917(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1918(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1765(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1766(.a(gate393inter0), .b(s_174), .O(gate393inter1));
  and2  gate1767(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1768(.a(s_174), .O(gate393inter3));
  inv1  gate1769(.a(s_175), .O(gate393inter4));
  nand2 gate1770(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1771(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1772(.a(G7), .O(gate393inter7));
  inv1  gate1773(.a(G1054), .O(gate393inter8));
  nand2 gate1774(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1775(.a(s_175), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1776(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1777(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1778(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate771(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate772(.a(gate394inter0), .b(s_32), .O(gate394inter1));
  and2  gate773(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate774(.a(s_32), .O(gate394inter3));
  inv1  gate775(.a(s_33), .O(gate394inter4));
  nand2 gate776(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate777(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate778(.a(G8), .O(gate394inter7));
  inv1  gate779(.a(G1057), .O(gate394inter8));
  nand2 gate780(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate781(.a(s_33), .b(gate394inter3), .O(gate394inter10));
  nor2  gate782(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate783(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate784(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1471(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1472(.a(gate398inter0), .b(s_132), .O(gate398inter1));
  and2  gate1473(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1474(.a(s_132), .O(gate398inter3));
  inv1  gate1475(.a(s_133), .O(gate398inter4));
  nand2 gate1476(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1477(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1478(.a(G12), .O(gate398inter7));
  inv1  gate1479(.a(G1069), .O(gate398inter8));
  nand2 gate1480(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1481(.a(s_133), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1482(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1483(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1484(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1835(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1836(.a(gate400inter0), .b(s_184), .O(gate400inter1));
  and2  gate1837(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1838(.a(s_184), .O(gate400inter3));
  inv1  gate1839(.a(s_185), .O(gate400inter4));
  nand2 gate1840(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1841(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1842(.a(G14), .O(gate400inter7));
  inv1  gate1843(.a(G1075), .O(gate400inter8));
  nand2 gate1844(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1845(.a(s_185), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1846(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1847(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1848(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate841(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate842(.a(gate401inter0), .b(s_42), .O(gate401inter1));
  and2  gate843(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate844(.a(s_42), .O(gate401inter3));
  inv1  gate845(.a(s_43), .O(gate401inter4));
  nand2 gate846(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate847(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate848(.a(G15), .O(gate401inter7));
  inv1  gate849(.a(G1078), .O(gate401inter8));
  nand2 gate850(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate851(.a(s_43), .b(gate401inter3), .O(gate401inter10));
  nor2  gate852(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate853(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate854(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate645(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate646(.a(gate402inter0), .b(s_14), .O(gate402inter1));
  and2  gate647(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate648(.a(s_14), .O(gate402inter3));
  inv1  gate649(.a(s_15), .O(gate402inter4));
  nand2 gate650(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate651(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate652(.a(G16), .O(gate402inter7));
  inv1  gate653(.a(G1081), .O(gate402inter8));
  nand2 gate654(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate655(.a(s_15), .b(gate402inter3), .O(gate402inter10));
  nor2  gate656(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate657(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate658(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate2087(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2088(.a(gate403inter0), .b(s_220), .O(gate403inter1));
  and2  gate2089(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2090(.a(s_220), .O(gate403inter3));
  inv1  gate2091(.a(s_221), .O(gate403inter4));
  nand2 gate2092(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2093(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2094(.a(G17), .O(gate403inter7));
  inv1  gate2095(.a(G1084), .O(gate403inter8));
  nand2 gate2096(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2097(.a(s_221), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2098(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2099(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2100(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1387(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1388(.a(gate404inter0), .b(s_120), .O(gate404inter1));
  and2  gate1389(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1390(.a(s_120), .O(gate404inter3));
  inv1  gate1391(.a(s_121), .O(gate404inter4));
  nand2 gate1392(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1393(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1394(.a(G18), .O(gate404inter7));
  inv1  gate1395(.a(G1087), .O(gate404inter8));
  nand2 gate1396(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1397(.a(s_121), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1398(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1399(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1400(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2409(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2410(.a(gate406inter0), .b(s_266), .O(gate406inter1));
  and2  gate2411(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2412(.a(s_266), .O(gate406inter3));
  inv1  gate2413(.a(s_267), .O(gate406inter4));
  nand2 gate2414(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2415(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2416(.a(G20), .O(gate406inter7));
  inv1  gate2417(.a(G1093), .O(gate406inter8));
  nand2 gate2418(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2419(.a(s_267), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2420(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2421(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2422(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1331(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1332(.a(gate407inter0), .b(s_112), .O(gate407inter1));
  and2  gate1333(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1334(.a(s_112), .O(gate407inter3));
  inv1  gate1335(.a(s_113), .O(gate407inter4));
  nand2 gate1336(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1337(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1338(.a(G21), .O(gate407inter7));
  inv1  gate1339(.a(G1096), .O(gate407inter8));
  nand2 gate1340(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1341(.a(s_113), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1342(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1343(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1344(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1737(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1738(.a(gate408inter0), .b(s_170), .O(gate408inter1));
  and2  gate1739(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1740(.a(s_170), .O(gate408inter3));
  inv1  gate1741(.a(s_171), .O(gate408inter4));
  nand2 gate1742(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1743(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1744(.a(G22), .O(gate408inter7));
  inv1  gate1745(.a(G1099), .O(gate408inter8));
  nand2 gate1746(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1747(.a(s_171), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1748(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1749(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1750(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1023(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1024(.a(gate413inter0), .b(s_68), .O(gate413inter1));
  and2  gate1025(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1026(.a(s_68), .O(gate413inter3));
  inv1  gate1027(.a(s_69), .O(gate413inter4));
  nand2 gate1028(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1029(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1030(.a(G27), .O(gate413inter7));
  inv1  gate1031(.a(G1114), .O(gate413inter8));
  nand2 gate1032(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1033(.a(s_69), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1034(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1035(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1036(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1653(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1654(.a(gate415inter0), .b(s_158), .O(gate415inter1));
  and2  gate1655(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1656(.a(s_158), .O(gate415inter3));
  inv1  gate1657(.a(s_159), .O(gate415inter4));
  nand2 gate1658(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1659(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1660(.a(G29), .O(gate415inter7));
  inv1  gate1661(.a(G1120), .O(gate415inter8));
  nand2 gate1662(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1663(.a(s_159), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1664(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1665(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1666(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1065(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1066(.a(gate420inter0), .b(s_74), .O(gate420inter1));
  and2  gate1067(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1068(.a(s_74), .O(gate420inter3));
  inv1  gate1069(.a(s_75), .O(gate420inter4));
  nand2 gate1070(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1071(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1072(.a(G1036), .O(gate420inter7));
  inv1  gate1073(.a(G1132), .O(gate420inter8));
  nand2 gate1074(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1075(.a(s_75), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1076(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1077(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1078(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2031(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2032(.a(gate421inter0), .b(s_212), .O(gate421inter1));
  and2  gate2033(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2034(.a(s_212), .O(gate421inter3));
  inv1  gate2035(.a(s_213), .O(gate421inter4));
  nand2 gate2036(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2037(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2038(.a(G2), .O(gate421inter7));
  inv1  gate2039(.a(G1135), .O(gate421inter8));
  nand2 gate2040(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2041(.a(s_213), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2042(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2043(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2044(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2073(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2074(.a(gate424inter0), .b(s_218), .O(gate424inter1));
  and2  gate2075(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2076(.a(s_218), .O(gate424inter3));
  inv1  gate2077(.a(s_219), .O(gate424inter4));
  nand2 gate2078(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2079(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2080(.a(G1042), .O(gate424inter7));
  inv1  gate2081(.a(G1138), .O(gate424inter8));
  nand2 gate2082(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2083(.a(s_219), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2084(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2085(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2086(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2227(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2228(.a(gate432inter0), .b(s_240), .O(gate432inter1));
  and2  gate2229(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2230(.a(s_240), .O(gate432inter3));
  inv1  gate2231(.a(s_241), .O(gate432inter4));
  nand2 gate2232(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2233(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2234(.a(G1054), .O(gate432inter7));
  inv1  gate2235(.a(G1150), .O(gate432inter8));
  nand2 gate2236(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2237(.a(s_241), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2238(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2239(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2240(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate687(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate688(.a(gate434inter0), .b(s_20), .O(gate434inter1));
  and2  gate689(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate690(.a(s_20), .O(gate434inter3));
  inv1  gate691(.a(s_21), .O(gate434inter4));
  nand2 gate692(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate693(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate694(.a(G1057), .O(gate434inter7));
  inv1  gate695(.a(G1153), .O(gate434inter8));
  nand2 gate696(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate697(.a(s_21), .b(gate434inter3), .O(gate434inter10));
  nor2  gate698(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate699(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate700(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate659(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate660(.a(gate436inter0), .b(s_16), .O(gate436inter1));
  and2  gate661(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate662(.a(s_16), .O(gate436inter3));
  inv1  gate663(.a(s_17), .O(gate436inter4));
  nand2 gate664(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate665(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate666(.a(G1060), .O(gate436inter7));
  inv1  gate667(.a(G1156), .O(gate436inter8));
  nand2 gate668(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate669(.a(s_17), .b(gate436inter3), .O(gate436inter10));
  nor2  gate670(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate671(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate672(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate883(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate884(.a(gate437inter0), .b(s_48), .O(gate437inter1));
  and2  gate885(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate886(.a(s_48), .O(gate437inter3));
  inv1  gate887(.a(s_49), .O(gate437inter4));
  nand2 gate888(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate889(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate890(.a(G10), .O(gate437inter7));
  inv1  gate891(.a(G1159), .O(gate437inter8));
  nand2 gate892(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate893(.a(s_49), .b(gate437inter3), .O(gate437inter10));
  nor2  gate894(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate895(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate896(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1079(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1080(.a(gate443inter0), .b(s_76), .O(gate443inter1));
  and2  gate1081(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1082(.a(s_76), .O(gate443inter3));
  inv1  gate1083(.a(s_77), .O(gate443inter4));
  nand2 gate1084(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1085(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1086(.a(G13), .O(gate443inter7));
  inv1  gate1087(.a(G1168), .O(gate443inter8));
  nand2 gate1088(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1089(.a(s_77), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1090(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1091(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1092(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1933(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1934(.a(gate444inter0), .b(s_198), .O(gate444inter1));
  and2  gate1935(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1936(.a(s_198), .O(gate444inter3));
  inv1  gate1937(.a(s_199), .O(gate444inter4));
  nand2 gate1938(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1939(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1940(.a(G1072), .O(gate444inter7));
  inv1  gate1941(.a(G1168), .O(gate444inter8));
  nand2 gate1942(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1943(.a(s_199), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1944(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1945(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1946(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1093(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1094(.a(gate451inter0), .b(s_78), .O(gate451inter1));
  and2  gate1095(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1096(.a(s_78), .O(gate451inter3));
  inv1  gate1097(.a(s_79), .O(gate451inter4));
  nand2 gate1098(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1099(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1100(.a(G17), .O(gate451inter7));
  inv1  gate1101(.a(G1180), .O(gate451inter8));
  nand2 gate1102(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1103(.a(s_79), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1104(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1105(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1106(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate729(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate730(.a(gate452inter0), .b(s_26), .O(gate452inter1));
  and2  gate731(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate732(.a(s_26), .O(gate452inter3));
  inv1  gate733(.a(s_27), .O(gate452inter4));
  nand2 gate734(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate735(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate736(.a(G1084), .O(gate452inter7));
  inv1  gate737(.a(G1180), .O(gate452inter8));
  nand2 gate738(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate739(.a(s_27), .b(gate452inter3), .O(gate452inter10));
  nor2  gate740(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate741(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate742(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate715(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate716(.a(gate456inter0), .b(s_24), .O(gate456inter1));
  and2  gate717(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate718(.a(s_24), .O(gate456inter3));
  inv1  gate719(.a(s_25), .O(gate456inter4));
  nand2 gate720(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate721(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate722(.a(G1090), .O(gate456inter7));
  inv1  gate723(.a(G1186), .O(gate456inter8));
  nand2 gate724(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate725(.a(s_25), .b(gate456inter3), .O(gate456inter10));
  nor2  gate726(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate727(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate728(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1345(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1346(.a(gate458inter0), .b(s_114), .O(gate458inter1));
  and2  gate1347(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1348(.a(s_114), .O(gate458inter3));
  inv1  gate1349(.a(s_115), .O(gate458inter4));
  nand2 gate1350(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1351(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1352(.a(G1093), .O(gate458inter7));
  inv1  gate1353(.a(G1189), .O(gate458inter8));
  nand2 gate1354(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1355(.a(s_115), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1356(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1357(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1358(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate743(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate744(.a(gate459inter0), .b(s_28), .O(gate459inter1));
  and2  gate745(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate746(.a(s_28), .O(gate459inter3));
  inv1  gate747(.a(s_29), .O(gate459inter4));
  nand2 gate748(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate749(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate750(.a(G21), .O(gate459inter7));
  inv1  gate751(.a(G1192), .O(gate459inter8));
  nand2 gate752(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate753(.a(s_29), .b(gate459inter3), .O(gate459inter10));
  nor2  gate754(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate755(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate756(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate757(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate758(.a(gate463inter0), .b(s_30), .O(gate463inter1));
  and2  gate759(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate760(.a(s_30), .O(gate463inter3));
  inv1  gate761(.a(s_31), .O(gate463inter4));
  nand2 gate762(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate763(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate764(.a(G23), .O(gate463inter7));
  inv1  gate765(.a(G1198), .O(gate463inter8));
  nand2 gate766(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate767(.a(s_31), .b(gate463inter3), .O(gate463inter10));
  nor2  gate768(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate769(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate770(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate855(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate856(.a(gate466inter0), .b(s_44), .O(gate466inter1));
  and2  gate857(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate858(.a(s_44), .O(gate466inter3));
  inv1  gate859(.a(s_45), .O(gate466inter4));
  nand2 gate860(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate861(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate862(.a(G1105), .O(gate466inter7));
  inv1  gate863(.a(G1201), .O(gate466inter8));
  nand2 gate864(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate865(.a(s_45), .b(gate466inter3), .O(gate466inter10));
  nor2  gate866(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate867(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate868(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1541(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1542(.a(gate471inter0), .b(s_142), .O(gate471inter1));
  and2  gate1543(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1544(.a(s_142), .O(gate471inter3));
  inv1  gate1545(.a(s_143), .O(gate471inter4));
  nand2 gate1546(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1547(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1548(.a(G27), .O(gate471inter7));
  inv1  gate1549(.a(G1210), .O(gate471inter8));
  nand2 gate1550(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1551(.a(s_143), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1552(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1553(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1554(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1191(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1192(.a(gate475inter0), .b(s_92), .O(gate475inter1));
  and2  gate1193(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1194(.a(s_92), .O(gate475inter3));
  inv1  gate1195(.a(s_93), .O(gate475inter4));
  nand2 gate1196(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1197(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1198(.a(G29), .O(gate475inter7));
  inv1  gate1199(.a(G1216), .O(gate475inter8));
  nand2 gate1200(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1201(.a(s_93), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1202(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1203(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1204(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1639(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1640(.a(gate476inter0), .b(s_156), .O(gate476inter1));
  and2  gate1641(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1642(.a(s_156), .O(gate476inter3));
  inv1  gate1643(.a(s_157), .O(gate476inter4));
  nand2 gate1644(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1645(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1646(.a(G1120), .O(gate476inter7));
  inv1  gate1647(.a(G1216), .O(gate476inter8));
  nand2 gate1648(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1649(.a(s_157), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1650(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1651(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1652(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2157(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2158(.a(gate480inter0), .b(s_230), .O(gate480inter1));
  and2  gate2159(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2160(.a(s_230), .O(gate480inter3));
  inv1  gate2161(.a(s_231), .O(gate480inter4));
  nand2 gate2162(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2163(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2164(.a(G1126), .O(gate480inter7));
  inv1  gate2165(.a(G1222), .O(gate480inter8));
  nand2 gate2166(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2167(.a(s_231), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2168(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2169(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2170(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate981(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate982(.a(gate502inter0), .b(s_62), .O(gate502inter1));
  and2  gate983(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate984(.a(s_62), .O(gate502inter3));
  inv1  gate985(.a(s_63), .O(gate502inter4));
  nand2 gate986(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate987(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate988(.a(G1266), .O(gate502inter7));
  inv1  gate989(.a(G1267), .O(gate502inter8));
  nand2 gate990(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate991(.a(s_63), .b(gate502inter3), .O(gate502inter10));
  nor2  gate992(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate993(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate994(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1821(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1822(.a(gate514inter0), .b(s_182), .O(gate514inter1));
  and2  gate1823(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1824(.a(s_182), .O(gate514inter3));
  inv1  gate1825(.a(s_183), .O(gate514inter4));
  nand2 gate1826(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1827(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1828(.a(G1290), .O(gate514inter7));
  inv1  gate1829(.a(G1291), .O(gate514inter8));
  nand2 gate1830(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1831(.a(s_183), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1832(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1833(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1834(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule