module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381, s_382, s_383, s_384, s_385, s_386, s_387, s_388, s_389, s_390, s_391;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1317(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1318(.a(gate9inter0), .b(s_110), .O(gate9inter1));
  and2  gate1319(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1320(.a(s_110), .O(gate9inter3));
  inv1  gate1321(.a(s_111), .O(gate9inter4));
  nand2 gate1322(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1323(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1324(.a(G1), .O(gate9inter7));
  inv1  gate1325(.a(G2), .O(gate9inter8));
  nand2 gate1326(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1327(.a(s_111), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1328(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1329(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1330(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1051(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1052(.a(gate10inter0), .b(s_72), .O(gate10inter1));
  and2  gate1053(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1054(.a(s_72), .O(gate10inter3));
  inv1  gate1055(.a(s_73), .O(gate10inter4));
  nand2 gate1056(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1057(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1058(.a(G3), .O(gate10inter7));
  inv1  gate1059(.a(G4), .O(gate10inter8));
  nand2 gate1060(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1061(.a(s_73), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1062(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1063(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1064(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2619(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2620(.a(gate12inter0), .b(s_296), .O(gate12inter1));
  and2  gate2621(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2622(.a(s_296), .O(gate12inter3));
  inv1  gate2623(.a(s_297), .O(gate12inter4));
  nand2 gate2624(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2625(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2626(.a(G7), .O(gate12inter7));
  inv1  gate2627(.a(G8), .O(gate12inter8));
  nand2 gate2628(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2629(.a(s_297), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2630(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2631(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2632(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2871(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2872(.a(gate15inter0), .b(s_332), .O(gate15inter1));
  and2  gate2873(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2874(.a(s_332), .O(gate15inter3));
  inv1  gate2875(.a(s_333), .O(gate15inter4));
  nand2 gate2876(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2877(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2878(.a(G13), .O(gate15inter7));
  inv1  gate2879(.a(G14), .O(gate15inter8));
  nand2 gate2880(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2881(.a(s_333), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2882(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2883(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2884(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1205(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1206(.a(gate17inter0), .b(s_94), .O(gate17inter1));
  and2  gate1207(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1208(.a(s_94), .O(gate17inter3));
  inv1  gate1209(.a(s_95), .O(gate17inter4));
  nand2 gate1210(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1211(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1212(.a(G17), .O(gate17inter7));
  inv1  gate1213(.a(G18), .O(gate17inter8));
  nand2 gate1214(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1215(.a(s_95), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1216(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1217(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1218(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate953(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate954(.a(gate19inter0), .b(s_58), .O(gate19inter1));
  and2  gate955(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate956(.a(s_58), .O(gate19inter3));
  inv1  gate957(.a(s_59), .O(gate19inter4));
  nand2 gate958(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate959(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate960(.a(G21), .O(gate19inter7));
  inv1  gate961(.a(G22), .O(gate19inter8));
  nand2 gate962(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate963(.a(s_59), .b(gate19inter3), .O(gate19inter10));
  nor2  gate964(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate965(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate966(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1681(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1682(.a(gate20inter0), .b(s_162), .O(gate20inter1));
  and2  gate1683(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1684(.a(s_162), .O(gate20inter3));
  inv1  gate1685(.a(s_163), .O(gate20inter4));
  nand2 gate1686(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1687(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1688(.a(G23), .O(gate20inter7));
  inv1  gate1689(.a(G24), .O(gate20inter8));
  nand2 gate1690(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1691(.a(s_163), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1692(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1693(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1694(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2955(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2956(.a(gate23inter0), .b(s_344), .O(gate23inter1));
  and2  gate2957(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2958(.a(s_344), .O(gate23inter3));
  inv1  gate2959(.a(s_345), .O(gate23inter4));
  nand2 gate2960(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2961(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2962(.a(G29), .O(gate23inter7));
  inv1  gate2963(.a(G30), .O(gate23inter8));
  nand2 gate2964(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2965(.a(s_345), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2966(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2967(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2968(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2283(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2284(.a(gate25inter0), .b(s_248), .O(gate25inter1));
  and2  gate2285(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2286(.a(s_248), .O(gate25inter3));
  inv1  gate2287(.a(s_249), .O(gate25inter4));
  nand2 gate2288(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2289(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2290(.a(G1), .O(gate25inter7));
  inv1  gate2291(.a(G5), .O(gate25inter8));
  nand2 gate2292(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2293(.a(s_249), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2294(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2295(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2296(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2003(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2004(.a(gate28inter0), .b(s_208), .O(gate28inter1));
  and2  gate2005(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2006(.a(s_208), .O(gate28inter3));
  inv1  gate2007(.a(s_209), .O(gate28inter4));
  nand2 gate2008(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2009(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2010(.a(G10), .O(gate28inter7));
  inv1  gate2011(.a(G14), .O(gate28inter8));
  nand2 gate2012(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2013(.a(s_209), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2014(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2015(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2016(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2199(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2200(.a(gate29inter0), .b(s_236), .O(gate29inter1));
  and2  gate2201(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2202(.a(s_236), .O(gate29inter3));
  inv1  gate2203(.a(s_237), .O(gate29inter4));
  nand2 gate2204(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2205(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2206(.a(G3), .O(gate29inter7));
  inv1  gate2207(.a(G7), .O(gate29inter8));
  nand2 gate2208(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2209(.a(s_237), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2210(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2211(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2212(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate2787(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate2788(.a(gate30inter0), .b(s_320), .O(gate30inter1));
  and2  gate2789(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate2790(.a(s_320), .O(gate30inter3));
  inv1  gate2791(.a(s_321), .O(gate30inter4));
  nand2 gate2792(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate2793(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate2794(.a(G11), .O(gate30inter7));
  inv1  gate2795(.a(G15), .O(gate30inter8));
  nand2 gate2796(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate2797(.a(s_321), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2798(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2799(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2800(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1331(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1332(.a(gate31inter0), .b(s_112), .O(gate31inter1));
  and2  gate1333(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1334(.a(s_112), .O(gate31inter3));
  inv1  gate1335(.a(s_113), .O(gate31inter4));
  nand2 gate1336(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1337(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1338(.a(G4), .O(gate31inter7));
  inv1  gate1339(.a(G8), .O(gate31inter8));
  nand2 gate1340(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1341(.a(s_113), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1342(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1343(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1344(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate813(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate814(.a(gate32inter0), .b(s_38), .O(gate32inter1));
  and2  gate815(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate816(.a(s_38), .O(gate32inter3));
  inv1  gate817(.a(s_39), .O(gate32inter4));
  nand2 gate818(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate819(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate820(.a(G12), .O(gate32inter7));
  inv1  gate821(.a(G16), .O(gate32inter8));
  nand2 gate822(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate823(.a(s_39), .b(gate32inter3), .O(gate32inter10));
  nor2  gate824(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate825(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate826(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1821(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1822(.a(gate36inter0), .b(s_182), .O(gate36inter1));
  and2  gate1823(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1824(.a(s_182), .O(gate36inter3));
  inv1  gate1825(.a(s_183), .O(gate36inter4));
  nand2 gate1826(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1827(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1828(.a(G26), .O(gate36inter7));
  inv1  gate1829(.a(G30), .O(gate36inter8));
  nand2 gate1830(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1831(.a(s_183), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1832(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1833(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1834(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1891(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1892(.a(gate38inter0), .b(s_192), .O(gate38inter1));
  and2  gate1893(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1894(.a(s_192), .O(gate38inter3));
  inv1  gate1895(.a(s_193), .O(gate38inter4));
  nand2 gate1896(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1897(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1898(.a(G27), .O(gate38inter7));
  inv1  gate1899(.a(G31), .O(gate38inter8));
  nand2 gate1900(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1901(.a(s_193), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1902(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1903(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1904(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate3221(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate3222(.a(gate44inter0), .b(s_382), .O(gate44inter1));
  and2  gate3223(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate3224(.a(s_382), .O(gate44inter3));
  inv1  gate3225(.a(s_383), .O(gate44inter4));
  nand2 gate3226(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate3227(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate3228(.a(G4), .O(gate44inter7));
  inv1  gate3229(.a(G269), .O(gate44inter8));
  nand2 gate3230(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate3231(.a(s_383), .b(gate44inter3), .O(gate44inter10));
  nor2  gate3232(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate3233(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate3234(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1709(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1710(.a(gate45inter0), .b(s_166), .O(gate45inter1));
  and2  gate1711(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1712(.a(s_166), .O(gate45inter3));
  inv1  gate1713(.a(s_167), .O(gate45inter4));
  nand2 gate1714(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1715(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1716(.a(G5), .O(gate45inter7));
  inv1  gate1717(.a(G272), .O(gate45inter8));
  nand2 gate1718(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1719(.a(s_167), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1720(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1721(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1722(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1933(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1934(.a(gate46inter0), .b(s_198), .O(gate46inter1));
  and2  gate1935(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1936(.a(s_198), .O(gate46inter3));
  inv1  gate1937(.a(s_199), .O(gate46inter4));
  nand2 gate1938(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1939(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1940(.a(G6), .O(gate46inter7));
  inv1  gate1941(.a(G272), .O(gate46inter8));
  nand2 gate1942(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1943(.a(s_199), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1944(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1945(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1946(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2437(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2438(.a(gate48inter0), .b(s_270), .O(gate48inter1));
  and2  gate2439(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2440(.a(s_270), .O(gate48inter3));
  inv1  gate2441(.a(s_271), .O(gate48inter4));
  nand2 gate2442(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2443(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2444(.a(G8), .O(gate48inter7));
  inv1  gate2445(.a(G275), .O(gate48inter8));
  nand2 gate2446(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2447(.a(s_271), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2448(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2449(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2450(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2227(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2228(.a(gate55inter0), .b(s_240), .O(gate55inter1));
  and2  gate2229(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2230(.a(s_240), .O(gate55inter3));
  inv1  gate2231(.a(s_241), .O(gate55inter4));
  nand2 gate2232(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2233(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2234(.a(G15), .O(gate55inter7));
  inv1  gate2235(.a(G287), .O(gate55inter8));
  nand2 gate2236(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2237(.a(s_241), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2238(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2239(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2240(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate3123(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate3124(.a(gate59inter0), .b(s_368), .O(gate59inter1));
  and2  gate3125(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate3126(.a(s_368), .O(gate59inter3));
  inv1  gate3127(.a(s_369), .O(gate59inter4));
  nand2 gate3128(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate3129(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate3130(.a(G19), .O(gate59inter7));
  inv1  gate3131(.a(G293), .O(gate59inter8));
  nand2 gate3132(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate3133(.a(s_369), .b(gate59inter3), .O(gate59inter10));
  nor2  gate3134(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate3135(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate3136(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2927(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2928(.a(gate61inter0), .b(s_340), .O(gate61inter1));
  and2  gate2929(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2930(.a(s_340), .O(gate61inter3));
  inv1  gate2931(.a(s_341), .O(gate61inter4));
  nand2 gate2932(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2933(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2934(.a(G21), .O(gate61inter7));
  inv1  gate2935(.a(G296), .O(gate61inter8));
  nand2 gate2936(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2937(.a(s_341), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2938(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2939(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2940(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate603(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate604(.a(gate63inter0), .b(s_8), .O(gate63inter1));
  and2  gate605(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate606(.a(s_8), .O(gate63inter3));
  inv1  gate607(.a(s_9), .O(gate63inter4));
  nand2 gate608(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate609(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate610(.a(G23), .O(gate63inter7));
  inv1  gate611(.a(G299), .O(gate63inter8));
  nand2 gate612(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate613(.a(s_9), .b(gate63inter3), .O(gate63inter10));
  nor2  gate614(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate615(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate616(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2423(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2424(.a(gate64inter0), .b(s_268), .O(gate64inter1));
  and2  gate2425(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2426(.a(s_268), .O(gate64inter3));
  inv1  gate2427(.a(s_269), .O(gate64inter4));
  nand2 gate2428(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2429(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2430(.a(G24), .O(gate64inter7));
  inv1  gate2431(.a(G299), .O(gate64inter8));
  nand2 gate2432(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2433(.a(s_269), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2434(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2435(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2436(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate2255(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2256(.a(gate65inter0), .b(s_244), .O(gate65inter1));
  and2  gate2257(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2258(.a(s_244), .O(gate65inter3));
  inv1  gate2259(.a(s_245), .O(gate65inter4));
  nand2 gate2260(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2261(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2262(.a(G25), .O(gate65inter7));
  inv1  gate2263(.a(G302), .O(gate65inter8));
  nand2 gate2264(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2265(.a(s_245), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2266(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2267(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2268(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate645(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate646(.a(gate66inter0), .b(s_14), .O(gate66inter1));
  and2  gate647(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate648(.a(s_14), .O(gate66inter3));
  inv1  gate649(.a(s_15), .O(gate66inter4));
  nand2 gate650(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate651(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate652(.a(G26), .O(gate66inter7));
  inv1  gate653(.a(G302), .O(gate66inter8));
  nand2 gate654(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate655(.a(s_15), .b(gate66inter3), .O(gate66inter10));
  nor2  gate656(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate657(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate658(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate659(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate660(.a(gate67inter0), .b(s_16), .O(gate67inter1));
  and2  gate661(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate662(.a(s_16), .O(gate67inter3));
  inv1  gate663(.a(s_17), .O(gate67inter4));
  nand2 gate664(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate665(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate666(.a(G27), .O(gate67inter7));
  inv1  gate667(.a(G305), .O(gate67inter8));
  nand2 gate668(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate669(.a(s_17), .b(gate67inter3), .O(gate67inter10));
  nor2  gate670(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate671(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate672(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate3025(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate3026(.a(gate72inter0), .b(s_354), .O(gate72inter1));
  and2  gate3027(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate3028(.a(s_354), .O(gate72inter3));
  inv1  gate3029(.a(s_355), .O(gate72inter4));
  nand2 gate3030(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate3031(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate3032(.a(G32), .O(gate72inter7));
  inv1  gate3033(.a(G311), .O(gate72inter8));
  nand2 gate3034(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate3035(.a(s_355), .b(gate72inter3), .O(gate72inter10));
  nor2  gate3036(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate3037(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate3038(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate3039(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate3040(.a(gate73inter0), .b(s_356), .O(gate73inter1));
  and2  gate3041(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate3042(.a(s_356), .O(gate73inter3));
  inv1  gate3043(.a(s_357), .O(gate73inter4));
  nand2 gate3044(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate3045(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate3046(.a(G1), .O(gate73inter7));
  inv1  gate3047(.a(G314), .O(gate73inter8));
  nand2 gate3048(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate3049(.a(s_357), .b(gate73inter3), .O(gate73inter10));
  nor2  gate3050(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate3051(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate3052(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1163(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1164(.a(gate75inter0), .b(s_88), .O(gate75inter1));
  and2  gate1165(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1166(.a(s_88), .O(gate75inter3));
  inv1  gate1167(.a(s_89), .O(gate75inter4));
  nand2 gate1168(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1169(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1170(.a(G9), .O(gate75inter7));
  inv1  gate1171(.a(G317), .O(gate75inter8));
  nand2 gate1172(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1173(.a(s_89), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1174(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1175(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1176(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2045(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2046(.a(gate78inter0), .b(s_214), .O(gate78inter1));
  and2  gate2047(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2048(.a(s_214), .O(gate78inter3));
  inv1  gate2049(.a(s_215), .O(gate78inter4));
  nand2 gate2050(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2051(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2052(.a(G6), .O(gate78inter7));
  inv1  gate2053(.a(G320), .O(gate78inter8));
  nand2 gate2054(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2055(.a(s_215), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2056(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2057(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2058(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2479(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2480(.a(gate79inter0), .b(s_276), .O(gate79inter1));
  and2  gate2481(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2482(.a(s_276), .O(gate79inter3));
  inv1  gate2483(.a(s_277), .O(gate79inter4));
  nand2 gate2484(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2485(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2486(.a(G10), .O(gate79inter7));
  inv1  gate2487(.a(G323), .O(gate79inter8));
  nand2 gate2488(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2489(.a(s_277), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2490(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2491(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2492(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1849(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1850(.a(gate80inter0), .b(s_186), .O(gate80inter1));
  and2  gate1851(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1852(.a(s_186), .O(gate80inter3));
  inv1  gate1853(.a(s_187), .O(gate80inter4));
  nand2 gate1854(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1855(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1856(.a(G14), .O(gate80inter7));
  inv1  gate1857(.a(G323), .O(gate80inter8));
  nand2 gate1858(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1859(.a(s_187), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1860(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1861(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1862(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate3235(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate3236(.a(gate81inter0), .b(s_384), .O(gate81inter1));
  and2  gate3237(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate3238(.a(s_384), .O(gate81inter3));
  inv1  gate3239(.a(s_385), .O(gate81inter4));
  nand2 gate3240(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate3241(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate3242(.a(G3), .O(gate81inter7));
  inv1  gate3243(.a(G326), .O(gate81inter8));
  nand2 gate3244(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate3245(.a(s_385), .b(gate81inter3), .O(gate81inter10));
  nor2  gate3246(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate3247(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate3248(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1023(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1024(.a(gate82inter0), .b(s_68), .O(gate82inter1));
  and2  gate1025(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1026(.a(s_68), .O(gate82inter3));
  inv1  gate1027(.a(s_69), .O(gate82inter4));
  nand2 gate1028(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1029(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1030(.a(G7), .O(gate82inter7));
  inv1  gate1031(.a(G326), .O(gate82inter8));
  nand2 gate1032(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1033(.a(s_69), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1034(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1035(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1036(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2213(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2214(.a(gate83inter0), .b(s_238), .O(gate83inter1));
  and2  gate2215(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2216(.a(s_238), .O(gate83inter3));
  inv1  gate2217(.a(s_239), .O(gate83inter4));
  nand2 gate2218(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2219(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2220(.a(G11), .O(gate83inter7));
  inv1  gate2221(.a(G329), .O(gate83inter8));
  nand2 gate2222(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2223(.a(s_239), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2224(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2225(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2226(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate827(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate828(.a(gate86inter0), .b(s_40), .O(gate86inter1));
  and2  gate829(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate830(.a(s_40), .O(gate86inter3));
  inv1  gate831(.a(s_41), .O(gate86inter4));
  nand2 gate832(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate833(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate834(.a(G8), .O(gate86inter7));
  inv1  gate835(.a(G332), .O(gate86inter8));
  nand2 gate836(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate837(.a(s_41), .b(gate86inter3), .O(gate86inter10));
  nor2  gate838(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate839(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate840(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2101(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2102(.a(gate87inter0), .b(s_222), .O(gate87inter1));
  and2  gate2103(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2104(.a(s_222), .O(gate87inter3));
  inv1  gate2105(.a(s_223), .O(gate87inter4));
  nand2 gate2106(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2107(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2108(.a(G12), .O(gate87inter7));
  inv1  gate2109(.a(G335), .O(gate87inter8));
  nand2 gate2110(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2111(.a(s_223), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2112(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2113(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2114(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1373(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1374(.a(gate89inter0), .b(s_118), .O(gate89inter1));
  and2  gate1375(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1376(.a(s_118), .O(gate89inter3));
  inv1  gate1377(.a(s_119), .O(gate89inter4));
  nand2 gate1378(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1379(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1380(.a(G17), .O(gate89inter7));
  inv1  gate1381(.a(G338), .O(gate89inter8));
  nand2 gate1382(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1383(.a(s_119), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1384(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1385(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1386(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2605(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2606(.a(gate91inter0), .b(s_294), .O(gate91inter1));
  and2  gate2607(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2608(.a(s_294), .O(gate91inter3));
  inv1  gate2609(.a(s_295), .O(gate91inter4));
  nand2 gate2610(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2611(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2612(.a(G25), .O(gate91inter7));
  inv1  gate2613(.a(G341), .O(gate91inter8));
  nand2 gate2614(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2615(.a(s_295), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2616(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2617(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2618(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1695(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1696(.a(gate92inter0), .b(s_164), .O(gate92inter1));
  and2  gate1697(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1698(.a(s_164), .O(gate92inter3));
  inv1  gate1699(.a(s_165), .O(gate92inter4));
  nand2 gate1700(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1701(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1702(.a(G29), .O(gate92inter7));
  inv1  gate1703(.a(G341), .O(gate92inter8));
  nand2 gate1704(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1705(.a(s_165), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1706(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1707(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1708(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2171(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2172(.a(gate94inter0), .b(s_232), .O(gate94inter1));
  and2  gate2173(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2174(.a(s_232), .O(gate94inter3));
  inv1  gate2175(.a(s_233), .O(gate94inter4));
  nand2 gate2176(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2177(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2178(.a(G22), .O(gate94inter7));
  inv1  gate2179(.a(G344), .O(gate94inter8));
  nand2 gate2180(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2181(.a(s_233), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2182(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2183(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2184(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate2717(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2718(.a(gate95inter0), .b(s_310), .O(gate95inter1));
  and2  gate2719(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2720(.a(s_310), .O(gate95inter3));
  inv1  gate2721(.a(s_311), .O(gate95inter4));
  nand2 gate2722(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2723(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2724(.a(G26), .O(gate95inter7));
  inv1  gate2725(.a(G347), .O(gate95inter8));
  nand2 gate2726(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2727(.a(s_311), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2728(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2729(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2730(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1387(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1388(.a(gate97inter0), .b(s_120), .O(gate97inter1));
  and2  gate1389(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1390(.a(s_120), .O(gate97inter3));
  inv1  gate1391(.a(s_121), .O(gate97inter4));
  nand2 gate1392(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1393(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1394(.a(G19), .O(gate97inter7));
  inv1  gate1395(.a(G350), .O(gate97inter8));
  nand2 gate1396(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1397(.a(s_121), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1398(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1399(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1400(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate715(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate716(.a(gate98inter0), .b(s_24), .O(gate98inter1));
  and2  gate717(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate718(.a(s_24), .O(gate98inter3));
  inv1  gate719(.a(s_25), .O(gate98inter4));
  nand2 gate720(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate721(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate722(.a(G23), .O(gate98inter7));
  inv1  gate723(.a(G350), .O(gate98inter8));
  nand2 gate724(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate725(.a(s_25), .b(gate98inter3), .O(gate98inter10));
  nor2  gate726(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate727(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate728(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2801(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2802(.a(gate99inter0), .b(s_322), .O(gate99inter1));
  and2  gate2803(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2804(.a(s_322), .O(gate99inter3));
  inv1  gate2805(.a(s_323), .O(gate99inter4));
  nand2 gate2806(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2807(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2808(.a(G27), .O(gate99inter7));
  inv1  gate2809(.a(G353), .O(gate99inter8));
  nand2 gate2810(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2811(.a(s_323), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2812(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2813(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2814(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate3277(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate3278(.a(gate100inter0), .b(s_390), .O(gate100inter1));
  and2  gate3279(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate3280(.a(s_390), .O(gate100inter3));
  inv1  gate3281(.a(s_391), .O(gate100inter4));
  nand2 gate3282(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate3283(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate3284(.a(G31), .O(gate100inter7));
  inv1  gate3285(.a(G353), .O(gate100inter8));
  nand2 gate3286(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate3287(.a(s_391), .b(gate100inter3), .O(gate100inter10));
  nor2  gate3288(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate3289(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate3290(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate3151(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate3152(.a(gate102inter0), .b(s_372), .O(gate102inter1));
  and2  gate3153(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate3154(.a(s_372), .O(gate102inter3));
  inv1  gate3155(.a(s_373), .O(gate102inter4));
  nand2 gate3156(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate3157(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate3158(.a(G24), .O(gate102inter7));
  inv1  gate3159(.a(G356), .O(gate102inter8));
  nand2 gate3160(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate3161(.a(s_373), .b(gate102inter3), .O(gate102inter10));
  nor2  gate3162(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate3163(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate3164(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1401(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1402(.a(gate103inter0), .b(s_122), .O(gate103inter1));
  and2  gate1403(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1404(.a(s_122), .O(gate103inter3));
  inv1  gate1405(.a(s_123), .O(gate103inter4));
  nand2 gate1406(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1407(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1408(.a(G28), .O(gate103inter7));
  inv1  gate1409(.a(G359), .O(gate103inter8));
  nand2 gate1410(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1411(.a(s_123), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1412(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1413(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1414(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1541(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1542(.a(gate104inter0), .b(s_142), .O(gate104inter1));
  and2  gate1543(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1544(.a(s_142), .O(gate104inter3));
  inv1  gate1545(.a(s_143), .O(gate104inter4));
  nand2 gate1546(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1547(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1548(.a(G32), .O(gate104inter7));
  inv1  gate1549(.a(G359), .O(gate104inter8));
  nand2 gate1550(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1551(.a(s_143), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1552(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1553(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1554(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1597(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1598(.a(gate105inter0), .b(s_150), .O(gate105inter1));
  and2  gate1599(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1600(.a(s_150), .O(gate105inter3));
  inv1  gate1601(.a(s_151), .O(gate105inter4));
  nand2 gate1602(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1603(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1604(.a(G362), .O(gate105inter7));
  inv1  gate1605(.a(G363), .O(gate105inter8));
  nand2 gate1606(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1607(.a(s_151), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1608(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1609(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1610(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate561(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate562(.a(gate107inter0), .b(s_2), .O(gate107inter1));
  and2  gate563(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate564(.a(s_2), .O(gate107inter3));
  inv1  gate565(.a(s_3), .O(gate107inter4));
  nand2 gate566(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate567(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate568(.a(G366), .O(gate107inter7));
  inv1  gate569(.a(G367), .O(gate107inter8));
  nand2 gate570(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate571(.a(s_3), .b(gate107inter3), .O(gate107inter10));
  nor2  gate572(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate573(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate574(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate2703(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2704(.a(gate109inter0), .b(s_308), .O(gate109inter1));
  and2  gate2705(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2706(.a(s_308), .O(gate109inter3));
  inv1  gate2707(.a(s_309), .O(gate109inter4));
  nand2 gate2708(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2709(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2710(.a(G370), .O(gate109inter7));
  inv1  gate2711(.a(G371), .O(gate109inter8));
  nand2 gate2712(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2713(.a(s_309), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2714(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2715(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2716(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2451(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2452(.a(gate111inter0), .b(s_272), .O(gate111inter1));
  and2  gate2453(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2454(.a(s_272), .O(gate111inter3));
  inv1  gate2455(.a(s_273), .O(gate111inter4));
  nand2 gate2456(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2457(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2458(.a(G374), .O(gate111inter7));
  inv1  gate2459(.a(G375), .O(gate111inter8));
  nand2 gate2460(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2461(.a(s_273), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2462(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2463(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2464(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate589(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate590(.a(gate112inter0), .b(s_6), .O(gate112inter1));
  and2  gate591(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate592(.a(s_6), .O(gate112inter3));
  inv1  gate593(.a(s_7), .O(gate112inter4));
  nand2 gate594(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate595(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate596(.a(G376), .O(gate112inter7));
  inv1  gate597(.a(G377), .O(gate112inter8));
  nand2 gate598(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate599(.a(s_7), .b(gate112inter3), .O(gate112inter10));
  nor2  gate600(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate601(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate602(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate2465(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2466(.a(gate113inter0), .b(s_274), .O(gate113inter1));
  and2  gate2467(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2468(.a(s_274), .O(gate113inter3));
  inv1  gate2469(.a(s_275), .O(gate113inter4));
  nand2 gate2470(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2471(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2472(.a(G378), .O(gate113inter7));
  inv1  gate2473(.a(G379), .O(gate113inter8));
  nand2 gate2474(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2475(.a(s_275), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2476(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2477(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2478(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate883(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate884(.a(gate114inter0), .b(s_48), .O(gate114inter1));
  and2  gate885(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate886(.a(s_48), .O(gate114inter3));
  inv1  gate887(.a(s_49), .O(gate114inter4));
  nand2 gate888(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate889(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate890(.a(G380), .O(gate114inter7));
  inv1  gate891(.a(G381), .O(gate114inter8));
  nand2 gate892(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate893(.a(s_49), .b(gate114inter3), .O(gate114inter10));
  nor2  gate894(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate895(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate896(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate3067(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate3068(.a(gate116inter0), .b(s_360), .O(gate116inter1));
  and2  gate3069(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate3070(.a(s_360), .O(gate116inter3));
  inv1  gate3071(.a(s_361), .O(gate116inter4));
  nand2 gate3072(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate3073(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate3074(.a(G384), .O(gate116inter7));
  inv1  gate3075(.a(G385), .O(gate116inter8));
  nand2 gate3076(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate3077(.a(s_361), .b(gate116inter3), .O(gate116inter10));
  nor2  gate3078(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate3079(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate3080(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate3137(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate3138(.a(gate118inter0), .b(s_370), .O(gate118inter1));
  and2  gate3139(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate3140(.a(s_370), .O(gate118inter3));
  inv1  gate3141(.a(s_371), .O(gate118inter4));
  nand2 gate3142(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate3143(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate3144(.a(G388), .O(gate118inter7));
  inv1  gate3145(.a(G389), .O(gate118inter8));
  nand2 gate3146(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate3147(.a(s_371), .b(gate118inter3), .O(gate118inter10));
  nor2  gate3148(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate3149(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate3150(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2395(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2396(.a(gate122inter0), .b(s_264), .O(gate122inter1));
  and2  gate2397(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2398(.a(s_264), .O(gate122inter3));
  inv1  gate2399(.a(s_265), .O(gate122inter4));
  nand2 gate2400(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2401(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2402(.a(G396), .O(gate122inter7));
  inv1  gate2403(.a(G397), .O(gate122inter8));
  nand2 gate2404(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2405(.a(s_265), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2406(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2407(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2408(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate673(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate674(.a(gate123inter0), .b(s_18), .O(gate123inter1));
  and2  gate675(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate676(.a(s_18), .O(gate123inter3));
  inv1  gate677(.a(s_19), .O(gate123inter4));
  nand2 gate678(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate679(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate680(.a(G398), .O(gate123inter7));
  inv1  gate681(.a(G399), .O(gate123inter8));
  nand2 gate682(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate683(.a(s_19), .b(gate123inter3), .O(gate123inter10));
  nor2  gate684(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate685(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate686(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate869(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate870(.a(gate128inter0), .b(s_46), .O(gate128inter1));
  and2  gate871(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate872(.a(s_46), .O(gate128inter3));
  inv1  gate873(.a(s_47), .O(gate128inter4));
  nand2 gate874(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate875(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate876(.a(G408), .O(gate128inter7));
  inv1  gate877(.a(G409), .O(gate128inter8));
  nand2 gate878(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate879(.a(s_47), .b(gate128inter3), .O(gate128inter10));
  nor2  gate880(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate881(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate882(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate2409(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2410(.a(gate129inter0), .b(s_266), .O(gate129inter1));
  and2  gate2411(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2412(.a(s_266), .O(gate129inter3));
  inv1  gate2413(.a(s_267), .O(gate129inter4));
  nand2 gate2414(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2415(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2416(.a(G410), .O(gate129inter7));
  inv1  gate2417(.a(G411), .O(gate129inter8));
  nand2 gate2418(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2419(.a(s_267), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2420(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2421(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2422(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1653(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1654(.a(gate132inter0), .b(s_158), .O(gate132inter1));
  and2  gate1655(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1656(.a(s_158), .O(gate132inter3));
  inv1  gate1657(.a(s_159), .O(gate132inter4));
  nand2 gate1658(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1659(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1660(.a(G416), .O(gate132inter7));
  inv1  gate1661(.a(G417), .O(gate132inter8));
  nand2 gate1662(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1663(.a(s_159), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1664(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1665(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1666(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1667(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1668(.a(gate133inter0), .b(s_160), .O(gate133inter1));
  and2  gate1669(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1670(.a(s_160), .O(gate133inter3));
  inv1  gate1671(.a(s_161), .O(gate133inter4));
  nand2 gate1672(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1673(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1674(.a(G418), .O(gate133inter7));
  inv1  gate1675(.a(G419), .O(gate133inter8));
  nand2 gate1676(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1677(.a(s_161), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1678(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1679(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1680(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1751(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1752(.a(gate134inter0), .b(s_172), .O(gate134inter1));
  and2  gate1753(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1754(.a(s_172), .O(gate134inter3));
  inv1  gate1755(.a(s_173), .O(gate134inter4));
  nand2 gate1756(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1757(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1758(.a(G420), .O(gate134inter7));
  inv1  gate1759(.a(G421), .O(gate134inter8));
  nand2 gate1760(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1761(.a(s_173), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1762(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1763(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1764(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2367(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2368(.a(gate138inter0), .b(s_260), .O(gate138inter1));
  and2  gate2369(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2370(.a(s_260), .O(gate138inter3));
  inv1  gate2371(.a(s_261), .O(gate138inter4));
  nand2 gate2372(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2373(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2374(.a(G432), .O(gate138inter7));
  inv1  gate2375(.a(G435), .O(gate138inter8));
  nand2 gate2376(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2377(.a(s_261), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2378(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2379(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2380(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2941(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2942(.a(gate142inter0), .b(s_342), .O(gate142inter1));
  and2  gate2943(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2944(.a(s_342), .O(gate142inter3));
  inv1  gate2945(.a(s_343), .O(gate142inter4));
  nand2 gate2946(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2947(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2948(.a(G456), .O(gate142inter7));
  inv1  gate2949(.a(G459), .O(gate142inter8));
  nand2 gate2950(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2951(.a(s_343), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2952(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2953(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2954(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2059(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2060(.a(gate153inter0), .b(s_216), .O(gate153inter1));
  and2  gate2061(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2062(.a(s_216), .O(gate153inter3));
  inv1  gate2063(.a(s_217), .O(gate153inter4));
  nand2 gate2064(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2065(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2066(.a(G426), .O(gate153inter7));
  inv1  gate2067(.a(G522), .O(gate153inter8));
  nand2 gate2068(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2069(.a(s_217), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2070(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2071(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2072(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1191(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1192(.a(gate155inter0), .b(s_92), .O(gate155inter1));
  and2  gate1193(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1194(.a(s_92), .O(gate155inter3));
  inv1  gate1195(.a(s_93), .O(gate155inter4));
  nand2 gate1196(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1197(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1198(.a(G432), .O(gate155inter7));
  inv1  gate1199(.a(G525), .O(gate155inter8));
  nand2 gate1200(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1201(.a(s_93), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1202(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1203(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1204(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate3053(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate3054(.a(gate156inter0), .b(s_358), .O(gate156inter1));
  and2  gate3055(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate3056(.a(s_358), .O(gate156inter3));
  inv1  gate3057(.a(s_359), .O(gate156inter4));
  nand2 gate3058(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate3059(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate3060(.a(G435), .O(gate156inter7));
  inv1  gate3061(.a(G525), .O(gate156inter8));
  nand2 gate3062(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate3063(.a(s_359), .b(gate156inter3), .O(gate156inter10));
  nor2  gate3064(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate3065(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate3066(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1723(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1724(.a(gate165inter0), .b(s_168), .O(gate165inter1));
  and2  gate1725(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1726(.a(s_168), .O(gate165inter3));
  inv1  gate1727(.a(s_169), .O(gate165inter4));
  nand2 gate1728(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1729(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1730(.a(G462), .O(gate165inter7));
  inv1  gate1731(.a(G540), .O(gate165inter8));
  nand2 gate1732(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1733(.a(s_169), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1734(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1735(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1736(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1107(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1108(.a(gate166inter0), .b(s_80), .O(gate166inter1));
  and2  gate1109(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1110(.a(s_80), .O(gate166inter3));
  inv1  gate1111(.a(s_81), .O(gate166inter4));
  nand2 gate1112(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1113(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1114(.a(G465), .O(gate166inter7));
  inv1  gate1115(.a(G540), .O(gate166inter8));
  nand2 gate1116(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1117(.a(s_81), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1118(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1119(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1120(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2507(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2508(.a(gate167inter0), .b(s_280), .O(gate167inter1));
  and2  gate2509(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2510(.a(s_280), .O(gate167inter3));
  inv1  gate2511(.a(s_281), .O(gate167inter4));
  nand2 gate2512(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2513(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2514(.a(G468), .O(gate167inter7));
  inv1  gate2515(.a(G543), .O(gate167inter8));
  nand2 gate2516(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2517(.a(s_281), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2518(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2519(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2520(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate841(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate842(.a(gate168inter0), .b(s_42), .O(gate168inter1));
  and2  gate843(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate844(.a(s_42), .O(gate168inter3));
  inv1  gate845(.a(s_43), .O(gate168inter4));
  nand2 gate846(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate847(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate848(.a(G471), .O(gate168inter7));
  inv1  gate849(.a(G543), .O(gate168inter8));
  nand2 gate850(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate851(.a(s_43), .b(gate168inter3), .O(gate168inter10));
  nor2  gate852(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate853(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate854(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1555(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1556(.a(gate169inter0), .b(s_144), .O(gate169inter1));
  and2  gate1557(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1558(.a(s_144), .O(gate169inter3));
  inv1  gate1559(.a(s_145), .O(gate169inter4));
  nand2 gate1560(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1561(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1562(.a(G474), .O(gate169inter7));
  inv1  gate1563(.a(G546), .O(gate169inter8));
  nand2 gate1564(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1565(.a(s_145), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1566(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1567(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1568(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1513(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1514(.a(gate172inter0), .b(s_138), .O(gate172inter1));
  and2  gate1515(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1516(.a(s_138), .O(gate172inter3));
  inv1  gate1517(.a(s_139), .O(gate172inter4));
  nand2 gate1518(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1519(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1520(.a(G483), .O(gate172inter7));
  inv1  gate1521(.a(G549), .O(gate172inter8));
  nand2 gate1522(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1523(.a(s_139), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1524(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1525(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1526(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate3263(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate3264(.a(gate174inter0), .b(s_388), .O(gate174inter1));
  and2  gate3265(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate3266(.a(s_388), .O(gate174inter3));
  inv1  gate3267(.a(s_389), .O(gate174inter4));
  nand2 gate3268(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate3269(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate3270(.a(G489), .O(gate174inter7));
  inv1  gate3271(.a(G552), .O(gate174inter8));
  nand2 gate3272(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate3273(.a(s_389), .b(gate174inter3), .O(gate174inter10));
  nor2  gate3274(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate3275(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate3276(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2115(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2116(.a(gate176inter0), .b(s_224), .O(gate176inter1));
  and2  gate2117(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2118(.a(s_224), .O(gate176inter3));
  inv1  gate2119(.a(s_225), .O(gate176inter4));
  nand2 gate2120(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2121(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2122(.a(G495), .O(gate176inter7));
  inv1  gate2123(.a(G555), .O(gate176inter8));
  nand2 gate2124(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2125(.a(s_225), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2126(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2127(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2128(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate3249(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate3250(.a(gate180inter0), .b(s_386), .O(gate180inter1));
  and2  gate3251(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate3252(.a(s_386), .O(gate180inter3));
  inv1  gate3253(.a(s_387), .O(gate180inter4));
  nand2 gate3254(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate3255(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate3256(.a(G507), .O(gate180inter7));
  inv1  gate3257(.a(G561), .O(gate180inter8));
  nand2 gate3258(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate3259(.a(s_387), .b(gate180inter3), .O(gate180inter10));
  nor2  gate3260(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate3261(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate3262(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate995(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate996(.a(gate181inter0), .b(s_64), .O(gate181inter1));
  and2  gate997(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate998(.a(s_64), .O(gate181inter3));
  inv1  gate999(.a(s_65), .O(gate181inter4));
  nand2 gate1000(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1001(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1002(.a(G510), .O(gate181inter7));
  inv1  gate1003(.a(G564), .O(gate181inter8));
  nand2 gate1004(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1005(.a(s_65), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1006(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1007(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1008(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate911(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate912(.a(gate184inter0), .b(s_52), .O(gate184inter1));
  and2  gate913(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate914(.a(s_52), .O(gate184inter3));
  inv1  gate915(.a(s_53), .O(gate184inter4));
  nand2 gate916(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate917(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate918(.a(G519), .O(gate184inter7));
  inv1  gate919(.a(G567), .O(gate184inter8));
  nand2 gate920(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate921(.a(s_53), .b(gate184inter3), .O(gate184inter10));
  nor2  gate922(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate923(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate924(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2759(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2760(.a(gate188inter0), .b(s_316), .O(gate188inter1));
  and2  gate2761(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2762(.a(s_316), .O(gate188inter3));
  inv1  gate2763(.a(s_317), .O(gate188inter4));
  nand2 gate2764(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2765(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2766(.a(G576), .O(gate188inter7));
  inv1  gate2767(.a(G577), .O(gate188inter8));
  nand2 gate2768(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2769(.a(s_317), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2770(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2771(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2772(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2913(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2914(.a(gate190inter0), .b(s_338), .O(gate190inter1));
  and2  gate2915(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2916(.a(s_338), .O(gate190inter3));
  inv1  gate2917(.a(s_339), .O(gate190inter4));
  nand2 gate2918(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2919(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2920(.a(G580), .O(gate190inter7));
  inv1  gate2921(.a(G581), .O(gate190inter8));
  nand2 gate2922(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2923(.a(s_339), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2924(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2925(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2926(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate3207(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate3208(.a(gate191inter0), .b(s_380), .O(gate191inter1));
  and2  gate3209(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate3210(.a(s_380), .O(gate191inter3));
  inv1  gate3211(.a(s_381), .O(gate191inter4));
  nand2 gate3212(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate3213(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate3214(.a(G582), .O(gate191inter7));
  inv1  gate3215(.a(G583), .O(gate191inter8));
  nand2 gate3216(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate3217(.a(s_381), .b(gate191inter3), .O(gate191inter10));
  nor2  gate3218(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate3219(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate3220(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1485(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1486(.a(gate192inter0), .b(s_134), .O(gate192inter1));
  and2  gate1487(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1488(.a(s_134), .O(gate192inter3));
  inv1  gate1489(.a(s_135), .O(gate192inter4));
  nand2 gate1490(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1491(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1492(.a(G584), .O(gate192inter7));
  inv1  gate1493(.a(G585), .O(gate192inter8));
  nand2 gate1494(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1495(.a(s_135), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1496(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1497(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1498(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1877(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1878(.a(gate196inter0), .b(s_190), .O(gate196inter1));
  and2  gate1879(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1880(.a(s_190), .O(gate196inter3));
  inv1  gate1881(.a(s_191), .O(gate196inter4));
  nand2 gate1882(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1883(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1884(.a(G592), .O(gate196inter7));
  inv1  gate1885(.a(G593), .O(gate196inter8));
  nand2 gate1886(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1887(.a(s_191), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1888(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1889(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1890(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate3179(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate3180(.a(gate197inter0), .b(s_376), .O(gate197inter1));
  and2  gate3181(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate3182(.a(s_376), .O(gate197inter3));
  inv1  gate3183(.a(s_377), .O(gate197inter4));
  nand2 gate3184(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate3185(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate3186(.a(G594), .O(gate197inter7));
  inv1  gate3187(.a(G595), .O(gate197inter8));
  nand2 gate3188(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate3189(.a(s_377), .b(gate197inter3), .O(gate197inter10));
  nor2  gate3190(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate3191(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate3192(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1149(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1150(.a(gate199inter0), .b(s_86), .O(gate199inter1));
  and2  gate1151(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1152(.a(s_86), .O(gate199inter3));
  inv1  gate1153(.a(s_87), .O(gate199inter4));
  nand2 gate1154(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1155(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1156(.a(G598), .O(gate199inter7));
  inv1  gate1157(.a(G599), .O(gate199inter8));
  nand2 gate1158(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1159(.a(s_87), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1160(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1161(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1162(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2563(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2564(.a(gate201inter0), .b(s_288), .O(gate201inter1));
  and2  gate2565(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2566(.a(s_288), .O(gate201inter3));
  inv1  gate2567(.a(s_289), .O(gate201inter4));
  nand2 gate2568(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2569(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2570(.a(G602), .O(gate201inter7));
  inv1  gate2571(.a(G607), .O(gate201inter8));
  nand2 gate2572(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2573(.a(s_289), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2574(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2575(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2576(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1737(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1738(.a(gate202inter0), .b(s_170), .O(gate202inter1));
  and2  gate1739(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1740(.a(s_170), .O(gate202inter3));
  inv1  gate1741(.a(s_171), .O(gate202inter4));
  nand2 gate1742(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1743(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1744(.a(G612), .O(gate202inter7));
  inv1  gate1745(.a(G617), .O(gate202inter8));
  nand2 gate1746(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1747(.a(s_171), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1748(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1749(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1750(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2983(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2984(.a(gate204inter0), .b(s_348), .O(gate204inter1));
  and2  gate2985(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2986(.a(s_348), .O(gate204inter3));
  inv1  gate2987(.a(s_349), .O(gate204inter4));
  nand2 gate2988(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2989(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2990(.a(G607), .O(gate204inter7));
  inv1  gate2991(.a(G617), .O(gate204inter8));
  nand2 gate2992(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2993(.a(s_349), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2994(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2995(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2996(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate617(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate618(.a(gate206inter0), .b(s_10), .O(gate206inter1));
  and2  gate619(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate620(.a(s_10), .O(gate206inter3));
  inv1  gate621(.a(s_11), .O(gate206inter4));
  nand2 gate622(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate623(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate624(.a(G632), .O(gate206inter7));
  inv1  gate625(.a(G637), .O(gate206inter8));
  nand2 gate626(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate627(.a(s_11), .b(gate206inter3), .O(gate206inter10));
  nor2  gate628(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate629(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate630(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2353(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2354(.a(gate210inter0), .b(s_258), .O(gate210inter1));
  and2  gate2355(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2356(.a(s_258), .O(gate210inter3));
  inv1  gate2357(.a(s_259), .O(gate210inter4));
  nand2 gate2358(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2359(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2360(.a(G607), .O(gate210inter7));
  inv1  gate2361(.a(G666), .O(gate210inter8));
  nand2 gate2362(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2363(.a(s_259), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2364(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2365(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2366(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1121(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1122(.a(gate211inter0), .b(s_82), .O(gate211inter1));
  and2  gate1123(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1124(.a(s_82), .O(gate211inter3));
  inv1  gate1125(.a(s_83), .O(gate211inter4));
  nand2 gate1126(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1127(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1128(.a(G612), .O(gate211inter7));
  inv1  gate1129(.a(G669), .O(gate211inter8));
  nand2 gate1130(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1131(.a(s_83), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1132(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1133(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1134(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate981(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate982(.a(gate213inter0), .b(s_62), .O(gate213inter1));
  and2  gate983(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate984(.a(s_62), .O(gate213inter3));
  inv1  gate985(.a(s_63), .O(gate213inter4));
  nand2 gate986(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate987(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate988(.a(G602), .O(gate213inter7));
  inv1  gate989(.a(G672), .O(gate213inter8));
  nand2 gate990(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate991(.a(s_63), .b(gate213inter3), .O(gate213inter10));
  nor2  gate992(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate993(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate994(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate575(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate576(.a(gate218inter0), .b(s_4), .O(gate218inter1));
  and2  gate577(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate578(.a(s_4), .O(gate218inter3));
  inv1  gate579(.a(s_5), .O(gate218inter4));
  nand2 gate580(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate581(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate582(.a(G627), .O(gate218inter7));
  inv1  gate583(.a(G678), .O(gate218inter8));
  nand2 gate584(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate585(.a(s_5), .b(gate218inter3), .O(gate218inter10));
  nor2  gate586(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate587(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate588(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate3165(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate3166(.a(gate220inter0), .b(s_374), .O(gate220inter1));
  and2  gate3167(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate3168(.a(s_374), .O(gate220inter3));
  inv1  gate3169(.a(s_375), .O(gate220inter4));
  nand2 gate3170(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate3171(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate3172(.a(G637), .O(gate220inter7));
  inv1  gate3173(.a(G681), .O(gate220inter8));
  nand2 gate3174(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate3175(.a(s_375), .b(gate220inter3), .O(gate220inter10));
  nor2  gate3176(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate3177(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate3178(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate3095(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate3096(.a(gate222inter0), .b(s_364), .O(gate222inter1));
  and2  gate3097(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate3098(.a(s_364), .O(gate222inter3));
  inv1  gate3099(.a(s_365), .O(gate222inter4));
  nand2 gate3100(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate3101(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate3102(.a(G632), .O(gate222inter7));
  inv1  gate3103(.a(G684), .O(gate222inter8));
  nand2 gate3104(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate3105(.a(s_365), .b(gate222inter3), .O(gate222inter10));
  nor2  gate3106(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate3107(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate3108(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate771(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate772(.a(gate226inter0), .b(s_32), .O(gate226inter1));
  and2  gate773(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate774(.a(s_32), .O(gate226inter3));
  inv1  gate775(.a(s_33), .O(gate226inter4));
  nand2 gate776(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate777(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate778(.a(G692), .O(gate226inter7));
  inv1  gate779(.a(G693), .O(gate226inter8));
  nand2 gate780(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate781(.a(s_33), .b(gate226inter3), .O(gate226inter10));
  nor2  gate782(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate783(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate784(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1863(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1864(.a(gate227inter0), .b(s_188), .O(gate227inter1));
  and2  gate1865(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1866(.a(s_188), .O(gate227inter3));
  inv1  gate1867(.a(s_189), .O(gate227inter4));
  nand2 gate1868(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1869(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1870(.a(G694), .O(gate227inter7));
  inv1  gate1871(.a(G695), .O(gate227inter8));
  nand2 gate1872(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1873(.a(s_189), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1874(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1875(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1876(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1415(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1416(.a(gate228inter0), .b(s_124), .O(gate228inter1));
  and2  gate1417(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1418(.a(s_124), .O(gate228inter3));
  inv1  gate1419(.a(s_125), .O(gate228inter4));
  nand2 gate1420(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1421(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1422(.a(G696), .O(gate228inter7));
  inv1  gate1423(.a(G697), .O(gate228inter8));
  nand2 gate1424(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1425(.a(s_125), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1426(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1427(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1428(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate757(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate758(.a(gate229inter0), .b(s_30), .O(gate229inter1));
  and2  gate759(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate760(.a(s_30), .O(gate229inter3));
  inv1  gate761(.a(s_31), .O(gate229inter4));
  nand2 gate762(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate763(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate764(.a(G698), .O(gate229inter7));
  inv1  gate765(.a(G699), .O(gate229inter8));
  nand2 gate766(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate767(.a(s_31), .b(gate229inter3), .O(gate229inter10));
  nor2  gate768(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate769(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate770(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate855(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate856(.a(gate230inter0), .b(s_44), .O(gate230inter1));
  and2  gate857(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate858(.a(s_44), .O(gate230inter3));
  inv1  gate859(.a(s_45), .O(gate230inter4));
  nand2 gate860(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate861(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate862(.a(G700), .O(gate230inter7));
  inv1  gate863(.a(G701), .O(gate230inter8));
  nand2 gate864(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate865(.a(s_45), .b(gate230inter3), .O(gate230inter10));
  nor2  gate866(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate867(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate868(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2689(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2690(.a(gate232inter0), .b(s_306), .O(gate232inter1));
  and2  gate2691(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2692(.a(s_306), .O(gate232inter3));
  inv1  gate2693(.a(s_307), .O(gate232inter4));
  nand2 gate2694(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2695(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2696(.a(G704), .O(gate232inter7));
  inv1  gate2697(.a(G705), .O(gate232inter8));
  nand2 gate2698(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2699(.a(s_307), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2700(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2701(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2702(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2325(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2326(.a(gate234inter0), .b(s_254), .O(gate234inter1));
  and2  gate2327(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2328(.a(s_254), .O(gate234inter3));
  inv1  gate2329(.a(s_255), .O(gate234inter4));
  nand2 gate2330(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2331(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2332(.a(G245), .O(gate234inter7));
  inv1  gate2333(.a(G721), .O(gate234inter8));
  nand2 gate2334(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2335(.a(s_255), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2336(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2337(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2338(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate799(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate800(.a(gate235inter0), .b(s_36), .O(gate235inter1));
  and2  gate801(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate802(.a(s_36), .O(gate235inter3));
  inv1  gate803(.a(s_37), .O(gate235inter4));
  nand2 gate804(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate805(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate806(.a(G248), .O(gate235inter7));
  inv1  gate807(.a(G724), .O(gate235inter8));
  nand2 gate808(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate809(.a(s_37), .b(gate235inter3), .O(gate235inter10));
  nor2  gate810(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate811(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate812(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate729(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate730(.a(gate238inter0), .b(s_26), .O(gate238inter1));
  and2  gate731(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate732(.a(s_26), .O(gate238inter3));
  inv1  gate733(.a(s_27), .O(gate238inter4));
  nand2 gate734(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate735(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate736(.a(G257), .O(gate238inter7));
  inv1  gate737(.a(G709), .O(gate238inter8));
  nand2 gate738(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate739(.a(s_27), .b(gate238inter3), .O(gate238inter10));
  nor2  gate740(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate741(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate742(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1471(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1472(.a(gate239inter0), .b(s_132), .O(gate239inter1));
  and2  gate1473(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1474(.a(s_132), .O(gate239inter3));
  inv1  gate1475(.a(s_133), .O(gate239inter4));
  nand2 gate1476(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1477(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1478(.a(G260), .O(gate239inter7));
  inv1  gate1479(.a(G712), .O(gate239inter8));
  nand2 gate1480(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1481(.a(s_133), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1482(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1483(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1484(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2241(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2242(.a(gate243inter0), .b(s_242), .O(gate243inter1));
  and2  gate2243(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2244(.a(s_242), .O(gate243inter3));
  inv1  gate2245(.a(s_243), .O(gate243inter4));
  nand2 gate2246(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2247(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2248(.a(G245), .O(gate243inter7));
  inv1  gate2249(.a(G733), .O(gate243inter8));
  nand2 gate2250(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2251(.a(s_243), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2252(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2253(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2254(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate925(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate926(.a(gate245inter0), .b(s_54), .O(gate245inter1));
  and2  gate927(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate928(.a(s_54), .O(gate245inter3));
  inv1  gate929(.a(s_55), .O(gate245inter4));
  nand2 gate930(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate931(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate932(.a(G248), .O(gate245inter7));
  inv1  gate933(.a(G736), .O(gate245inter8));
  nand2 gate934(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate935(.a(s_55), .b(gate245inter3), .O(gate245inter10));
  nor2  gate936(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate937(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate938(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2731(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2732(.a(gate249inter0), .b(s_312), .O(gate249inter1));
  and2  gate2733(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2734(.a(s_312), .O(gate249inter3));
  inv1  gate2735(.a(s_313), .O(gate249inter4));
  nand2 gate2736(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2737(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2738(.a(G254), .O(gate249inter7));
  inv1  gate2739(.a(G742), .O(gate249inter8));
  nand2 gate2740(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2741(.a(s_313), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2742(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2743(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2744(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2087(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2088(.a(gate250inter0), .b(s_220), .O(gate250inter1));
  and2  gate2089(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2090(.a(s_220), .O(gate250inter3));
  inv1  gate2091(.a(s_221), .O(gate250inter4));
  nand2 gate2092(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2093(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2094(.a(G706), .O(gate250inter7));
  inv1  gate2095(.a(G742), .O(gate250inter8));
  nand2 gate2096(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2097(.a(s_221), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2098(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2099(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2100(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2829(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2830(.a(gate251inter0), .b(s_326), .O(gate251inter1));
  and2  gate2831(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2832(.a(s_326), .O(gate251inter3));
  inv1  gate2833(.a(s_327), .O(gate251inter4));
  nand2 gate2834(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2835(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2836(.a(G257), .O(gate251inter7));
  inv1  gate2837(.a(G745), .O(gate251inter8));
  nand2 gate2838(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2839(.a(s_327), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2840(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2841(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2842(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1989(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1990(.a(gate252inter0), .b(s_206), .O(gate252inter1));
  and2  gate1991(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1992(.a(s_206), .O(gate252inter3));
  inv1  gate1993(.a(s_207), .O(gate252inter4));
  nand2 gate1994(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1995(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1996(.a(G709), .O(gate252inter7));
  inv1  gate1997(.a(G745), .O(gate252inter8));
  nand2 gate1998(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1999(.a(s_207), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2000(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2001(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2002(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate1429(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1430(.a(gate253inter0), .b(s_126), .O(gate253inter1));
  and2  gate1431(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1432(.a(s_126), .O(gate253inter3));
  inv1  gate1433(.a(s_127), .O(gate253inter4));
  nand2 gate1434(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1435(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1436(.a(G260), .O(gate253inter7));
  inv1  gate1437(.a(G748), .O(gate253inter8));
  nand2 gate1438(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1439(.a(s_127), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1440(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1441(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1442(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2577(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2578(.a(gate256inter0), .b(s_290), .O(gate256inter1));
  and2  gate2579(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2580(.a(s_290), .O(gate256inter3));
  inv1  gate2581(.a(s_291), .O(gate256inter4));
  nand2 gate2582(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2583(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2584(.a(G715), .O(gate256inter7));
  inv1  gate2585(.a(G751), .O(gate256inter8));
  nand2 gate2586(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2587(.a(s_291), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2588(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2589(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2590(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate2773(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2774(.a(gate259inter0), .b(s_318), .O(gate259inter1));
  and2  gate2775(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2776(.a(s_318), .O(gate259inter3));
  inv1  gate2777(.a(s_319), .O(gate259inter4));
  nand2 gate2778(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2779(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2780(.a(G758), .O(gate259inter7));
  inv1  gate2781(.a(G759), .O(gate259inter8));
  nand2 gate2782(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2783(.a(s_319), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2784(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2785(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2786(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2815(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2816(.a(gate262inter0), .b(s_324), .O(gate262inter1));
  and2  gate2817(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2818(.a(s_324), .O(gate262inter3));
  inv1  gate2819(.a(s_325), .O(gate262inter4));
  nand2 gate2820(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2821(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2822(.a(G764), .O(gate262inter7));
  inv1  gate2823(.a(G765), .O(gate262inter8));
  nand2 gate2824(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2825(.a(s_325), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2826(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2827(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2828(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2311(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2312(.a(gate263inter0), .b(s_252), .O(gate263inter1));
  and2  gate2313(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2314(.a(s_252), .O(gate263inter3));
  inv1  gate2315(.a(s_253), .O(gate263inter4));
  nand2 gate2316(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2317(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2318(.a(G766), .O(gate263inter7));
  inv1  gate2319(.a(G767), .O(gate263inter8));
  nand2 gate2320(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2321(.a(s_253), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2322(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2323(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2324(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1009(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1010(.a(gate266inter0), .b(s_66), .O(gate266inter1));
  and2  gate1011(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1012(.a(s_66), .O(gate266inter3));
  inv1  gate1013(.a(s_67), .O(gate266inter4));
  nand2 gate1014(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1015(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1016(.a(G645), .O(gate266inter7));
  inv1  gate1017(.a(G773), .O(gate266inter8));
  nand2 gate1018(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1019(.a(s_67), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1020(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1021(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1022(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2521(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2522(.a(gate267inter0), .b(s_282), .O(gate267inter1));
  and2  gate2523(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2524(.a(s_282), .O(gate267inter3));
  inv1  gate2525(.a(s_283), .O(gate267inter4));
  nand2 gate2526(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2527(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2528(.a(G648), .O(gate267inter7));
  inv1  gate2529(.a(G776), .O(gate267inter8));
  nand2 gate2530(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2531(.a(s_283), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2532(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2533(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2534(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2843(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2844(.a(gate269inter0), .b(s_328), .O(gate269inter1));
  and2  gate2845(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2846(.a(s_328), .O(gate269inter3));
  inv1  gate2847(.a(s_329), .O(gate269inter4));
  nand2 gate2848(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2849(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2850(.a(G654), .O(gate269inter7));
  inv1  gate2851(.a(G782), .O(gate269inter8));
  nand2 gate2852(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2853(.a(s_329), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2854(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2855(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2856(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1835(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1836(.a(gate271inter0), .b(s_184), .O(gate271inter1));
  and2  gate1837(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1838(.a(s_184), .O(gate271inter3));
  inv1  gate1839(.a(s_185), .O(gate271inter4));
  nand2 gate1840(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1841(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1842(.a(G660), .O(gate271inter7));
  inv1  gate1843(.a(G788), .O(gate271inter8));
  nand2 gate1844(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1845(.a(s_185), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1846(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1847(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1848(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1793(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1794(.a(gate274inter0), .b(s_178), .O(gate274inter1));
  and2  gate1795(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1796(.a(s_178), .O(gate274inter3));
  inv1  gate1797(.a(s_179), .O(gate274inter4));
  nand2 gate1798(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1799(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1800(.a(G770), .O(gate274inter7));
  inv1  gate1801(.a(G794), .O(gate274inter8));
  nand2 gate1802(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1803(.a(s_179), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1804(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1805(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1806(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1177(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1178(.a(gate275inter0), .b(s_90), .O(gate275inter1));
  and2  gate1179(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1180(.a(s_90), .O(gate275inter3));
  inv1  gate1181(.a(s_91), .O(gate275inter4));
  nand2 gate1182(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1183(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1184(.a(G645), .O(gate275inter7));
  inv1  gate1185(.a(G797), .O(gate275inter8));
  nand2 gate1186(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1187(.a(s_91), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1188(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1189(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1190(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2269(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2270(.a(gate277inter0), .b(s_246), .O(gate277inter1));
  and2  gate2271(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2272(.a(s_246), .O(gate277inter3));
  inv1  gate2273(.a(s_247), .O(gate277inter4));
  nand2 gate2274(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2275(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2276(.a(G648), .O(gate277inter7));
  inv1  gate2277(.a(G800), .O(gate277inter8));
  nand2 gate2278(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2279(.a(s_247), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2280(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2281(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2282(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1807(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1808(.a(gate279inter0), .b(s_180), .O(gate279inter1));
  and2  gate1809(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1810(.a(s_180), .O(gate279inter3));
  inv1  gate1811(.a(s_181), .O(gate279inter4));
  nand2 gate1812(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1813(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1814(.a(G651), .O(gate279inter7));
  inv1  gate1815(.a(G803), .O(gate279inter8));
  nand2 gate1816(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1817(.a(s_181), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1818(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1819(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1820(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1975(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1976(.a(gate280inter0), .b(s_204), .O(gate280inter1));
  and2  gate1977(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1978(.a(s_204), .O(gate280inter3));
  inv1  gate1979(.a(s_205), .O(gate280inter4));
  nand2 gate1980(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1981(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1982(.a(G779), .O(gate280inter7));
  inv1  gate1983(.a(G803), .O(gate280inter8));
  nand2 gate1984(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1985(.a(s_205), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1986(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1987(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1988(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1499(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1500(.a(gate284inter0), .b(s_136), .O(gate284inter1));
  and2  gate1501(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1502(.a(s_136), .O(gate284inter3));
  inv1  gate1503(.a(s_137), .O(gate284inter4));
  nand2 gate1504(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1505(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1506(.a(G785), .O(gate284inter7));
  inv1  gate1507(.a(G809), .O(gate284inter8));
  nand2 gate1508(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1509(.a(s_137), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1510(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1511(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1512(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1275(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1276(.a(gate285inter0), .b(s_104), .O(gate285inter1));
  and2  gate1277(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1278(.a(s_104), .O(gate285inter3));
  inv1  gate1279(.a(s_105), .O(gate285inter4));
  nand2 gate1280(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1281(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1282(.a(G660), .O(gate285inter7));
  inv1  gate1283(.a(G812), .O(gate285inter8));
  nand2 gate1284(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1285(.a(s_105), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1286(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1287(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1288(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2185(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2186(.a(gate286inter0), .b(s_234), .O(gate286inter1));
  and2  gate2187(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2188(.a(s_234), .O(gate286inter3));
  inv1  gate2189(.a(s_235), .O(gate286inter4));
  nand2 gate2190(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2191(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2192(.a(G788), .O(gate286inter7));
  inv1  gate2193(.a(G812), .O(gate286inter8));
  nand2 gate2194(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2195(.a(s_235), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2196(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2197(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2198(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2339(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2340(.a(gate287inter0), .b(s_256), .O(gate287inter1));
  and2  gate2341(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2342(.a(s_256), .O(gate287inter3));
  inv1  gate2343(.a(s_257), .O(gate287inter4));
  nand2 gate2344(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2345(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2346(.a(G663), .O(gate287inter7));
  inv1  gate2347(.a(G815), .O(gate287inter8));
  nand2 gate2348(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2349(.a(s_257), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2350(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2351(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2352(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2857(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2858(.a(gate289inter0), .b(s_330), .O(gate289inter1));
  and2  gate2859(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2860(.a(s_330), .O(gate289inter3));
  inv1  gate2861(.a(s_331), .O(gate289inter4));
  nand2 gate2862(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2863(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2864(.a(G818), .O(gate289inter7));
  inv1  gate2865(.a(G819), .O(gate289inter8));
  nand2 gate2866(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2867(.a(s_331), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2868(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2869(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2870(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate3081(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate3082(.a(gate290inter0), .b(s_362), .O(gate290inter1));
  and2  gate3083(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate3084(.a(s_362), .O(gate290inter3));
  inv1  gate3085(.a(s_363), .O(gate290inter4));
  nand2 gate3086(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate3087(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate3088(.a(G820), .O(gate290inter7));
  inv1  gate3089(.a(G821), .O(gate290inter8));
  nand2 gate3090(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate3091(.a(s_363), .b(gate290inter3), .O(gate290inter10));
  nor2  gate3092(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate3093(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate3094(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1625(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1626(.a(gate291inter0), .b(s_154), .O(gate291inter1));
  and2  gate1627(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1628(.a(s_154), .O(gate291inter3));
  inv1  gate1629(.a(s_155), .O(gate291inter4));
  nand2 gate1630(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1631(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1632(.a(G822), .O(gate291inter7));
  inv1  gate1633(.a(G823), .O(gate291inter8));
  nand2 gate1634(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1635(.a(s_155), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1636(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1637(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1638(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate3109(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate3110(.a(gate294inter0), .b(s_366), .O(gate294inter1));
  and2  gate3111(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate3112(.a(s_366), .O(gate294inter3));
  inv1  gate3113(.a(s_367), .O(gate294inter4));
  nand2 gate3114(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate3115(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate3116(.a(G832), .O(gate294inter7));
  inv1  gate3117(.a(G833), .O(gate294inter8));
  nand2 gate3118(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate3119(.a(s_367), .b(gate294inter3), .O(gate294inter10));
  nor2  gate3120(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate3121(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate3122(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2633(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2634(.a(gate296inter0), .b(s_298), .O(gate296inter1));
  and2  gate2635(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2636(.a(s_298), .O(gate296inter3));
  inv1  gate2637(.a(s_299), .O(gate296inter4));
  nand2 gate2638(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2639(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2640(.a(G826), .O(gate296inter7));
  inv1  gate2641(.a(G827), .O(gate296inter8));
  nand2 gate2642(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2643(.a(s_299), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2644(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2645(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2646(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate687(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate688(.a(gate387inter0), .b(s_20), .O(gate387inter1));
  and2  gate689(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate690(.a(s_20), .O(gate387inter3));
  inv1  gate691(.a(s_21), .O(gate387inter4));
  nand2 gate692(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate693(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate694(.a(G1), .O(gate387inter7));
  inv1  gate695(.a(G1036), .O(gate387inter8));
  nand2 gate696(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate697(.a(s_21), .b(gate387inter3), .O(gate387inter10));
  nor2  gate698(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate699(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate700(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate3011(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate3012(.a(gate392inter0), .b(s_352), .O(gate392inter1));
  and2  gate3013(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate3014(.a(s_352), .O(gate392inter3));
  inv1  gate3015(.a(s_353), .O(gate392inter4));
  nand2 gate3016(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate3017(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate3018(.a(G6), .O(gate392inter7));
  inv1  gate3019(.a(G1051), .O(gate392inter8));
  nand2 gate3020(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate3021(.a(s_353), .b(gate392inter3), .O(gate392inter10));
  nor2  gate3022(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate3023(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate3024(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate2157(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate2158(.a(gate393inter0), .b(s_230), .O(gate393inter1));
  and2  gate2159(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate2160(.a(s_230), .O(gate393inter3));
  inv1  gate2161(.a(s_231), .O(gate393inter4));
  nand2 gate2162(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate2163(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate2164(.a(G7), .O(gate393inter7));
  inv1  gate2165(.a(G1054), .O(gate393inter8));
  nand2 gate2166(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate2167(.a(s_231), .b(gate393inter3), .O(gate393inter10));
  nor2  gate2168(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate2169(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate2170(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2549(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2550(.a(gate394inter0), .b(s_286), .O(gate394inter1));
  and2  gate2551(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2552(.a(s_286), .O(gate394inter3));
  inv1  gate2553(.a(s_287), .O(gate394inter4));
  nand2 gate2554(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2555(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2556(.a(G8), .O(gate394inter7));
  inv1  gate2557(.a(G1057), .O(gate394inter8));
  nand2 gate2558(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2559(.a(s_287), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2560(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2561(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2562(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate2031(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2032(.a(gate395inter0), .b(s_212), .O(gate395inter1));
  and2  gate2033(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2034(.a(s_212), .O(gate395inter3));
  inv1  gate2035(.a(s_213), .O(gate395inter4));
  nand2 gate2036(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2037(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2038(.a(G9), .O(gate395inter7));
  inv1  gate2039(.a(G1060), .O(gate395inter8));
  nand2 gate2040(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2041(.a(s_213), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2042(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2043(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2044(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2493(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2494(.a(gate396inter0), .b(s_278), .O(gate396inter1));
  and2  gate2495(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2496(.a(s_278), .O(gate396inter3));
  inv1  gate2497(.a(s_279), .O(gate396inter4));
  nand2 gate2498(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2499(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2500(.a(G10), .O(gate396inter7));
  inv1  gate2501(.a(G1063), .O(gate396inter8));
  nand2 gate2502(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2503(.a(s_279), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2504(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2505(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2506(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate1261(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1262(.a(gate397inter0), .b(s_102), .O(gate397inter1));
  and2  gate1263(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1264(.a(s_102), .O(gate397inter3));
  inv1  gate1265(.a(s_103), .O(gate397inter4));
  nand2 gate1266(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1267(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1268(.a(G11), .O(gate397inter7));
  inv1  gate1269(.a(G1066), .O(gate397inter8));
  nand2 gate1270(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1271(.a(s_103), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1272(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1273(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1274(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate743(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate744(.a(gate399inter0), .b(s_28), .O(gate399inter1));
  and2  gate745(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate746(.a(s_28), .O(gate399inter3));
  inv1  gate747(.a(s_29), .O(gate399inter4));
  nand2 gate748(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate749(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate750(.a(G13), .O(gate399inter7));
  inv1  gate751(.a(G1072), .O(gate399inter8));
  nand2 gate752(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate753(.a(s_29), .b(gate399inter3), .O(gate399inter10));
  nor2  gate754(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate755(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate756(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1079(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1080(.a(gate402inter0), .b(s_76), .O(gate402inter1));
  and2  gate1081(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1082(.a(s_76), .O(gate402inter3));
  inv1  gate1083(.a(s_77), .O(gate402inter4));
  nand2 gate1084(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1085(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1086(.a(G16), .O(gate402inter7));
  inv1  gate1087(.a(G1081), .O(gate402inter8));
  nand2 gate1088(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1089(.a(s_77), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1090(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1091(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1092(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1611(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1612(.a(gate403inter0), .b(s_152), .O(gate403inter1));
  and2  gate1613(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1614(.a(s_152), .O(gate403inter3));
  inv1  gate1615(.a(s_153), .O(gate403inter4));
  nand2 gate1616(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1617(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1618(.a(G17), .O(gate403inter7));
  inv1  gate1619(.a(G1084), .O(gate403inter8));
  nand2 gate1620(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1621(.a(s_153), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1622(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1623(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1624(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1639(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1640(.a(gate404inter0), .b(s_156), .O(gate404inter1));
  and2  gate1641(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1642(.a(s_156), .O(gate404inter3));
  inv1  gate1643(.a(s_157), .O(gate404inter4));
  nand2 gate1644(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1645(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1646(.a(G18), .O(gate404inter7));
  inv1  gate1647(.a(G1087), .O(gate404inter8));
  nand2 gate1648(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1649(.a(s_157), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1650(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1651(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1652(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate3193(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate3194(.a(gate406inter0), .b(s_378), .O(gate406inter1));
  and2  gate3195(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate3196(.a(s_378), .O(gate406inter3));
  inv1  gate3197(.a(s_379), .O(gate406inter4));
  nand2 gate3198(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate3199(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate3200(.a(G20), .O(gate406inter7));
  inv1  gate3201(.a(G1093), .O(gate406inter8));
  nand2 gate3202(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate3203(.a(s_379), .b(gate406inter3), .O(gate406inter10));
  nor2  gate3204(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate3205(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate3206(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2129(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2130(.a(gate408inter0), .b(s_226), .O(gate408inter1));
  and2  gate2131(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2132(.a(s_226), .O(gate408inter3));
  inv1  gate2133(.a(s_227), .O(gate408inter4));
  nand2 gate2134(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2135(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2136(.a(G22), .O(gate408inter7));
  inv1  gate2137(.a(G1099), .O(gate408inter8));
  nand2 gate2138(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2139(.a(s_227), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2140(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2141(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2142(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate2143(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2144(.a(gate409inter0), .b(s_228), .O(gate409inter1));
  and2  gate2145(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2146(.a(s_228), .O(gate409inter3));
  inv1  gate2147(.a(s_229), .O(gate409inter4));
  nand2 gate2148(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2149(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2150(.a(G23), .O(gate409inter7));
  inv1  gate2151(.a(G1102), .O(gate409inter8));
  nand2 gate2152(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2153(.a(s_229), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2154(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2155(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2156(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1457(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1458(.a(gate410inter0), .b(s_130), .O(gate410inter1));
  and2  gate1459(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1460(.a(s_130), .O(gate410inter3));
  inv1  gate1461(.a(s_131), .O(gate410inter4));
  nand2 gate1462(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1463(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1464(.a(G24), .O(gate410inter7));
  inv1  gate1465(.a(G1105), .O(gate410inter8));
  nand2 gate1466(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1467(.a(s_131), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1468(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1469(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1470(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate785(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate786(.a(gate412inter0), .b(s_34), .O(gate412inter1));
  and2  gate787(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate788(.a(s_34), .O(gate412inter3));
  inv1  gate789(.a(s_35), .O(gate412inter4));
  nand2 gate790(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate791(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate792(.a(G26), .O(gate412inter7));
  inv1  gate793(.a(G1111), .O(gate412inter8));
  nand2 gate794(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate795(.a(s_35), .b(gate412inter3), .O(gate412inter10));
  nor2  gate796(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate797(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate798(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate967(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate968(.a(gate413inter0), .b(s_60), .O(gate413inter1));
  and2  gate969(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate970(.a(s_60), .O(gate413inter3));
  inv1  gate971(.a(s_61), .O(gate413inter4));
  nand2 gate972(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate973(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate974(.a(G27), .O(gate413inter7));
  inv1  gate975(.a(G1114), .O(gate413inter8));
  nand2 gate976(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate977(.a(s_61), .b(gate413inter3), .O(gate413inter10));
  nor2  gate978(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate979(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate980(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate1135(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1136(.a(gate414inter0), .b(s_84), .O(gate414inter1));
  and2  gate1137(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1138(.a(s_84), .O(gate414inter3));
  inv1  gate1139(.a(s_85), .O(gate414inter4));
  nand2 gate1140(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1141(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1142(.a(G28), .O(gate414inter7));
  inv1  gate1143(.a(G1117), .O(gate414inter8));
  nand2 gate1144(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1145(.a(s_85), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1146(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1147(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1148(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate2899(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2900(.a(gate415inter0), .b(s_336), .O(gate415inter1));
  and2  gate2901(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2902(.a(s_336), .O(gate415inter3));
  inv1  gate2903(.a(s_337), .O(gate415inter4));
  nand2 gate2904(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2905(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2906(.a(G29), .O(gate415inter7));
  inv1  gate2907(.a(G1120), .O(gate415inter8));
  nand2 gate2908(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2909(.a(s_337), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2910(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2911(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2912(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2997(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2998(.a(gate418inter0), .b(s_350), .O(gate418inter1));
  and2  gate2999(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate3000(.a(s_350), .O(gate418inter3));
  inv1  gate3001(.a(s_351), .O(gate418inter4));
  nand2 gate3002(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate3003(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate3004(.a(G32), .O(gate418inter7));
  inv1  gate3005(.a(G1129), .O(gate418inter8));
  nand2 gate3006(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate3007(.a(s_351), .b(gate418inter3), .O(gate418inter10));
  nor2  gate3008(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate3009(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate3010(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate2381(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2382(.a(gate422inter0), .b(s_262), .O(gate422inter1));
  and2  gate2383(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2384(.a(s_262), .O(gate422inter3));
  inv1  gate2385(.a(s_263), .O(gate422inter4));
  nand2 gate2386(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2387(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2388(.a(G1039), .O(gate422inter7));
  inv1  gate2389(.a(G1135), .O(gate422inter8));
  nand2 gate2390(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2391(.a(s_263), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2392(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2393(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2394(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate897(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate898(.a(gate425inter0), .b(s_50), .O(gate425inter1));
  and2  gate899(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate900(.a(s_50), .O(gate425inter3));
  inv1  gate901(.a(s_51), .O(gate425inter4));
  nand2 gate902(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate903(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate904(.a(G4), .O(gate425inter7));
  inv1  gate905(.a(G1141), .O(gate425inter8));
  nand2 gate906(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate907(.a(s_51), .b(gate425inter3), .O(gate425inter10));
  nor2  gate908(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate909(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate910(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1219(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1220(.a(gate426inter0), .b(s_96), .O(gate426inter1));
  and2  gate1221(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1222(.a(s_96), .O(gate426inter3));
  inv1  gate1223(.a(s_97), .O(gate426inter4));
  nand2 gate1224(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1225(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1226(.a(G1045), .O(gate426inter7));
  inv1  gate1227(.a(G1141), .O(gate426inter8));
  nand2 gate1228(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1229(.a(s_97), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1230(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1231(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1232(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1289(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1290(.a(gate429inter0), .b(s_106), .O(gate429inter1));
  and2  gate1291(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1292(.a(s_106), .O(gate429inter3));
  inv1  gate1293(.a(s_107), .O(gate429inter4));
  nand2 gate1294(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1295(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1296(.a(G6), .O(gate429inter7));
  inv1  gate1297(.a(G1147), .O(gate429inter8));
  nand2 gate1298(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1299(.a(s_107), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1300(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1301(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1302(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1093(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1094(.a(gate431inter0), .b(s_78), .O(gate431inter1));
  and2  gate1095(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1096(.a(s_78), .O(gate431inter3));
  inv1  gate1097(.a(s_79), .O(gate431inter4));
  nand2 gate1098(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1099(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1100(.a(G7), .O(gate431inter7));
  inv1  gate1101(.a(G1150), .O(gate431inter8));
  nand2 gate1102(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1103(.a(s_79), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1104(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1105(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1106(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate2745(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2746(.a(gate433inter0), .b(s_314), .O(gate433inter1));
  and2  gate2747(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2748(.a(s_314), .O(gate433inter3));
  inv1  gate2749(.a(s_315), .O(gate433inter4));
  nand2 gate2750(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2751(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2752(.a(G8), .O(gate433inter7));
  inv1  gate2753(.a(G1153), .O(gate433inter8));
  nand2 gate2754(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2755(.a(s_315), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2756(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2757(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2758(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1037(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1038(.a(gate434inter0), .b(s_70), .O(gate434inter1));
  and2  gate1039(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1040(.a(s_70), .O(gate434inter3));
  inv1  gate1041(.a(s_71), .O(gate434inter4));
  nand2 gate1042(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1043(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1044(.a(G1057), .O(gate434inter7));
  inv1  gate1045(.a(G1153), .O(gate434inter8));
  nand2 gate1046(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1047(.a(s_71), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1048(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1049(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1050(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1961(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1962(.a(gate440inter0), .b(s_202), .O(gate440inter1));
  and2  gate1963(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1964(.a(s_202), .O(gate440inter3));
  inv1  gate1965(.a(s_203), .O(gate440inter4));
  nand2 gate1966(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1967(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1968(.a(G1066), .O(gate440inter7));
  inv1  gate1969(.a(G1162), .O(gate440inter8));
  nand2 gate1970(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1971(.a(s_203), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1972(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1973(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1974(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1583(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1584(.a(gate443inter0), .b(s_148), .O(gate443inter1));
  and2  gate1585(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1586(.a(s_148), .O(gate443inter3));
  inv1  gate1587(.a(s_149), .O(gate443inter4));
  nand2 gate1588(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1589(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1590(.a(G13), .O(gate443inter7));
  inv1  gate1591(.a(G1168), .O(gate443inter8));
  nand2 gate1592(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1593(.a(s_149), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1594(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1595(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1596(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1443(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1444(.a(gate445inter0), .b(s_128), .O(gate445inter1));
  and2  gate1445(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1446(.a(s_128), .O(gate445inter3));
  inv1  gate1447(.a(s_129), .O(gate445inter4));
  nand2 gate1448(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1449(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1450(.a(G14), .O(gate445inter7));
  inv1  gate1451(.a(G1171), .O(gate445inter8));
  nand2 gate1452(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1453(.a(s_129), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1454(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1455(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1456(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate631(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate632(.a(gate446inter0), .b(s_12), .O(gate446inter1));
  and2  gate633(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate634(.a(s_12), .O(gate446inter3));
  inv1  gate635(.a(s_13), .O(gate446inter4));
  nand2 gate636(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate637(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate638(.a(G1075), .O(gate446inter7));
  inv1  gate639(.a(G1171), .O(gate446inter8));
  nand2 gate640(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate641(.a(s_13), .b(gate446inter3), .O(gate446inter10));
  nor2  gate642(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate643(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate644(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1765(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1766(.a(gate448inter0), .b(s_174), .O(gate448inter1));
  and2  gate1767(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1768(.a(s_174), .O(gate448inter3));
  inv1  gate1769(.a(s_175), .O(gate448inter4));
  nand2 gate1770(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1771(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1772(.a(G1078), .O(gate448inter7));
  inv1  gate1773(.a(G1174), .O(gate448inter8));
  nand2 gate1774(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1775(.a(s_175), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1776(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1777(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1778(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2885(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2886(.a(gate449inter0), .b(s_334), .O(gate449inter1));
  and2  gate2887(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2888(.a(s_334), .O(gate449inter3));
  inv1  gate2889(.a(s_335), .O(gate449inter4));
  nand2 gate2890(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2891(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2892(.a(G16), .O(gate449inter7));
  inv1  gate2893(.a(G1177), .O(gate449inter8));
  nand2 gate2894(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2895(.a(s_335), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2896(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2897(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2898(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate2661(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2662(.a(gate457inter0), .b(s_302), .O(gate457inter1));
  and2  gate2663(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2664(.a(s_302), .O(gate457inter3));
  inv1  gate2665(.a(s_303), .O(gate457inter4));
  nand2 gate2666(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2667(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2668(.a(G20), .O(gate457inter7));
  inv1  gate2669(.a(G1189), .O(gate457inter8));
  nand2 gate2670(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2671(.a(s_303), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2672(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2673(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2674(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate547(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate548(.a(gate459inter0), .b(s_0), .O(gate459inter1));
  and2  gate549(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate550(.a(s_0), .O(gate459inter3));
  inv1  gate551(.a(s_1), .O(gate459inter4));
  nand2 gate552(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate553(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate554(.a(G21), .O(gate459inter7));
  inv1  gate555(.a(G1192), .O(gate459inter8));
  nand2 gate556(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate557(.a(s_1), .b(gate459inter3), .O(gate459inter10));
  nor2  gate558(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate559(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate560(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2675(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2676(.a(gate461inter0), .b(s_304), .O(gate461inter1));
  and2  gate2677(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2678(.a(s_304), .O(gate461inter3));
  inv1  gate2679(.a(s_305), .O(gate461inter4));
  nand2 gate2680(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2681(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2682(.a(G22), .O(gate461inter7));
  inv1  gate2683(.a(G1195), .O(gate461inter8));
  nand2 gate2684(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2685(.a(s_305), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2686(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2687(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2688(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2969(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2970(.a(gate464inter0), .b(s_346), .O(gate464inter1));
  and2  gate2971(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2972(.a(s_346), .O(gate464inter3));
  inv1  gate2973(.a(s_347), .O(gate464inter4));
  nand2 gate2974(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2975(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2976(.a(G1102), .O(gate464inter7));
  inv1  gate2977(.a(G1198), .O(gate464inter8));
  nand2 gate2978(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2979(.a(s_347), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2980(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2981(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2982(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1527(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1528(.a(gate465inter0), .b(s_140), .O(gate465inter1));
  and2  gate1529(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1530(.a(s_140), .O(gate465inter3));
  inv1  gate1531(.a(s_141), .O(gate465inter4));
  nand2 gate1532(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1533(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1534(.a(G24), .O(gate465inter7));
  inv1  gate1535(.a(G1201), .O(gate465inter8));
  nand2 gate1536(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1537(.a(s_141), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1538(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1539(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1540(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1065(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1066(.a(gate466inter0), .b(s_74), .O(gate466inter1));
  and2  gate1067(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1068(.a(s_74), .O(gate466inter3));
  inv1  gate1069(.a(s_75), .O(gate466inter4));
  nand2 gate1070(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1071(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1072(.a(G1105), .O(gate466inter7));
  inv1  gate1073(.a(G1201), .O(gate466inter8));
  nand2 gate1074(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1075(.a(s_75), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1076(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1077(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1078(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1947(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1948(.a(gate467inter0), .b(s_200), .O(gate467inter1));
  and2  gate1949(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1950(.a(s_200), .O(gate467inter3));
  inv1  gate1951(.a(s_201), .O(gate467inter4));
  nand2 gate1952(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1953(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1954(.a(G25), .O(gate467inter7));
  inv1  gate1955(.a(G1204), .O(gate467inter8));
  nand2 gate1956(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1957(.a(s_201), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1958(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1959(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1960(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2647(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2648(.a(gate469inter0), .b(s_300), .O(gate469inter1));
  and2  gate2649(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2650(.a(s_300), .O(gate469inter3));
  inv1  gate2651(.a(s_301), .O(gate469inter4));
  nand2 gate2652(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2653(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2654(.a(G26), .O(gate469inter7));
  inv1  gate2655(.a(G1207), .O(gate469inter8));
  nand2 gate2656(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2657(.a(s_301), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2658(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2659(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2660(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate701(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate702(.a(gate470inter0), .b(s_22), .O(gate470inter1));
  and2  gate703(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate704(.a(s_22), .O(gate470inter3));
  inv1  gate705(.a(s_23), .O(gate470inter4));
  nand2 gate706(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate707(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate708(.a(G1111), .O(gate470inter7));
  inv1  gate709(.a(G1207), .O(gate470inter8));
  nand2 gate710(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate711(.a(s_23), .b(gate470inter3), .O(gate470inter10));
  nor2  gate712(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate713(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate714(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate2591(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2592(.a(gate472inter0), .b(s_292), .O(gate472inter1));
  and2  gate2593(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2594(.a(s_292), .O(gate472inter3));
  inv1  gate2595(.a(s_293), .O(gate472inter4));
  nand2 gate2596(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2597(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2598(.a(G1114), .O(gate472inter7));
  inv1  gate2599(.a(G1210), .O(gate472inter8));
  nand2 gate2600(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2601(.a(s_293), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2602(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2603(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2604(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1233(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1234(.a(gate485inter0), .b(s_98), .O(gate485inter1));
  and2  gate1235(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1236(.a(s_98), .O(gate485inter3));
  inv1  gate1237(.a(s_99), .O(gate485inter4));
  nand2 gate1238(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1239(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1240(.a(G1232), .O(gate485inter7));
  inv1  gate1241(.a(G1233), .O(gate485inter8));
  nand2 gate1242(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1243(.a(s_99), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1244(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1245(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1246(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1345(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1346(.a(gate487inter0), .b(s_114), .O(gate487inter1));
  and2  gate1347(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1348(.a(s_114), .O(gate487inter3));
  inv1  gate1349(.a(s_115), .O(gate487inter4));
  nand2 gate1350(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1351(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1352(.a(G1236), .O(gate487inter7));
  inv1  gate1353(.a(G1237), .O(gate487inter8));
  nand2 gate1354(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1355(.a(s_115), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1356(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1357(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1358(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate939(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate940(.a(gate493inter0), .b(s_56), .O(gate493inter1));
  and2  gate941(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate942(.a(s_56), .O(gate493inter3));
  inv1  gate943(.a(s_57), .O(gate493inter4));
  nand2 gate944(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate945(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate946(.a(G1248), .O(gate493inter7));
  inv1  gate947(.a(G1249), .O(gate493inter8));
  nand2 gate948(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate949(.a(s_57), .b(gate493inter3), .O(gate493inter10));
  nor2  gate950(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate951(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate952(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1779(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1780(.a(gate494inter0), .b(s_176), .O(gate494inter1));
  and2  gate1781(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1782(.a(s_176), .O(gate494inter3));
  inv1  gate1783(.a(s_177), .O(gate494inter4));
  nand2 gate1784(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1785(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1786(.a(G1250), .O(gate494inter7));
  inv1  gate1787(.a(G1251), .O(gate494inter8));
  nand2 gate1788(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1789(.a(s_177), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1790(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1791(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1792(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2073(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2074(.a(gate497inter0), .b(s_218), .O(gate497inter1));
  and2  gate2075(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2076(.a(s_218), .O(gate497inter3));
  inv1  gate2077(.a(s_219), .O(gate497inter4));
  nand2 gate2078(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2079(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2080(.a(G1256), .O(gate497inter7));
  inv1  gate2081(.a(G1257), .O(gate497inter8));
  nand2 gate2082(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2083(.a(s_219), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2084(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2085(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2086(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1905(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1906(.a(gate498inter0), .b(s_194), .O(gate498inter1));
  and2  gate1907(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1908(.a(s_194), .O(gate498inter3));
  inv1  gate1909(.a(s_195), .O(gate498inter4));
  nand2 gate1910(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1911(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1912(.a(G1258), .O(gate498inter7));
  inv1  gate1913(.a(G1259), .O(gate498inter8));
  nand2 gate1914(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1915(.a(s_195), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1916(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1917(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1918(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1359(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1360(.a(gate499inter0), .b(s_116), .O(gate499inter1));
  and2  gate1361(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1362(.a(s_116), .O(gate499inter3));
  inv1  gate1363(.a(s_117), .O(gate499inter4));
  nand2 gate1364(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1365(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1366(.a(G1260), .O(gate499inter7));
  inv1  gate1367(.a(G1261), .O(gate499inter8));
  nand2 gate1368(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1369(.a(s_117), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1370(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1371(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1372(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1303(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1304(.a(gate501inter0), .b(s_108), .O(gate501inter1));
  and2  gate1305(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1306(.a(s_108), .O(gate501inter3));
  inv1  gate1307(.a(s_109), .O(gate501inter4));
  nand2 gate1308(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1309(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1310(.a(G1264), .O(gate501inter7));
  inv1  gate1311(.a(G1265), .O(gate501inter8));
  nand2 gate1312(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1313(.a(s_109), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1314(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1315(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1316(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1919(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1920(.a(gate502inter0), .b(s_196), .O(gate502inter1));
  and2  gate1921(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1922(.a(s_196), .O(gate502inter3));
  inv1  gate1923(.a(s_197), .O(gate502inter4));
  nand2 gate1924(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1925(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1926(.a(G1266), .O(gate502inter7));
  inv1  gate1927(.a(G1267), .O(gate502inter8));
  nand2 gate1928(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1929(.a(s_197), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1930(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1931(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1932(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate2297(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2298(.a(gate504inter0), .b(s_250), .O(gate504inter1));
  and2  gate2299(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2300(.a(s_250), .O(gate504inter3));
  inv1  gate2301(.a(s_251), .O(gate504inter4));
  nand2 gate2302(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2303(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2304(.a(G1270), .O(gate504inter7));
  inv1  gate2305(.a(G1271), .O(gate504inter8));
  nand2 gate2306(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2307(.a(s_251), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2308(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2309(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2310(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2535(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2536(.a(gate507inter0), .b(s_284), .O(gate507inter1));
  and2  gate2537(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2538(.a(s_284), .O(gate507inter3));
  inv1  gate2539(.a(s_285), .O(gate507inter4));
  nand2 gate2540(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2541(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2542(.a(G1276), .O(gate507inter7));
  inv1  gate2543(.a(G1277), .O(gate507inter8));
  nand2 gate2544(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2545(.a(s_285), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2546(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2547(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2548(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1569(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1570(.a(gate508inter0), .b(s_146), .O(gate508inter1));
  and2  gate1571(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1572(.a(s_146), .O(gate508inter3));
  inv1  gate1573(.a(s_147), .O(gate508inter4));
  nand2 gate1574(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1575(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1576(.a(G1278), .O(gate508inter7));
  inv1  gate1577(.a(G1279), .O(gate508inter8));
  nand2 gate1578(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1579(.a(s_147), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1580(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1581(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1582(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2017(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2018(.a(gate510inter0), .b(s_210), .O(gate510inter1));
  and2  gate2019(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2020(.a(s_210), .O(gate510inter3));
  inv1  gate2021(.a(s_211), .O(gate510inter4));
  nand2 gate2022(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2023(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2024(.a(G1282), .O(gate510inter7));
  inv1  gate2025(.a(G1283), .O(gate510inter8));
  nand2 gate2026(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2027(.a(s_211), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2028(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2029(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2030(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1247(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1248(.a(gate513inter0), .b(s_100), .O(gate513inter1));
  and2  gate1249(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1250(.a(s_100), .O(gate513inter3));
  inv1  gate1251(.a(s_101), .O(gate513inter4));
  nand2 gate1252(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1253(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1254(.a(G1288), .O(gate513inter7));
  inv1  gate1255(.a(G1289), .O(gate513inter8));
  nand2 gate1256(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1257(.a(s_101), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1258(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1259(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1260(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule