module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate2675(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2676(.a(gate10inter0), .b(s_304), .O(gate10inter1));
  and2  gate2677(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2678(.a(s_304), .O(gate10inter3));
  inv1  gate2679(.a(s_305), .O(gate10inter4));
  nand2 gate2680(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2681(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2682(.a(G3), .O(gate10inter7));
  inv1  gate2683(.a(G4), .O(gate10inter8));
  nand2 gate2684(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2685(.a(s_305), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2686(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2687(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2688(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1331(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1332(.a(gate12inter0), .b(s_112), .O(gate12inter1));
  and2  gate1333(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1334(.a(s_112), .O(gate12inter3));
  inv1  gate1335(.a(s_113), .O(gate12inter4));
  nand2 gate1336(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1337(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1338(.a(G7), .O(gate12inter7));
  inv1  gate1339(.a(G8), .O(gate12inter8));
  nand2 gate1340(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1341(.a(s_113), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1342(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1343(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1344(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1485(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1486(.a(gate13inter0), .b(s_134), .O(gate13inter1));
  and2  gate1487(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1488(.a(s_134), .O(gate13inter3));
  inv1  gate1489(.a(s_135), .O(gate13inter4));
  nand2 gate1490(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1491(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1492(.a(G9), .O(gate13inter7));
  inv1  gate1493(.a(G10), .O(gate13inter8));
  nand2 gate1494(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1495(.a(s_135), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1496(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1497(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1498(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate617(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate618(.a(gate22inter0), .b(s_10), .O(gate22inter1));
  and2  gate619(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate620(.a(s_10), .O(gate22inter3));
  inv1  gate621(.a(s_11), .O(gate22inter4));
  nand2 gate622(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate623(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate624(.a(G27), .O(gate22inter7));
  inv1  gate625(.a(G28), .O(gate22inter8));
  nand2 gate626(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate627(.a(s_11), .b(gate22inter3), .O(gate22inter10));
  nor2  gate628(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate629(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate630(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2661(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2662(.a(gate25inter0), .b(s_302), .O(gate25inter1));
  and2  gate2663(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2664(.a(s_302), .O(gate25inter3));
  inv1  gate2665(.a(s_303), .O(gate25inter4));
  nand2 gate2666(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2667(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2668(.a(G1), .O(gate25inter7));
  inv1  gate2669(.a(G5), .O(gate25inter8));
  nand2 gate2670(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2671(.a(s_303), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2672(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2673(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2674(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate813(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate814(.a(gate31inter0), .b(s_38), .O(gate31inter1));
  and2  gate815(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate816(.a(s_38), .O(gate31inter3));
  inv1  gate817(.a(s_39), .O(gate31inter4));
  nand2 gate818(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate819(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate820(.a(G4), .O(gate31inter7));
  inv1  gate821(.a(G8), .O(gate31inter8));
  nand2 gate822(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate823(.a(s_39), .b(gate31inter3), .O(gate31inter10));
  nor2  gate824(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate825(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate826(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1569(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1570(.a(gate32inter0), .b(s_146), .O(gate32inter1));
  and2  gate1571(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1572(.a(s_146), .O(gate32inter3));
  inv1  gate1573(.a(s_147), .O(gate32inter4));
  nand2 gate1574(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1575(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1576(.a(G12), .O(gate32inter7));
  inv1  gate1577(.a(G16), .O(gate32inter8));
  nand2 gate1578(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1579(.a(s_147), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1580(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1581(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1582(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2311(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2312(.a(gate34inter0), .b(s_252), .O(gate34inter1));
  and2  gate2313(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2314(.a(s_252), .O(gate34inter3));
  inv1  gate2315(.a(s_253), .O(gate34inter4));
  nand2 gate2316(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2317(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2318(.a(G25), .O(gate34inter7));
  inv1  gate2319(.a(G29), .O(gate34inter8));
  nand2 gate2320(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2321(.a(s_253), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2322(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2323(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2324(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1723(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1724(.a(gate36inter0), .b(s_168), .O(gate36inter1));
  and2  gate1725(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1726(.a(s_168), .O(gate36inter3));
  inv1  gate1727(.a(s_169), .O(gate36inter4));
  nand2 gate1728(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1729(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1730(.a(G26), .O(gate36inter7));
  inv1  gate1731(.a(G30), .O(gate36inter8));
  nand2 gate1732(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1733(.a(s_169), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1734(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1735(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1736(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate2255(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2256(.a(gate40inter0), .b(s_244), .O(gate40inter1));
  and2  gate2257(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2258(.a(s_244), .O(gate40inter3));
  inv1  gate2259(.a(s_245), .O(gate40inter4));
  nand2 gate2260(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2261(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2262(.a(G28), .O(gate40inter7));
  inv1  gate2263(.a(G32), .O(gate40inter8));
  nand2 gate2264(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2265(.a(s_245), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2266(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2267(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2268(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2647(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2648(.a(gate42inter0), .b(s_300), .O(gate42inter1));
  and2  gate2649(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2650(.a(s_300), .O(gate42inter3));
  inv1  gate2651(.a(s_301), .O(gate42inter4));
  nand2 gate2652(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2653(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2654(.a(G2), .O(gate42inter7));
  inv1  gate2655(.a(G266), .O(gate42inter8));
  nand2 gate2656(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2657(.a(s_301), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2658(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2659(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2660(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2367(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2368(.a(gate46inter0), .b(s_260), .O(gate46inter1));
  and2  gate2369(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2370(.a(s_260), .O(gate46inter3));
  inv1  gate2371(.a(s_261), .O(gate46inter4));
  nand2 gate2372(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2373(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2374(.a(G6), .O(gate46inter7));
  inv1  gate2375(.a(G272), .O(gate46inter8));
  nand2 gate2376(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2377(.a(s_261), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2378(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2379(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2380(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1247(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1248(.a(gate51inter0), .b(s_100), .O(gate51inter1));
  and2  gate1249(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1250(.a(s_100), .O(gate51inter3));
  inv1  gate1251(.a(s_101), .O(gate51inter4));
  nand2 gate1252(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1253(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1254(.a(G11), .O(gate51inter7));
  inv1  gate1255(.a(G281), .O(gate51inter8));
  nand2 gate1256(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1257(.a(s_101), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1258(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1259(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1260(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2269(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2270(.a(gate58inter0), .b(s_246), .O(gate58inter1));
  and2  gate2271(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2272(.a(s_246), .O(gate58inter3));
  inv1  gate2273(.a(s_247), .O(gate58inter4));
  nand2 gate2274(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2275(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2276(.a(G18), .O(gate58inter7));
  inv1  gate2277(.a(G290), .O(gate58inter8));
  nand2 gate2278(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2279(.a(s_247), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2280(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2281(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2282(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1149(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1150(.a(gate65inter0), .b(s_86), .O(gate65inter1));
  and2  gate1151(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1152(.a(s_86), .O(gate65inter3));
  inv1  gate1153(.a(s_87), .O(gate65inter4));
  nand2 gate1154(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1155(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1156(.a(G25), .O(gate65inter7));
  inv1  gate1157(.a(G302), .O(gate65inter8));
  nand2 gate1158(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1159(.a(s_87), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1160(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1161(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1162(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate2423(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2424(.a(gate66inter0), .b(s_268), .O(gate66inter1));
  and2  gate2425(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2426(.a(s_268), .O(gate66inter3));
  inv1  gate2427(.a(s_269), .O(gate66inter4));
  nand2 gate2428(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2429(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2430(.a(G26), .O(gate66inter7));
  inv1  gate2431(.a(G302), .O(gate66inter8));
  nand2 gate2432(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2433(.a(s_269), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2434(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2435(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2436(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1793(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1794(.a(gate67inter0), .b(s_178), .O(gate67inter1));
  and2  gate1795(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1796(.a(s_178), .O(gate67inter3));
  inv1  gate1797(.a(s_179), .O(gate67inter4));
  nand2 gate1798(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1799(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1800(.a(G27), .O(gate67inter7));
  inv1  gate1801(.a(G305), .O(gate67inter8));
  nand2 gate1802(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1803(.a(s_179), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1804(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1805(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1806(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate2017(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2018(.a(gate68inter0), .b(s_210), .O(gate68inter1));
  and2  gate2019(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2020(.a(s_210), .O(gate68inter3));
  inv1  gate2021(.a(s_211), .O(gate68inter4));
  nand2 gate2022(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2023(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2024(.a(G28), .O(gate68inter7));
  inv1  gate2025(.a(G305), .O(gate68inter8));
  nand2 gate2026(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2027(.a(s_211), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2028(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2029(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2030(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate673(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate674(.a(gate69inter0), .b(s_18), .O(gate69inter1));
  and2  gate675(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate676(.a(s_18), .O(gate69inter3));
  inv1  gate677(.a(s_19), .O(gate69inter4));
  nand2 gate678(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate679(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate680(.a(G29), .O(gate69inter7));
  inv1  gate681(.a(G308), .O(gate69inter8));
  nand2 gate682(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate683(.a(s_19), .b(gate69inter3), .O(gate69inter10));
  nor2  gate684(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate685(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate686(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2003(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2004(.a(gate71inter0), .b(s_208), .O(gate71inter1));
  and2  gate2005(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2006(.a(s_208), .O(gate71inter3));
  inv1  gate2007(.a(s_209), .O(gate71inter4));
  nand2 gate2008(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2009(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2010(.a(G31), .O(gate71inter7));
  inv1  gate2011(.a(G311), .O(gate71inter8));
  nand2 gate2012(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2013(.a(s_209), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2014(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2015(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2016(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate2353(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2354(.a(gate75inter0), .b(s_258), .O(gate75inter1));
  and2  gate2355(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2356(.a(s_258), .O(gate75inter3));
  inv1  gate2357(.a(s_259), .O(gate75inter4));
  nand2 gate2358(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2359(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2360(.a(G9), .O(gate75inter7));
  inv1  gate2361(.a(G317), .O(gate75inter8));
  nand2 gate2362(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2363(.a(s_259), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2364(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2365(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2366(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2241(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2242(.a(gate79inter0), .b(s_242), .O(gate79inter1));
  and2  gate2243(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2244(.a(s_242), .O(gate79inter3));
  inv1  gate2245(.a(s_243), .O(gate79inter4));
  nand2 gate2246(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2247(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2248(.a(G10), .O(gate79inter7));
  inv1  gate2249(.a(G323), .O(gate79inter8));
  nand2 gate2250(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2251(.a(s_243), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2252(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2253(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2254(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate575(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate576(.a(gate80inter0), .b(s_4), .O(gate80inter1));
  and2  gate577(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate578(.a(s_4), .O(gate80inter3));
  inv1  gate579(.a(s_5), .O(gate80inter4));
  nand2 gate580(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate581(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate582(.a(G14), .O(gate80inter7));
  inv1  gate583(.a(G323), .O(gate80inter8));
  nand2 gate584(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate585(.a(s_5), .b(gate80inter3), .O(gate80inter10));
  nor2  gate586(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate587(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate588(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2101(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2102(.a(gate82inter0), .b(s_222), .O(gate82inter1));
  and2  gate2103(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2104(.a(s_222), .O(gate82inter3));
  inv1  gate2105(.a(s_223), .O(gate82inter4));
  nand2 gate2106(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2107(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2108(.a(G7), .O(gate82inter7));
  inv1  gate2109(.a(G326), .O(gate82inter8));
  nand2 gate2110(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2111(.a(s_223), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2112(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2113(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2114(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate1905(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1906(.a(gate83inter0), .b(s_194), .O(gate83inter1));
  and2  gate1907(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1908(.a(s_194), .O(gate83inter3));
  inv1  gate1909(.a(s_195), .O(gate83inter4));
  nand2 gate1910(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1911(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1912(.a(G11), .O(gate83inter7));
  inv1  gate1913(.a(G329), .O(gate83inter8));
  nand2 gate1914(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1915(.a(s_195), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1916(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1917(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1918(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1429(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1430(.a(gate86inter0), .b(s_126), .O(gate86inter1));
  and2  gate1431(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1432(.a(s_126), .O(gate86inter3));
  inv1  gate1433(.a(s_127), .O(gate86inter4));
  nand2 gate1434(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1435(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1436(.a(G8), .O(gate86inter7));
  inv1  gate1437(.a(G332), .O(gate86inter8));
  nand2 gate1438(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1439(.a(s_127), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1440(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1441(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1442(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2563(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2564(.a(gate87inter0), .b(s_288), .O(gate87inter1));
  and2  gate2565(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2566(.a(s_288), .O(gate87inter3));
  inv1  gate2567(.a(s_289), .O(gate87inter4));
  nand2 gate2568(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2569(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2570(.a(G12), .O(gate87inter7));
  inv1  gate2571(.a(G335), .O(gate87inter8));
  nand2 gate2572(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2573(.a(s_289), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2574(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2575(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2576(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2479(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2480(.a(gate90inter0), .b(s_276), .O(gate90inter1));
  and2  gate2481(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2482(.a(s_276), .O(gate90inter3));
  inv1  gate2483(.a(s_277), .O(gate90inter4));
  nand2 gate2484(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2485(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2486(.a(G21), .O(gate90inter7));
  inv1  gate2487(.a(G338), .O(gate90inter8));
  nand2 gate2488(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2489(.a(s_277), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2490(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2491(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2492(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1695(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1696(.a(gate94inter0), .b(s_164), .O(gate94inter1));
  and2  gate1697(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1698(.a(s_164), .O(gate94inter3));
  inv1  gate1699(.a(s_165), .O(gate94inter4));
  nand2 gate1700(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1701(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1702(.a(G22), .O(gate94inter7));
  inv1  gate1703(.a(G344), .O(gate94inter8));
  nand2 gate1704(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1705(.a(s_165), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1706(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1707(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1708(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate687(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate688(.a(gate95inter0), .b(s_20), .O(gate95inter1));
  and2  gate689(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate690(.a(s_20), .O(gate95inter3));
  inv1  gate691(.a(s_21), .O(gate95inter4));
  nand2 gate692(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate693(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate694(.a(G26), .O(gate95inter7));
  inv1  gate695(.a(G347), .O(gate95inter8));
  nand2 gate696(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate697(.a(s_21), .b(gate95inter3), .O(gate95inter10));
  nor2  gate698(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate699(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate700(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1863(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1864(.a(gate100inter0), .b(s_188), .O(gate100inter1));
  and2  gate1865(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1866(.a(s_188), .O(gate100inter3));
  inv1  gate1867(.a(s_189), .O(gate100inter4));
  nand2 gate1868(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1869(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1870(.a(G31), .O(gate100inter7));
  inv1  gate1871(.a(G353), .O(gate100inter8));
  nand2 gate1872(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1873(.a(s_189), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1874(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1875(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1876(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate799(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate800(.a(gate101inter0), .b(s_36), .O(gate101inter1));
  and2  gate801(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate802(.a(s_36), .O(gate101inter3));
  inv1  gate803(.a(s_37), .O(gate101inter4));
  nand2 gate804(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate805(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate806(.a(G20), .O(gate101inter7));
  inv1  gate807(.a(G356), .O(gate101inter8));
  nand2 gate808(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate809(.a(s_37), .b(gate101inter3), .O(gate101inter10));
  nor2  gate810(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate811(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate812(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate771(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate772(.a(gate102inter0), .b(s_32), .O(gate102inter1));
  and2  gate773(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate774(.a(s_32), .O(gate102inter3));
  inv1  gate775(.a(s_33), .O(gate102inter4));
  nand2 gate776(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate777(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate778(.a(G24), .O(gate102inter7));
  inv1  gate779(.a(G356), .O(gate102inter8));
  nand2 gate780(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate781(.a(s_33), .b(gate102inter3), .O(gate102inter10));
  nor2  gate782(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate783(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate784(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1513(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1514(.a(gate107inter0), .b(s_138), .O(gate107inter1));
  and2  gate1515(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1516(.a(s_138), .O(gate107inter3));
  inv1  gate1517(.a(s_139), .O(gate107inter4));
  nand2 gate1518(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1519(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1520(.a(G366), .O(gate107inter7));
  inv1  gate1521(.a(G367), .O(gate107inter8));
  nand2 gate1522(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1523(.a(s_139), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1524(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1525(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1526(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate2843(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2844(.a(gate108inter0), .b(s_328), .O(gate108inter1));
  and2  gate2845(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2846(.a(s_328), .O(gate108inter3));
  inv1  gate2847(.a(s_329), .O(gate108inter4));
  nand2 gate2848(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2849(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2850(.a(G368), .O(gate108inter7));
  inv1  gate2851(.a(G369), .O(gate108inter8));
  nand2 gate2852(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2853(.a(s_329), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2854(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2855(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2856(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate2129(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2130(.a(gate109inter0), .b(s_226), .O(gate109inter1));
  and2  gate2131(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2132(.a(s_226), .O(gate109inter3));
  inv1  gate2133(.a(s_227), .O(gate109inter4));
  nand2 gate2134(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2135(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2136(.a(G370), .O(gate109inter7));
  inv1  gate2137(.a(G371), .O(gate109inter8));
  nand2 gate2138(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2139(.a(s_227), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2140(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2141(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2142(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1373(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1374(.a(gate110inter0), .b(s_118), .O(gate110inter1));
  and2  gate1375(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1376(.a(s_118), .O(gate110inter3));
  inv1  gate1377(.a(s_119), .O(gate110inter4));
  nand2 gate1378(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1379(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1380(.a(G372), .O(gate110inter7));
  inv1  gate1381(.a(G373), .O(gate110inter8));
  nand2 gate1382(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1383(.a(s_119), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1384(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1385(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1386(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1009(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1010(.a(gate116inter0), .b(s_66), .O(gate116inter1));
  and2  gate1011(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1012(.a(s_66), .O(gate116inter3));
  inv1  gate1013(.a(s_67), .O(gate116inter4));
  nand2 gate1014(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1015(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1016(.a(G384), .O(gate116inter7));
  inv1  gate1017(.a(G385), .O(gate116inter8));
  nand2 gate1018(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1019(.a(s_67), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1020(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1021(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1022(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2717(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2718(.a(gate118inter0), .b(s_310), .O(gate118inter1));
  and2  gate2719(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2720(.a(s_310), .O(gate118inter3));
  inv1  gate2721(.a(s_311), .O(gate118inter4));
  nand2 gate2722(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2723(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2724(.a(G388), .O(gate118inter7));
  inv1  gate2725(.a(G389), .O(gate118inter8));
  nand2 gate2726(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2727(.a(s_311), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2728(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2729(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2730(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1807(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1808(.a(gate121inter0), .b(s_180), .O(gate121inter1));
  and2  gate1809(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1810(.a(s_180), .O(gate121inter3));
  inv1  gate1811(.a(s_181), .O(gate121inter4));
  nand2 gate1812(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1813(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1814(.a(G394), .O(gate121inter7));
  inv1  gate1815(.a(G395), .O(gate121inter8));
  nand2 gate1816(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1817(.a(s_181), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1818(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1819(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1820(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1527(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1528(.a(gate125inter0), .b(s_140), .O(gate125inter1));
  and2  gate1529(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1530(.a(s_140), .O(gate125inter3));
  inv1  gate1531(.a(s_141), .O(gate125inter4));
  nand2 gate1532(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1533(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1534(.a(G402), .O(gate125inter7));
  inv1  gate1535(.a(G403), .O(gate125inter8));
  nand2 gate1536(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1537(.a(s_141), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1538(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1539(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1540(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate2745(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2746(.a(gate126inter0), .b(s_314), .O(gate126inter1));
  and2  gate2747(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2748(.a(s_314), .O(gate126inter3));
  inv1  gate2749(.a(s_315), .O(gate126inter4));
  nand2 gate2750(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2751(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2752(.a(G404), .O(gate126inter7));
  inv1  gate2753(.a(G405), .O(gate126inter8));
  nand2 gate2754(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2755(.a(s_315), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2756(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2757(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2758(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate2213(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2214(.a(gate127inter0), .b(s_238), .O(gate127inter1));
  and2  gate2215(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2216(.a(s_238), .O(gate127inter3));
  inv1  gate2217(.a(s_239), .O(gate127inter4));
  nand2 gate2218(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2219(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2220(.a(G406), .O(gate127inter7));
  inv1  gate2221(.a(G407), .O(gate127inter8));
  nand2 gate2222(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2223(.a(s_239), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2224(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2225(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2226(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate939(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate940(.a(gate131inter0), .b(s_56), .O(gate131inter1));
  and2  gate941(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate942(.a(s_56), .O(gate131inter3));
  inv1  gate943(.a(s_57), .O(gate131inter4));
  nand2 gate944(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate945(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate946(.a(G414), .O(gate131inter7));
  inv1  gate947(.a(G415), .O(gate131inter8));
  nand2 gate948(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate949(.a(s_57), .b(gate131inter3), .O(gate131inter10));
  nor2  gate950(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate951(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate952(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate953(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate954(.a(gate135inter0), .b(s_58), .O(gate135inter1));
  and2  gate955(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate956(.a(s_58), .O(gate135inter3));
  inv1  gate957(.a(s_59), .O(gate135inter4));
  nand2 gate958(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate959(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate960(.a(G422), .O(gate135inter7));
  inv1  gate961(.a(G423), .O(gate135inter8));
  nand2 gate962(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate963(.a(s_59), .b(gate135inter3), .O(gate135inter10));
  nor2  gate964(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate965(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate966(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1023(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1024(.a(gate138inter0), .b(s_68), .O(gate138inter1));
  and2  gate1025(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1026(.a(s_68), .O(gate138inter3));
  inv1  gate1027(.a(s_69), .O(gate138inter4));
  nand2 gate1028(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1029(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1030(.a(G432), .O(gate138inter7));
  inv1  gate1031(.a(G435), .O(gate138inter8));
  nand2 gate1032(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1033(.a(s_69), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1034(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1035(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1036(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate701(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate702(.a(gate139inter0), .b(s_22), .O(gate139inter1));
  and2  gate703(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate704(.a(s_22), .O(gate139inter3));
  inv1  gate705(.a(s_23), .O(gate139inter4));
  nand2 gate706(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate707(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate708(.a(G438), .O(gate139inter7));
  inv1  gate709(.a(G441), .O(gate139inter8));
  nand2 gate710(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate711(.a(s_23), .b(gate139inter3), .O(gate139inter10));
  nor2  gate712(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate713(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate714(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1625(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1626(.a(gate140inter0), .b(s_154), .O(gate140inter1));
  and2  gate1627(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1628(.a(s_154), .O(gate140inter3));
  inv1  gate1629(.a(s_155), .O(gate140inter4));
  nand2 gate1630(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1631(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1632(.a(G444), .O(gate140inter7));
  inv1  gate1633(.a(G447), .O(gate140inter8));
  nand2 gate1634(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1635(.a(s_155), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1636(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1637(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1638(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1737(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1738(.a(gate141inter0), .b(s_170), .O(gate141inter1));
  and2  gate1739(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1740(.a(s_170), .O(gate141inter3));
  inv1  gate1741(.a(s_171), .O(gate141inter4));
  nand2 gate1742(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1743(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1744(.a(G450), .O(gate141inter7));
  inv1  gate1745(.a(G453), .O(gate141inter8));
  nand2 gate1746(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1747(.a(s_171), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1748(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1749(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1750(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate925(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate926(.a(gate150inter0), .b(s_54), .O(gate150inter1));
  and2  gate927(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate928(.a(s_54), .O(gate150inter3));
  inv1  gate929(.a(s_55), .O(gate150inter4));
  nand2 gate930(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate931(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate932(.a(G504), .O(gate150inter7));
  inv1  gate933(.a(G507), .O(gate150inter8));
  nand2 gate934(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate935(.a(s_55), .b(gate150inter3), .O(gate150inter10));
  nor2  gate936(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate937(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate938(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1401(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1402(.a(gate155inter0), .b(s_122), .O(gate155inter1));
  and2  gate1403(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1404(.a(s_122), .O(gate155inter3));
  inv1  gate1405(.a(s_123), .O(gate155inter4));
  nand2 gate1406(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1407(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1408(.a(G432), .O(gate155inter7));
  inv1  gate1409(.a(G525), .O(gate155inter8));
  nand2 gate1410(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1411(.a(s_123), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1412(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1413(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1414(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1205(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1206(.a(gate156inter0), .b(s_94), .O(gate156inter1));
  and2  gate1207(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1208(.a(s_94), .O(gate156inter3));
  inv1  gate1209(.a(s_95), .O(gate156inter4));
  nand2 gate1210(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1211(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1212(.a(G435), .O(gate156inter7));
  inv1  gate1213(.a(G525), .O(gate156inter8));
  nand2 gate1214(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1215(.a(s_95), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1216(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1217(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1218(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2619(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2620(.a(gate161inter0), .b(s_296), .O(gate161inter1));
  and2  gate2621(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2622(.a(s_296), .O(gate161inter3));
  inv1  gate2623(.a(s_297), .O(gate161inter4));
  nand2 gate2624(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2625(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2626(.a(G450), .O(gate161inter7));
  inv1  gate2627(.a(G534), .O(gate161inter8));
  nand2 gate2628(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2629(.a(s_297), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2630(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2631(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2632(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate2409(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2410(.a(gate162inter0), .b(s_266), .O(gate162inter1));
  and2  gate2411(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2412(.a(s_266), .O(gate162inter3));
  inv1  gate2413(.a(s_267), .O(gate162inter4));
  nand2 gate2414(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2415(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2416(.a(G453), .O(gate162inter7));
  inv1  gate2417(.a(G534), .O(gate162inter8));
  nand2 gate2418(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2419(.a(s_267), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2420(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2421(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2422(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate547(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate548(.a(gate166inter0), .b(s_0), .O(gate166inter1));
  and2  gate549(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate550(.a(s_0), .O(gate166inter3));
  inv1  gate551(.a(s_1), .O(gate166inter4));
  nand2 gate552(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate553(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate554(.a(G465), .O(gate166inter7));
  inv1  gate555(.a(G540), .O(gate166inter8));
  nand2 gate556(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate557(.a(s_1), .b(gate166inter3), .O(gate166inter10));
  nor2  gate558(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate559(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate560(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate981(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate982(.a(gate168inter0), .b(s_62), .O(gate168inter1));
  and2  gate983(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate984(.a(s_62), .O(gate168inter3));
  inv1  gate985(.a(s_63), .O(gate168inter4));
  nand2 gate986(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate987(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate988(.a(G471), .O(gate168inter7));
  inv1  gate989(.a(G543), .O(gate168inter8));
  nand2 gate990(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate991(.a(s_63), .b(gate168inter3), .O(gate168inter10));
  nor2  gate992(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate993(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate994(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1975(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1976(.a(gate171inter0), .b(s_204), .O(gate171inter1));
  and2  gate1977(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1978(.a(s_204), .O(gate171inter3));
  inv1  gate1979(.a(s_205), .O(gate171inter4));
  nand2 gate1980(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1981(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1982(.a(G480), .O(gate171inter7));
  inv1  gate1983(.a(G549), .O(gate171inter8));
  nand2 gate1984(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1985(.a(s_205), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1986(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1987(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1988(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1289(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1290(.a(gate173inter0), .b(s_106), .O(gate173inter1));
  and2  gate1291(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1292(.a(s_106), .O(gate173inter3));
  inv1  gate1293(.a(s_107), .O(gate173inter4));
  nand2 gate1294(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1295(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1296(.a(G486), .O(gate173inter7));
  inv1  gate1297(.a(G552), .O(gate173inter8));
  nand2 gate1298(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1299(.a(s_107), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1300(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1301(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1302(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate967(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate968(.a(gate180inter0), .b(s_60), .O(gate180inter1));
  and2  gate969(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate970(.a(s_60), .O(gate180inter3));
  inv1  gate971(.a(s_61), .O(gate180inter4));
  nand2 gate972(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate973(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate974(.a(G507), .O(gate180inter7));
  inv1  gate975(.a(G561), .O(gate180inter8));
  nand2 gate976(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate977(.a(s_61), .b(gate180inter3), .O(gate180inter10));
  nor2  gate978(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate979(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate980(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1471(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1472(.a(gate181inter0), .b(s_132), .O(gate181inter1));
  and2  gate1473(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1474(.a(s_132), .O(gate181inter3));
  inv1  gate1475(.a(s_133), .O(gate181inter4));
  nand2 gate1476(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1477(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1478(.a(G510), .O(gate181inter7));
  inv1  gate1479(.a(G564), .O(gate181inter8));
  nand2 gate1480(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1481(.a(s_133), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1482(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1483(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1484(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2731(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2732(.a(gate182inter0), .b(s_312), .O(gate182inter1));
  and2  gate2733(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2734(.a(s_312), .O(gate182inter3));
  inv1  gate2735(.a(s_313), .O(gate182inter4));
  nand2 gate2736(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2737(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2738(.a(G513), .O(gate182inter7));
  inv1  gate2739(.a(G564), .O(gate182inter8));
  nand2 gate2740(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2741(.a(s_313), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2742(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2743(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2744(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate2521(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2522(.a(gate184inter0), .b(s_282), .O(gate184inter1));
  and2  gate2523(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2524(.a(s_282), .O(gate184inter3));
  inv1  gate2525(.a(s_283), .O(gate184inter4));
  nand2 gate2526(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2527(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2528(.a(G519), .O(gate184inter7));
  inv1  gate2529(.a(G567), .O(gate184inter8));
  nand2 gate2530(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2531(.a(s_283), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2532(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2533(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2534(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2199(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2200(.a(gate190inter0), .b(s_236), .O(gate190inter1));
  and2  gate2201(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2202(.a(s_236), .O(gate190inter3));
  inv1  gate2203(.a(s_237), .O(gate190inter4));
  nand2 gate2204(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2205(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2206(.a(G580), .O(gate190inter7));
  inv1  gate2207(.a(G581), .O(gate190inter8));
  nand2 gate2208(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2209(.a(s_237), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2210(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2211(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2212(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate1891(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1892(.a(gate191inter0), .b(s_192), .O(gate191inter1));
  and2  gate1893(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1894(.a(s_192), .O(gate191inter3));
  inv1  gate1895(.a(s_193), .O(gate191inter4));
  nand2 gate1896(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1897(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1898(.a(G582), .O(gate191inter7));
  inv1  gate1899(.a(G583), .O(gate191inter8));
  nand2 gate1900(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1901(.a(s_193), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1902(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1903(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1904(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1499(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1500(.a(gate192inter0), .b(s_136), .O(gate192inter1));
  and2  gate1501(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1502(.a(s_136), .O(gate192inter3));
  inv1  gate1503(.a(s_137), .O(gate192inter4));
  nand2 gate1504(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1505(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1506(.a(G584), .O(gate192inter7));
  inv1  gate1507(.a(G585), .O(gate192inter8));
  nand2 gate1508(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1509(.a(s_137), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1510(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1511(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1512(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2283(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2284(.a(gate198inter0), .b(s_248), .O(gate198inter1));
  and2  gate2285(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2286(.a(s_248), .O(gate198inter3));
  inv1  gate2287(.a(s_249), .O(gate198inter4));
  nand2 gate2288(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2289(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2290(.a(G596), .O(gate198inter7));
  inv1  gate2291(.a(G597), .O(gate198inter8));
  nand2 gate2292(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2293(.a(s_249), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2294(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2295(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2296(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1275(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1276(.a(gate199inter0), .b(s_104), .O(gate199inter1));
  and2  gate1277(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1278(.a(s_104), .O(gate199inter3));
  inv1  gate1279(.a(s_105), .O(gate199inter4));
  nand2 gate1280(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1281(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1282(.a(G598), .O(gate199inter7));
  inv1  gate1283(.a(G599), .O(gate199inter8));
  nand2 gate1284(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1285(.a(s_105), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1286(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1287(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1288(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1387(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1388(.a(gate200inter0), .b(s_120), .O(gate200inter1));
  and2  gate1389(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1390(.a(s_120), .O(gate200inter3));
  inv1  gate1391(.a(s_121), .O(gate200inter4));
  nand2 gate1392(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1393(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1394(.a(G600), .O(gate200inter7));
  inv1  gate1395(.a(G601), .O(gate200inter8));
  nand2 gate1396(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1397(.a(s_121), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1398(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1399(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1400(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate2031(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2032(.a(gate201inter0), .b(s_212), .O(gate201inter1));
  and2  gate2033(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2034(.a(s_212), .O(gate201inter3));
  inv1  gate2035(.a(s_213), .O(gate201inter4));
  nand2 gate2036(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2037(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2038(.a(G602), .O(gate201inter7));
  inv1  gate2039(.a(G607), .O(gate201inter8));
  nand2 gate2040(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2041(.a(s_213), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2042(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2043(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2044(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1933(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1934(.a(gate202inter0), .b(s_198), .O(gate202inter1));
  and2  gate1935(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1936(.a(s_198), .O(gate202inter3));
  inv1  gate1937(.a(s_199), .O(gate202inter4));
  nand2 gate1938(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1939(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1940(.a(G612), .O(gate202inter7));
  inv1  gate1941(.a(G617), .O(gate202inter8));
  nand2 gate1942(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1943(.a(s_199), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1944(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1945(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1946(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate659(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate660(.a(gate203inter0), .b(s_16), .O(gate203inter1));
  and2  gate661(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate662(.a(s_16), .O(gate203inter3));
  inv1  gate663(.a(s_17), .O(gate203inter4));
  nand2 gate664(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate665(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate666(.a(G602), .O(gate203inter7));
  inv1  gate667(.a(G612), .O(gate203inter8));
  nand2 gate668(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate669(.a(s_17), .b(gate203inter3), .O(gate203inter10));
  nor2  gate670(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate671(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate672(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1415(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1416(.a(gate206inter0), .b(s_124), .O(gate206inter1));
  and2  gate1417(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1418(.a(s_124), .O(gate206inter3));
  inv1  gate1419(.a(s_125), .O(gate206inter4));
  nand2 gate1420(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1421(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1422(.a(G632), .O(gate206inter7));
  inv1  gate1423(.a(G637), .O(gate206inter8));
  nand2 gate1424(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1425(.a(s_125), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1426(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1427(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1428(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1177(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1178(.a(gate209inter0), .b(s_90), .O(gate209inter1));
  and2  gate1179(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1180(.a(s_90), .O(gate209inter3));
  inv1  gate1181(.a(s_91), .O(gate209inter4));
  nand2 gate1182(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1183(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1184(.a(G602), .O(gate209inter7));
  inv1  gate1185(.a(G666), .O(gate209inter8));
  nand2 gate1186(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1187(.a(s_91), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1188(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1189(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1190(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2227(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2228(.a(gate213inter0), .b(s_240), .O(gate213inter1));
  and2  gate2229(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2230(.a(s_240), .O(gate213inter3));
  inv1  gate2231(.a(s_241), .O(gate213inter4));
  nand2 gate2232(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2233(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2234(.a(G602), .O(gate213inter7));
  inv1  gate2235(.a(G672), .O(gate213inter8));
  nand2 gate2236(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2237(.a(s_241), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2238(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2239(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2240(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2591(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2592(.a(gate214inter0), .b(s_292), .O(gate214inter1));
  and2  gate2593(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2594(.a(s_292), .O(gate214inter3));
  inv1  gate2595(.a(s_293), .O(gate214inter4));
  nand2 gate2596(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2597(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2598(.a(G612), .O(gate214inter7));
  inv1  gate2599(.a(G672), .O(gate214inter8));
  nand2 gate2600(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2601(.a(s_293), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2602(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2603(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2604(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate883(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate884(.a(gate216inter0), .b(s_48), .O(gate216inter1));
  and2  gate885(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate886(.a(s_48), .O(gate216inter3));
  inv1  gate887(.a(s_49), .O(gate216inter4));
  nand2 gate888(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate889(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate890(.a(G617), .O(gate216inter7));
  inv1  gate891(.a(G675), .O(gate216inter8));
  nand2 gate892(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate893(.a(s_49), .b(gate216inter3), .O(gate216inter10));
  nor2  gate894(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate895(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate896(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate995(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate996(.a(gate218inter0), .b(s_64), .O(gate218inter1));
  and2  gate997(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate998(.a(s_64), .O(gate218inter3));
  inv1  gate999(.a(s_65), .O(gate218inter4));
  nand2 gate1000(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1001(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1002(.a(G627), .O(gate218inter7));
  inv1  gate1003(.a(G678), .O(gate218inter8));
  nand2 gate1004(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1005(.a(s_65), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1006(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1007(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1008(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate589(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate590(.a(gate222inter0), .b(s_6), .O(gate222inter1));
  and2  gate591(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate592(.a(s_6), .O(gate222inter3));
  inv1  gate593(.a(s_7), .O(gate222inter4));
  nand2 gate594(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate595(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate596(.a(G632), .O(gate222inter7));
  inv1  gate597(.a(G684), .O(gate222inter8));
  nand2 gate598(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate599(.a(s_7), .b(gate222inter3), .O(gate222inter10));
  nor2  gate600(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate601(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate602(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1051(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1052(.a(gate224inter0), .b(s_72), .O(gate224inter1));
  and2  gate1053(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1054(.a(s_72), .O(gate224inter3));
  inv1  gate1055(.a(s_73), .O(gate224inter4));
  nand2 gate1056(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1057(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1058(.a(G637), .O(gate224inter7));
  inv1  gate1059(.a(G687), .O(gate224inter8));
  nand2 gate1060(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1061(.a(s_73), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1062(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1063(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1064(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate2143(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2144(.a(gate225inter0), .b(s_228), .O(gate225inter1));
  and2  gate2145(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2146(.a(s_228), .O(gate225inter3));
  inv1  gate2147(.a(s_229), .O(gate225inter4));
  nand2 gate2148(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2149(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2150(.a(G690), .O(gate225inter7));
  inv1  gate2151(.a(G691), .O(gate225inter8));
  nand2 gate2152(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2153(.a(s_229), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2154(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2155(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2156(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1233(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1234(.a(gate227inter0), .b(s_98), .O(gate227inter1));
  and2  gate1235(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1236(.a(s_98), .O(gate227inter3));
  inv1  gate1237(.a(s_99), .O(gate227inter4));
  nand2 gate1238(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1239(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1240(.a(G694), .O(gate227inter7));
  inv1  gate1241(.a(G695), .O(gate227inter8));
  nand2 gate1242(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1243(.a(s_99), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1244(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1245(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1246(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate827(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate828(.a(gate228inter0), .b(s_40), .O(gate228inter1));
  and2  gate829(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate830(.a(s_40), .O(gate228inter3));
  inv1  gate831(.a(s_41), .O(gate228inter4));
  nand2 gate832(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate833(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate834(.a(G696), .O(gate228inter7));
  inv1  gate835(.a(G697), .O(gate228inter8));
  nand2 gate836(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate837(.a(s_41), .b(gate228inter3), .O(gate228inter10));
  nor2  gate838(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate839(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate840(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1667(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1668(.a(gate231inter0), .b(s_160), .O(gate231inter1));
  and2  gate1669(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1670(.a(s_160), .O(gate231inter3));
  inv1  gate1671(.a(s_161), .O(gate231inter4));
  nand2 gate1672(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1673(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1674(.a(G702), .O(gate231inter7));
  inv1  gate1675(.a(G703), .O(gate231inter8));
  nand2 gate1676(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1677(.a(s_161), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1678(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1679(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1680(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1457(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1458(.a(gate233inter0), .b(s_130), .O(gate233inter1));
  and2  gate1459(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1460(.a(s_130), .O(gate233inter3));
  inv1  gate1461(.a(s_131), .O(gate233inter4));
  nand2 gate1462(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1463(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1464(.a(G242), .O(gate233inter7));
  inv1  gate1465(.a(G718), .O(gate233inter8));
  nand2 gate1466(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1467(.a(s_131), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1468(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1469(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1470(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate785(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate786(.a(gate234inter0), .b(s_34), .O(gate234inter1));
  and2  gate787(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate788(.a(s_34), .O(gate234inter3));
  inv1  gate789(.a(s_35), .O(gate234inter4));
  nand2 gate790(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate791(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate792(.a(G245), .O(gate234inter7));
  inv1  gate793(.a(G721), .O(gate234inter8));
  nand2 gate794(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate795(.a(s_35), .b(gate234inter3), .O(gate234inter10));
  nor2  gate796(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate797(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate798(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2829(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2830(.a(gate235inter0), .b(s_326), .O(gate235inter1));
  and2  gate2831(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2832(.a(s_326), .O(gate235inter3));
  inv1  gate2833(.a(s_327), .O(gate235inter4));
  nand2 gate2834(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2835(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2836(.a(G248), .O(gate235inter7));
  inv1  gate2837(.a(G724), .O(gate235inter8));
  nand2 gate2838(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2839(.a(s_327), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2840(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2841(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2842(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate715(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate716(.a(gate236inter0), .b(s_24), .O(gate236inter1));
  and2  gate717(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate718(.a(s_24), .O(gate236inter3));
  inv1  gate719(.a(s_25), .O(gate236inter4));
  nand2 gate720(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate721(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate722(.a(G251), .O(gate236inter7));
  inv1  gate723(.a(G727), .O(gate236inter8));
  nand2 gate724(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate725(.a(s_25), .b(gate236inter3), .O(gate236inter10));
  nor2  gate726(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate727(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate728(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1835(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1836(.a(gate237inter0), .b(s_184), .O(gate237inter1));
  and2  gate1837(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1838(.a(s_184), .O(gate237inter3));
  inv1  gate1839(.a(s_185), .O(gate237inter4));
  nand2 gate1840(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1841(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1842(.a(G254), .O(gate237inter7));
  inv1  gate1843(.a(G706), .O(gate237inter8));
  nand2 gate1844(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1845(.a(s_185), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1846(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1847(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1848(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1345(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1346(.a(gate238inter0), .b(s_114), .O(gate238inter1));
  and2  gate1347(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1348(.a(s_114), .O(gate238inter3));
  inv1  gate1349(.a(s_115), .O(gate238inter4));
  nand2 gate1350(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1351(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1352(.a(G257), .O(gate238inter7));
  inv1  gate1353(.a(G709), .O(gate238inter8));
  nand2 gate1354(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1355(.a(s_115), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1356(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1357(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1358(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1303(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1304(.a(gate243inter0), .b(s_108), .O(gate243inter1));
  and2  gate1305(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1306(.a(s_108), .O(gate243inter3));
  inv1  gate1307(.a(s_109), .O(gate243inter4));
  nand2 gate1308(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1309(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1310(.a(G245), .O(gate243inter7));
  inv1  gate1311(.a(G733), .O(gate243inter8));
  nand2 gate1312(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1313(.a(s_109), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1314(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1315(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1316(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1093(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1094(.a(gate244inter0), .b(s_78), .O(gate244inter1));
  and2  gate1095(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1096(.a(s_78), .O(gate244inter3));
  inv1  gate1097(.a(s_79), .O(gate244inter4));
  nand2 gate1098(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1099(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1100(.a(G721), .O(gate244inter7));
  inv1  gate1101(.a(G733), .O(gate244inter8));
  nand2 gate1102(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1103(.a(s_79), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1104(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1105(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1106(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate2437(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2438(.a(gate247inter0), .b(s_270), .O(gate247inter1));
  and2  gate2439(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2440(.a(s_270), .O(gate247inter3));
  inv1  gate2441(.a(s_271), .O(gate247inter4));
  nand2 gate2442(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2443(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2444(.a(G251), .O(gate247inter7));
  inv1  gate2445(.a(G739), .O(gate247inter8));
  nand2 gate2446(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2447(.a(s_271), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2448(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2449(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2450(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1919(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1920(.a(gate248inter0), .b(s_196), .O(gate248inter1));
  and2  gate1921(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1922(.a(s_196), .O(gate248inter3));
  inv1  gate1923(.a(s_197), .O(gate248inter4));
  nand2 gate1924(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1925(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1926(.a(G727), .O(gate248inter7));
  inv1  gate1927(.a(G739), .O(gate248inter8));
  nand2 gate1928(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1929(.a(s_197), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1930(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1931(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1932(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2815(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2816(.a(gate252inter0), .b(s_324), .O(gate252inter1));
  and2  gate2817(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2818(.a(s_324), .O(gate252inter3));
  inv1  gate2819(.a(s_325), .O(gate252inter4));
  nand2 gate2820(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2821(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2822(.a(G709), .O(gate252inter7));
  inv1  gate2823(.a(G745), .O(gate252inter8));
  nand2 gate2824(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2825(.a(s_325), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2826(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2827(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2828(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate645(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate646(.a(gate253inter0), .b(s_14), .O(gate253inter1));
  and2  gate647(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate648(.a(s_14), .O(gate253inter3));
  inv1  gate649(.a(s_15), .O(gate253inter4));
  nand2 gate650(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate651(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate652(.a(G260), .O(gate253inter7));
  inv1  gate653(.a(G748), .O(gate253inter8));
  nand2 gate654(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate655(.a(s_15), .b(gate253inter3), .O(gate253inter10));
  nor2  gate656(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate657(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate658(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1849(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1850(.a(gate257inter0), .b(s_186), .O(gate257inter1));
  and2  gate1851(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1852(.a(s_186), .O(gate257inter3));
  inv1  gate1853(.a(s_187), .O(gate257inter4));
  nand2 gate1854(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1855(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1856(.a(G754), .O(gate257inter7));
  inv1  gate1857(.a(G755), .O(gate257inter8));
  nand2 gate1858(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1859(.a(s_187), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1860(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1861(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1862(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate2115(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2116(.a(gate258inter0), .b(s_224), .O(gate258inter1));
  and2  gate2117(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2118(.a(s_224), .O(gate258inter3));
  inv1  gate2119(.a(s_225), .O(gate258inter4));
  nand2 gate2120(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2121(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2122(.a(G756), .O(gate258inter7));
  inv1  gate2123(.a(G757), .O(gate258inter8));
  nand2 gate2124(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2125(.a(s_225), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2126(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2127(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2128(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1359(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1360(.a(gate263inter0), .b(s_116), .O(gate263inter1));
  and2  gate1361(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1362(.a(s_116), .O(gate263inter3));
  inv1  gate1363(.a(s_117), .O(gate263inter4));
  nand2 gate1364(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1365(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1366(.a(G766), .O(gate263inter7));
  inv1  gate1367(.a(G767), .O(gate263inter8));
  nand2 gate1368(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1369(.a(s_117), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1370(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1371(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1372(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1163(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1164(.a(gate266inter0), .b(s_88), .O(gate266inter1));
  and2  gate1165(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1166(.a(s_88), .O(gate266inter3));
  inv1  gate1167(.a(s_89), .O(gate266inter4));
  nand2 gate1168(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1169(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1170(.a(G645), .O(gate266inter7));
  inv1  gate1171(.a(G773), .O(gate266inter8));
  nand2 gate1172(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1173(.a(s_89), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1174(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1175(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1176(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2087(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2088(.a(gate269inter0), .b(s_220), .O(gate269inter1));
  and2  gate2089(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2090(.a(s_220), .O(gate269inter3));
  inv1  gate2091(.a(s_221), .O(gate269inter4));
  nand2 gate2092(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2093(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2094(.a(G654), .O(gate269inter7));
  inv1  gate2095(.a(G782), .O(gate269inter8));
  nand2 gate2096(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2097(.a(s_221), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2098(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2099(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2100(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate1135(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1136(.a(gate270inter0), .b(s_84), .O(gate270inter1));
  and2  gate1137(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1138(.a(s_84), .O(gate270inter3));
  inv1  gate1139(.a(s_85), .O(gate270inter4));
  nand2 gate1140(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1141(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1142(.a(G657), .O(gate270inter7));
  inv1  gate1143(.a(G785), .O(gate270inter8));
  nand2 gate1144(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1145(.a(s_85), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1146(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1147(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1148(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1709(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1710(.a(gate276inter0), .b(s_166), .O(gate276inter1));
  and2  gate1711(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1712(.a(s_166), .O(gate276inter3));
  inv1  gate1713(.a(s_167), .O(gate276inter4));
  nand2 gate1714(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1715(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1716(.a(G773), .O(gate276inter7));
  inv1  gate1717(.a(G797), .O(gate276inter8));
  nand2 gate1718(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1719(.a(s_167), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1720(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1721(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1722(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1751(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1752(.a(gate277inter0), .b(s_172), .O(gate277inter1));
  and2  gate1753(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1754(.a(s_172), .O(gate277inter3));
  inv1  gate1755(.a(s_173), .O(gate277inter4));
  nand2 gate1756(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1757(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1758(.a(G648), .O(gate277inter7));
  inv1  gate1759(.a(G800), .O(gate277inter8));
  nand2 gate1760(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1761(.a(s_173), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1762(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1763(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1764(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate2381(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2382(.a(gate278inter0), .b(s_262), .O(gate278inter1));
  and2  gate2383(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2384(.a(s_262), .O(gate278inter3));
  inv1  gate2385(.a(s_263), .O(gate278inter4));
  nand2 gate2386(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2387(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2388(.a(G776), .O(gate278inter7));
  inv1  gate2389(.a(G800), .O(gate278inter8));
  nand2 gate2390(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2391(.a(s_263), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2392(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2393(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2394(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2185(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2186(.a(gate281inter0), .b(s_234), .O(gate281inter1));
  and2  gate2187(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2188(.a(s_234), .O(gate281inter3));
  inv1  gate2189(.a(s_235), .O(gate281inter4));
  nand2 gate2190(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2191(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2192(.a(G654), .O(gate281inter7));
  inv1  gate2193(.a(G806), .O(gate281inter8));
  nand2 gate2194(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2195(.a(s_235), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2196(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2197(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2198(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate911(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate912(.a(gate284inter0), .b(s_52), .O(gate284inter1));
  and2  gate913(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate914(.a(s_52), .O(gate284inter3));
  inv1  gate915(.a(s_53), .O(gate284inter4));
  nand2 gate916(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate917(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate918(.a(G785), .O(gate284inter7));
  inv1  gate919(.a(G809), .O(gate284inter8));
  nand2 gate920(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate921(.a(s_53), .b(gate284inter3), .O(gate284inter10));
  nor2  gate922(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate923(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate924(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2857(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2858(.a(gate287inter0), .b(s_330), .O(gate287inter1));
  and2  gate2859(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2860(.a(s_330), .O(gate287inter3));
  inv1  gate2861(.a(s_331), .O(gate287inter4));
  nand2 gate2862(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2863(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2864(.a(G663), .O(gate287inter7));
  inv1  gate2865(.a(G815), .O(gate287inter8));
  nand2 gate2866(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2867(.a(s_331), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2868(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2869(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2870(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate2689(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2690(.a(gate288inter0), .b(s_306), .O(gate288inter1));
  and2  gate2691(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2692(.a(s_306), .O(gate288inter3));
  inv1  gate2693(.a(s_307), .O(gate288inter4));
  nand2 gate2694(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2695(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2696(.a(G791), .O(gate288inter7));
  inv1  gate2697(.a(G815), .O(gate288inter8));
  nand2 gate2698(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2699(.a(s_307), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2700(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2701(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2702(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate729(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate730(.a(gate289inter0), .b(s_26), .O(gate289inter1));
  and2  gate731(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate732(.a(s_26), .O(gate289inter3));
  inv1  gate733(.a(s_27), .O(gate289inter4));
  nand2 gate734(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate735(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate736(.a(G818), .O(gate289inter7));
  inv1  gate737(.a(G819), .O(gate289inter8));
  nand2 gate738(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate739(.a(s_27), .b(gate289inter3), .O(gate289inter10));
  nor2  gate740(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate741(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate742(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2605(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2606(.a(gate291inter0), .b(s_294), .O(gate291inter1));
  and2  gate2607(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2608(.a(s_294), .O(gate291inter3));
  inv1  gate2609(.a(s_295), .O(gate291inter4));
  nand2 gate2610(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2611(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2612(.a(G822), .O(gate291inter7));
  inv1  gate2613(.a(G823), .O(gate291inter8));
  nand2 gate2614(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2615(.a(s_295), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2616(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2617(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2618(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate2535(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2536(.a(gate292inter0), .b(s_284), .O(gate292inter1));
  and2  gate2537(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2538(.a(s_284), .O(gate292inter3));
  inv1  gate2539(.a(s_285), .O(gate292inter4));
  nand2 gate2540(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2541(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2542(.a(G824), .O(gate292inter7));
  inv1  gate2543(.a(G825), .O(gate292inter8));
  nand2 gate2544(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2545(.a(s_285), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2546(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2547(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2548(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1443(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1444(.a(gate293inter0), .b(s_128), .O(gate293inter1));
  and2  gate1445(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1446(.a(s_128), .O(gate293inter3));
  inv1  gate1447(.a(s_129), .O(gate293inter4));
  nand2 gate1448(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1449(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1450(.a(G828), .O(gate293inter7));
  inv1  gate1451(.a(G829), .O(gate293inter8));
  nand2 gate1452(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1453(.a(s_129), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1454(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1455(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1456(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1219(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1220(.a(gate388inter0), .b(s_96), .O(gate388inter1));
  and2  gate1221(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1222(.a(s_96), .O(gate388inter3));
  inv1  gate1223(.a(s_97), .O(gate388inter4));
  nand2 gate1224(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1225(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1226(.a(G2), .O(gate388inter7));
  inv1  gate1227(.a(G1039), .O(gate388inter8));
  nand2 gate1228(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1229(.a(s_97), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1230(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1231(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1232(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate2073(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2074(.a(gate390inter0), .b(s_218), .O(gate390inter1));
  and2  gate2075(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2076(.a(s_218), .O(gate390inter3));
  inv1  gate2077(.a(s_219), .O(gate390inter4));
  nand2 gate2078(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2079(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2080(.a(G4), .O(gate390inter7));
  inv1  gate2081(.a(G1045), .O(gate390inter8));
  nand2 gate2082(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2083(.a(s_219), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2084(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2085(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2086(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate2507(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2508(.a(gate391inter0), .b(s_280), .O(gate391inter1));
  and2  gate2509(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2510(.a(s_280), .O(gate391inter3));
  inv1  gate2511(.a(s_281), .O(gate391inter4));
  nand2 gate2512(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2513(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2514(.a(G5), .O(gate391inter7));
  inv1  gate2515(.a(G1048), .O(gate391inter8));
  nand2 gate2516(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2517(.a(s_281), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2518(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2519(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2520(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate743(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate744(.a(gate394inter0), .b(s_28), .O(gate394inter1));
  and2  gate745(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate746(.a(s_28), .O(gate394inter3));
  inv1  gate747(.a(s_29), .O(gate394inter4));
  nand2 gate748(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate749(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate750(.a(G8), .O(gate394inter7));
  inv1  gate751(.a(G1057), .O(gate394inter8));
  nand2 gate752(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate753(.a(s_29), .b(gate394inter3), .O(gate394inter10));
  nor2  gate754(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate755(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate756(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1681(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1682(.a(gate396inter0), .b(s_162), .O(gate396inter1));
  and2  gate1683(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1684(.a(s_162), .O(gate396inter3));
  inv1  gate1685(.a(s_163), .O(gate396inter4));
  nand2 gate1686(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1687(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1688(.a(G10), .O(gate396inter7));
  inv1  gate1689(.a(G1063), .O(gate396inter8));
  nand2 gate1690(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1691(.a(s_163), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1692(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1693(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1694(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1989(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1990(.a(gate398inter0), .b(s_206), .O(gate398inter1));
  and2  gate1991(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1992(.a(s_206), .O(gate398inter3));
  inv1  gate1993(.a(s_207), .O(gate398inter4));
  nand2 gate1994(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1995(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1996(.a(G12), .O(gate398inter7));
  inv1  gate1997(.a(G1069), .O(gate398inter8));
  nand2 gate1998(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1999(.a(s_207), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2000(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2001(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2002(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1583(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1584(.a(gate400inter0), .b(s_148), .O(gate400inter1));
  and2  gate1585(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1586(.a(s_148), .O(gate400inter3));
  inv1  gate1587(.a(s_149), .O(gate400inter4));
  nand2 gate1588(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1589(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1590(.a(G14), .O(gate400inter7));
  inv1  gate1591(.a(G1075), .O(gate400inter8));
  nand2 gate1592(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1593(.a(s_149), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1594(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1595(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1596(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1877(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1878(.a(gate404inter0), .b(s_190), .O(gate404inter1));
  and2  gate1879(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1880(.a(s_190), .O(gate404inter3));
  inv1  gate1881(.a(s_191), .O(gate404inter4));
  nand2 gate1882(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1883(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1884(.a(G18), .O(gate404inter7));
  inv1  gate1885(.a(G1087), .O(gate404inter8));
  nand2 gate1886(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1887(.a(s_191), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1888(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1889(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1890(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1121(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1122(.a(gate408inter0), .b(s_82), .O(gate408inter1));
  and2  gate1123(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1124(.a(s_82), .O(gate408inter3));
  inv1  gate1125(.a(s_83), .O(gate408inter4));
  nand2 gate1126(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1127(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1128(.a(G22), .O(gate408inter7));
  inv1  gate1129(.a(G1099), .O(gate408inter8));
  nand2 gate1130(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1131(.a(s_83), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1132(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1133(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1134(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1821(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1822(.a(gate409inter0), .b(s_182), .O(gate409inter1));
  and2  gate1823(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1824(.a(s_182), .O(gate409inter3));
  inv1  gate1825(.a(s_183), .O(gate409inter4));
  nand2 gate1826(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1827(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1828(.a(G23), .O(gate409inter7));
  inv1  gate1829(.a(G1102), .O(gate409inter8));
  nand2 gate1830(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1831(.a(s_183), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1832(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1833(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1834(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2549(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2550(.a(gate410inter0), .b(s_286), .O(gate410inter1));
  and2  gate2551(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2552(.a(s_286), .O(gate410inter3));
  inv1  gate2553(.a(s_287), .O(gate410inter4));
  nand2 gate2554(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2555(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2556(.a(G24), .O(gate410inter7));
  inv1  gate2557(.a(G1105), .O(gate410inter8));
  nand2 gate2558(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2559(.a(s_287), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2560(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2561(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2562(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1947(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1948(.a(gate413inter0), .b(s_200), .O(gate413inter1));
  and2  gate1949(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1950(.a(s_200), .O(gate413inter3));
  inv1  gate1951(.a(s_201), .O(gate413inter4));
  nand2 gate1952(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1953(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1954(.a(G27), .O(gate413inter7));
  inv1  gate1955(.a(G1114), .O(gate413inter8));
  nand2 gate1956(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1957(.a(s_201), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1958(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1959(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1960(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate561(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate562(.a(gate414inter0), .b(s_2), .O(gate414inter1));
  and2  gate563(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate564(.a(s_2), .O(gate414inter3));
  inv1  gate565(.a(s_3), .O(gate414inter4));
  nand2 gate566(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate567(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate568(.a(G28), .O(gate414inter7));
  inv1  gate569(.a(G1117), .O(gate414inter8));
  nand2 gate570(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate571(.a(s_3), .b(gate414inter3), .O(gate414inter10));
  nor2  gate572(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate573(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate574(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1779(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1780(.a(gate415inter0), .b(s_176), .O(gate415inter1));
  and2  gate1781(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1782(.a(s_176), .O(gate415inter3));
  inv1  gate1783(.a(s_177), .O(gate415inter4));
  nand2 gate1784(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1785(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1786(.a(G29), .O(gate415inter7));
  inv1  gate1787(.a(G1120), .O(gate415inter8));
  nand2 gate1788(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1789(.a(s_177), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1790(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1791(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1792(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate841(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate842(.a(gate416inter0), .b(s_42), .O(gate416inter1));
  and2  gate843(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate844(.a(s_42), .O(gate416inter3));
  inv1  gate845(.a(s_43), .O(gate416inter4));
  nand2 gate846(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate847(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate848(.a(G30), .O(gate416inter7));
  inv1  gate849(.a(G1123), .O(gate416inter8));
  nand2 gate850(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate851(.a(s_43), .b(gate416inter3), .O(gate416inter10));
  nor2  gate852(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate853(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate854(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1555(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1556(.a(gate420inter0), .b(s_144), .O(gate420inter1));
  and2  gate1557(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1558(.a(s_144), .O(gate420inter3));
  inv1  gate1559(.a(s_145), .O(gate420inter4));
  nand2 gate1560(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1561(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1562(.a(G1036), .O(gate420inter7));
  inv1  gate1563(.a(G1132), .O(gate420inter8));
  nand2 gate1564(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1565(.a(s_145), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1566(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1567(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1568(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1191(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1192(.a(gate423inter0), .b(s_92), .O(gate423inter1));
  and2  gate1193(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1194(.a(s_92), .O(gate423inter3));
  inv1  gate1195(.a(s_93), .O(gate423inter4));
  nand2 gate1196(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1197(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1198(.a(G3), .O(gate423inter7));
  inv1  gate1199(.a(G1138), .O(gate423inter8));
  nand2 gate1200(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1201(.a(s_93), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1202(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1203(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1204(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1961(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1962(.a(gate424inter0), .b(s_202), .O(gate424inter1));
  and2  gate1963(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1964(.a(s_202), .O(gate424inter3));
  inv1  gate1965(.a(s_203), .O(gate424inter4));
  nand2 gate1966(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1967(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1968(.a(G1042), .O(gate424inter7));
  inv1  gate1969(.a(G1138), .O(gate424inter8));
  nand2 gate1970(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1971(.a(s_203), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1972(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1973(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1974(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1261(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1262(.a(gate425inter0), .b(s_102), .O(gate425inter1));
  and2  gate1263(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1264(.a(s_102), .O(gate425inter3));
  inv1  gate1265(.a(s_103), .O(gate425inter4));
  nand2 gate1266(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1267(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1268(.a(G4), .O(gate425inter7));
  inv1  gate1269(.a(G1141), .O(gate425inter8));
  nand2 gate1270(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1271(.a(s_103), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1272(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1273(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1274(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2045(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2046(.a(gate426inter0), .b(s_214), .O(gate426inter1));
  and2  gate2047(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2048(.a(s_214), .O(gate426inter3));
  inv1  gate2049(.a(s_215), .O(gate426inter4));
  nand2 gate2050(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2051(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2052(.a(G1045), .O(gate426inter7));
  inv1  gate2053(.a(G1141), .O(gate426inter8));
  nand2 gate2054(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2055(.a(s_215), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2056(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2057(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2058(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2451(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2452(.a(gate427inter0), .b(s_272), .O(gate427inter1));
  and2  gate2453(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2454(.a(s_272), .O(gate427inter3));
  inv1  gate2455(.a(s_273), .O(gate427inter4));
  nand2 gate2456(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2457(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2458(.a(G5), .O(gate427inter7));
  inv1  gate2459(.a(G1144), .O(gate427inter8));
  nand2 gate2460(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2461(.a(s_273), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2462(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2463(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2464(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2465(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2466(.a(gate429inter0), .b(s_274), .O(gate429inter1));
  and2  gate2467(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2468(.a(s_274), .O(gate429inter3));
  inv1  gate2469(.a(s_275), .O(gate429inter4));
  nand2 gate2470(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2471(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2472(.a(G6), .O(gate429inter7));
  inv1  gate2473(.a(G1147), .O(gate429inter8));
  nand2 gate2474(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2475(.a(s_275), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2476(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2477(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2478(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1611(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1612(.a(gate432inter0), .b(s_152), .O(gate432inter1));
  and2  gate1613(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1614(.a(s_152), .O(gate432inter3));
  inv1  gate1615(.a(s_153), .O(gate432inter4));
  nand2 gate1616(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1617(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1618(.a(G1054), .O(gate432inter7));
  inv1  gate1619(.a(G1150), .O(gate432inter8));
  nand2 gate1620(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1621(.a(s_153), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1622(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1623(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1624(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2577(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2578(.a(gate433inter0), .b(s_290), .O(gate433inter1));
  and2  gate2579(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2580(.a(s_290), .O(gate433inter3));
  inv1  gate2581(.a(s_291), .O(gate433inter4));
  nand2 gate2582(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2583(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2584(.a(G8), .O(gate433inter7));
  inv1  gate2585(.a(G1153), .O(gate433inter8));
  nand2 gate2586(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2587(.a(s_291), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2588(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2589(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2590(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2297(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2298(.a(gate435inter0), .b(s_250), .O(gate435inter1));
  and2  gate2299(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2300(.a(s_250), .O(gate435inter3));
  inv1  gate2301(.a(s_251), .O(gate435inter4));
  nand2 gate2302(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2303(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2304(.a(G9), .O(gate435inter7));
  inv1  gate2305(.a(G1156), .O(gate435inter8));
  nand2 gate2306(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2307(.a(s_251), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2308(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2309(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2310(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate757(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate758(.a(gate437inter0), .b(s_30), .O(gate437inter1));
  and2  gate759(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate760(.a(s_30), .O(gate437inter3));
  inv1  gate761(.a(s_31), .O(gate437inter4));
  nand2 gate762(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate763(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate764(.a(G10), .O(gate437inter7));
  inv1  gate765(.a(G1159), .O(gate437inter8));
  nand2 gate766(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate767(.a(s_31), .b(gate437inter3), .O(gate437inter10));
  nor2  gate768(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate769(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate770(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2339(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2340(.a(gate438inter0), .b(s_256), .O(gate438inter1));
  and2  gate2341(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2342(.a(s_256), .O(gate438inter3));
  inv1  gate2343(.a(s_257), .O(gate438inter4));
  nand2 gate2344(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2345(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2346(.a(G1063), .O(gate438inter7));
  inv1  gate2347(.a(G1159), .O(gate438inter8));
  nand2 gate2348(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2349(.a(s_257), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2350(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2351(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2352(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2759(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2760(.a(gate441inter0), .b(s_316), .O(gate441inter1));
  and2  gate2761(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2762(.a(s_316), .O(gate441inter3));
  inv1  gate2763(.a(s_317), .O(gate441inter4));
  nand2 gate2764(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2765(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2766(.a(G12), .O(gate441inter7));
  inv1  gate2767(.a(G1165), .O(gate441inter8));
  nand2 gate2768(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2769(.a(s_317), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2770(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2771(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2772(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2493(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2494(.a(gate442inter0), .b(s_278), .O(gate442inter1));
  and2  gate2495(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2496(.a(s_278), .O(gate442inter3));
  inv1  gate2497(.a(s_279), .O(gate442inter4));
  nand2 gate2498(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2499(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2500(.a(G1069), .O(gate442inter7));
  inv1  gate2501(.a(G1165), .O(gate442inter8));
  nand2 gate2502(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2503(.a(s_279), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2504(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2505(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2506(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate603(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate604(.a(gate444inter0), .b(s_8), .O(gate444inter1));
  and2  gate605(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate606(.a(s_8), .O(gate444inter3));
  inv1  gate607(.a(s_9), .O(gate444inter4));
  nand2 gate608(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate609(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate610(.a(G1072), .O(gate444inter7));
  inv1  gate611(.a(G1168), .O(gate444inter8));
  nand2 gate612(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate613(.a(s_9), .b(gate444inter3), .O(gate444inter10));
  nor2  gate614(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate615(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate616(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate2633(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2634(.a(gate445inter0), .b(s_298), .O(gate445inter1));
  and2  gate2635(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2636(.a(s_298), .O(gate445inter3));
  inv1  gate2637(.a(s_299), .O(gate445inter4));
  nand2 gate2638(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2639(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2640(.a(G14), .O(gate445inter7));
  inv1  gate2641(.a(G1171), .O(gate445inter8));
  nand2 gate2642(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2643(.a(s_299), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2644(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2645(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2646(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1597(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1598(.a(gate449inter0), .b(s_150), .O(gate449inter1));
  and2  gate1599(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1600(.a(s_150), .O(gate449inter3));
  inv1  gate1601(.a(s_151), .O(gate449inter4));
  nand2 gate1602(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1603(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1604(.a(G16), .O(gate449inter7));
  inv1  gate1605(.a(G1177), .O(gate449inter8));
  nand2 gate1606(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1607(.a(s_151), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1608(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1609(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1610(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate631(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate632(.a(gate450inter0), .b(s_12), .O(gate450inter1));
  and2  gate633(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate634(.a(s_12), .O(gate450inter3));
  inv1  gate635(.a(s_13), .O(gate450inter4));
  nand2 gate636(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate637(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate638(.a(G1081), .O(gate450inter7));
  inv1  gate639(.a(G1177), .O(gate450inter8));
  nand2 gate640(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate641(.a(s_13), .b(gate450inter3), .O(gate450inter10));
  nor2  gate642(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate643(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate644(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1765(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1766(.a(gate454inter0), .b(s_174), .O(gate454inter1));
  and2  gate1767(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1768(.a(s_174), .O(gate454inter3));
  inv1  gate1769(.a(s_175), .O(gate454inter4));
  nand2 gate1770(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1771(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1772(.a(G1087), .O(gate454inter7));
  inv1  gate1773(.a(G1183), .O(gate454inter8));
  nand2 gate1774(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1775(.a(s_175), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1776(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1777(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1778(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1639(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1640(.a(gate456inter0), .b(s_156), .O(gate456inter1));
  and2  gate1641(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1642(.a(s_156), .O(gate456inter3));
  inv1  gate1643(.a(s_157), .O(gate456inter4));
  nand2 gate1644(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1645(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1646(.a(G1090), .O(gate456inter7));
  inv1  gate1647(.a(G1186), .O(gate456inter8));
  nand2 gate1648(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1649(.a(s_157), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1650(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1651(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1652(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2773(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2774(.a(gate459inter0), .b(s_318), .O(gate459inter1));
  and2  gate2775(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2776(.a(s_318), .O(gate459inter3));
  inv1  gate2777(.a(s_319), .O(gate459inter4));
  nand2 gate2778(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2779(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2780(.a(G21), .O(gate459inter7));
  inv1  gate2781(.a(G1192), .O(gate459inter8));
  nand2 gate2782(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2783(.a(s_319), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2784(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2785(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2786(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2395(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2396(.a(gate461inter0), .b(s_264), .O(gate461inter1));
  and2  gate2397(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2398(.a(s_264), .O(gate461inter3));
  inv1  gate2399(.a(s_265), .O(gate461inter4));
  nand2 gate2400(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2401(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2402(.a(G22), .O(gate461inter7));
  inv1  gate2403(.a(G1195), .O(gate461inter8));
  nand2 gate2404(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2405(.a(s_265), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2406(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2407(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2408(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2325(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2326(.a(gate462inter0), .b(s_254), .O(gate462inter1));
  and2  gate2327(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2328(.a(s_254), .O(gate462inter3));
  inv1  gate2329(.a(s_255), .O(gate462inter4));
  nand2 gate2330(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2331(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2332(.a(G1099), .O(gate462inter7));
  inv1  gate2333(.a(G1195), .O(gate462inter8));
  nand2 gate2334(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2335(.a(s_255), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2336(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2337(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2338(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate897(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate898(.a(gate463inter0), .b(s_50), .O(gate463inter1));
  and2  gate899(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate900(.a(s_50), .O(gate463inter3));
  inv1  gate901(.a(s_51), .O(gate463inter4));
  nand2 gate902(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate903(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate904(.a(G23), .O(gate463inter7));
  inv1  gate905(.a(G1198), .O(gate463inter8));
  nand2 gate906(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate907(.a(s_51), .b(gate463inter3), .O(gate463inter10));
  nor2  gate908(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate909(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate910(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1107(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1108(.a(gate464inter0), .b(s_80), .O(gate464inter1));
  and2  gate1109(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1110(.a(s_80), .O(gate464inter3));
  inv1  gate1111(.a(s_81), .O(gate464inter4));
  nand2 gate1112(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1113(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1114(.a(G1102), .O(gate464inter7));
  inv1  gate1115(.a(G1198), .O(gate464inter8));
  nand2 gate1116(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1117(.a(s_81), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1118(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1119(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1120(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2059(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2060(.a(gate466inter0), .b(s_216), .O(gate466inter1));
  and2  gate2061(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2062(.a(s_216), .O(gate466inter3));
  inv1  gate2063(.a(s_217), .O(gate466inter4));
  nand2 gate2064(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2065(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2066(.a(G1105), .O(gate466inter7));
  inv1  gate2067(.a(G1201), .O(gate466inter8));
  nand2 gate2068(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2069(.a(s_217), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2070(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2071(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2072(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1541(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1542(.a(gate470inter0), .b(s_142), .O(gate470inter1));
  and2  gate1543(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1544(.a(s_142), .O(gate470inter3));
  inv1  gate1545(.a(s_143), .O(gate470inter4));
  nand2 gate1546(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1547(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1548(.a(G1111), .O(gate470inter7));
  inv1  gate1549(.a(G1207), .O(gate470inter8));
  nand2 gate1550(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1551(.a(s_143), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1552(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1553(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1554(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2703(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2704(.a(gate471inter0), .b(s_308), .O(gate471inter1));
  and2  gate2705(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2706(.a(s_308), .O(gate471inter3));
  inv1  gate2707(.a(s_309), .O(gate471inter4));
  nand2 gate2708(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2709(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2710(.a(G27), .O(gate471inter7));
  inv1  gate2711(.a(G1210), .O(gate471inter8));
  nand2 gate2712(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2713(.a(s_309), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2714(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2715(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2716(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1065(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1066(.a(gate472inter0), .b(s_74), .O(gate472inter1));
  and2  gate1067(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1068(.a(s_74), .O(gate472inter3));
  inv1  gate1069(.a(s_75), .O(gate472inter4));
  nand2 gate1070(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1071(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1072(.a(G1114), .O(gate472inter7));
  inv1  gate1073(.a(G1210), .O(gate472inter8));
  nand2 gate1074(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1075(.a(s_75), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1076(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1077(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1078(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2801(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2802(.a(gate478inter0), .b(s_322), .O(gate478inter1));
  and2  gate2803(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2804(.a(s_322), .O(gate478inter3));
  inv1  gate2805(.a(s_323), .O(gate478inter4));
  nand2 gate2806(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2807(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2808(.a(G1123), .O(gate478inter7));
  inv1  gate2809(.a(G1219), .O(gate478inter8));
  nand2 gate2810(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2811(.a(s_323), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2812(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2813(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2814(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1317(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1318(.a(gate481inter0), .b(s_110), .O(gate481inter1));
  and2  gate1319(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1320(.a(s_110), .O(gate481inter3));
  inv1  gate1321(.a(s_111), .O(gate481inter4));
  nand2 gate1322(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1323(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1324(.a(G32), .O(gate481inter7));
  inv1  gate1325(.a(G1225), .O(gate481inter8));
  nand2 gate1326(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1327(.a(s_111), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1328(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1329(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1330(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1037(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1038(.a(gate486inter0), .b(s_70), .O(gate486inter1));
  and2  gate1039(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1040(.a(s_70), .O(gate486inter3));
  inv1  gate1041(.a(s_71), .O(gate486inter4));
  nand2 gate1042(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1043(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1044(.a(G1234), .O(gate486inter7));
  inv1  gate1045(.a(G1235), .O(gate486inter8));
  nand2 gate1046(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1047(.a(s_71), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1048(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1049(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1050(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2171(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2172(.a(gate489inter0), .b(s_232), .O(gate489inter1));
  and2  gate2173(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2174(.a(s_232), .O(gate489inter3));
  inv1  gate2175(.a(s_233), .O(gate489inter4));
  nand2 gate2176(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2177(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2178(.a(G1240), .O(gate489inter7));
  inv1  gate2179(.a(G1241), .O(gate489inter8));
  nand2 gate2180(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2181(.a(s_233), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2182(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2183(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2184(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2157(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2158(.a(gate491inter0), .b(s_230), .O(gate491inter1));
  and2  gate2159(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2160(.a(s_230), .O(gate491inter3));
  inv1  gate2161(.a(s_231), .O(gate491inter4));
  nand2 gate2162(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2163(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2164(.a(G1244), .O(gate491inter7));
  inv1  gate2165(.a(G1245), .O(gate491inter8));
  nand2 gate2166(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2167(.a(s_231), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2168(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2169(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2170(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate869(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate870(.a(gate492inter0), .b(s_46), .O(gate492inter1));
  and2  gate871(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate872(.a(s_46), .O(gate492inter3));
  inv1  gate873(.a(s_47), .O(gate492inter4));
  nand2 gate874(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate875(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate876(.a(G1246), .O(gate492inter7));
  inv1  gate877(.a(G1247), .O(gate492inter8));
  nand2 gate878(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate879(.a(s_47), .b(gate492inter3), .O(gate492inter10));
  nor2  gate880(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate881(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate882(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1079(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1080(.a(gate493inter0), .b(s_76), .O(gate493inter1));
  and2  gate1081(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1082(.a(s_76), .O(gate493inter3));
  inv1  gate1083(.a(s_77), .O(gate493inter4));
  nand2 gate1084(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1085(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1086(.a(G1248), .O(gate493inter7));
  inv1  gate1087(.a(G1249), .O(gate493inter8));
  nand2 gate1088(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1089(.a(s_77), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1090(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1091(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1092(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate855(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate856(.a(gate495inter0), .b(s_44), .O(gate495inter1));
  and2  gate857(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate858(.a(s_44), .O(gate495inter3));
  inv1  gate859(.a(s_45), .O(gate495inter4));
  nand2 gate860(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate861(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate862(.a(G1252), .O(gate495inter7));
  inv1  gate863(.a(G1253), .O(gate495inter8));
  nand2 gate864(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate865(.a(s_45), .b(gate495inter3), .O(gate495inter10));
  nor2  gate866(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate867(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate868(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2787(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2788(.a(gate499inter0), .b(s_320), .O(gate499inter1));
  and2  gate2789(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2790(.a(s_320), .O(gate499inter3));
  inv1  gate2791(.a(s_321), .O(gate499inter4));
  nand2 gate2792(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2793(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2794(.a(G1260), .O(gate499inter7));
  inv1  gate2795(.a(G1261), .O(gate499inter8));
  nand2 gate2796(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2797(.a(s_321), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2798(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2799(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2800(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1653(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1654(.a(gate501inter0), .b(s_158), .O(gate501inter1));
  and2  gate1655(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1656(.a(s_158), .O(gate501inter3));
  inv1  gate1657(.a(s_159), .O(gate501inter4));
  nand2 gate1658(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1659(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1660(.a(G1264), .O(gate501inter7));
  inv1  gate1661(.a(G1265), .O(gate501inter8));
  nand2 gate1662(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1663(.a(s_159), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1664(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1665(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1666(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule