module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate939(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate940(.a(gate15inter0), .b(s_56), .O(gate15inter1));
  and2  gate941(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate942(.a(s_56), .O(gate15inter3));
  inv1  gate943(.a(s_57), .O(gate15inter4));
  nand2 gate944(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate945(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate946(.a(G13), .O(gate15inter7));
  inv1  gate947(.a(G14), .O(gate15inter8));
  nand2 gate948(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate949(.a(s_57), .b(gate15inter3), .O(gate15inter10));
  nor2  gate950(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate951(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate952(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate771(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate772(.a(gate17inter0), .b(s_32), .O(gate17inter1));
  and2  gate773(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate774(.a(s_32), .O(gate17inter3));
  inv1  gate775(.a(s_33), .O(gate17inter4));
  nand2 gate776(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate777(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate778(.a(G17), .O(gate17inter7));
  inv1  gate779(.a(G18), .O(gate17inter8));
  nand2 gate780(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate781(.a(s_33), .b(gate17inter3), .O(gate17inter10));
  nor2  gate782(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate783(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate784(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate645(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate646(.a(gate24inter0), .b(s_14), .O(gate24inter1));
  and2  gate647(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate648(.a(s_14), .O(gate24inter3));
  inv1  gate649(.a(s_15), .O(gate24inter4));
  nand2 gate650(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate651(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate652(.a(G31), .O(gate24inter7));
  inv1  gate653(.a(G32), .O(gate24inter8));
  nand2 gate654(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate655(.a(s_15), .b(gate24inter3), .O(gate24inter10));
  nor2  gate656(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate657(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate658(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1485(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1486(.a(gate27inter0), .b(s_134), .O(gate27inter1));
  and2  gate1487(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1488(.a(s_134), .O(gate27inter3));
  inv1  gate1489(.a(s_135), .O(gate27inter4));
  nand2 gate1490(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1491(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1492(.a(G2), .O(gate27inter7));
  inv1  gate1493(.a(G6), .O(gate27inter8));
  nand2 gate1494(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1495(.a(s_135), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1496(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1497(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1498(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1625(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1626(.a(gate34inter0), .b(s_154), .O(gate34inter1));
  and2  gate1627(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1628(.a(s_154), .O(gate34inter3));
  inv1  gate1629(.a(s_155), .O(gate34inter4));
  nand2 gate1630(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1631(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1632(.a(G25), .O(gate34inter7));
  inv1  gate1633(.a(G29), .O(gate34inter8));
  nand2 gate1634(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1635(.a(s_155), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1636(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1637(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1638(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1919(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1920(.a(gate36inter0), .b(s_196), .O(gate36inter1));
  and2  gate1921(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1922(.a(s_196), .O(gate36inter3));
  inv1  gate1923(.a(s_197), .O(gate36inter4));
  nand2 gate1924(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1925(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1926(.a(G26), .O(gate36inter7));
  inv1  gate1927(.a(G30), .O(gate36inter8));
  nand2 gate1928(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1929(.a(s_197), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1930(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1931(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1932(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate911(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate912(.a(gate37inter0), .b(s_52), .O(gate37inter1));
  and2  gate913(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate914(.a(s_52), .O(gate37inter3));
  inv1  gate915(.a(s_53), .O(gate37inter4));
  nand2 gate916(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate917(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate918(.a(G19), .O(gate37inter7));
  inv1  gate919(.a(G23), .O(gate37inter8));
  nand2 gate920(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate921(.a(s_53), .b(gate37inter3), .O(gate37inter10));
  nor2  gate922(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate923(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate924(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1121(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1122(.a(gate41inter0), .b(s_82), .O(gate41inter1));
  and2  gate1123(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1124(.a(s_82), .O(gate41inter3));
  inv1  gate1125(.a(s_83), .O(gate41inter4));
  nand2 gate1126(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1127(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1128(.a(G1), .O(gate41inter7));
  inv1  gate1129(.a(G266), .O(gate41inter8));
  nand2 gate1130(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1131(.a(s_83), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1132(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1133(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1134(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1009(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1010(.a(gate42inter0), .b(s_66), .O(gate42inter1));
  and2  gate1011(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1012(.a(s_66), .O(gate42inter3));
  inv1  gate1013(.a(s_67), .O(gate42inter4));
  nand2 gate1014(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1015(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1016(.a(G2), .O(gate42inter7));
  inv1  gate1017(.a(G266), .O(gate42inter8));
  nand2 gate1018(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1019(.a(s_67), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1020(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1021(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1022(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate729(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate730(.a(gate57inter0), .b(s_26), .O(gate57inter1));
  and2  gate731(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate732(.a(s_26), .O(gate57inter3));
  inv1  gate733(.a(s_27), .O(gate57inter4));
  nand2 gate734(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate735(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate736(.a(G17), .O(gate57inter7));
  inv1  gate737(.a(G290), .O(gate57inter8));
  nand2 gate738(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate739(.a(s_27), .b(gate57inter3), .O(gate57inter10));
  nor2  gate740(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate741(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate742(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1541(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1542(.a(gate61inter0), .b(s_142), .O(gate61inter1));
  and2  gate1543(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1544(.a(s_142), .O(gate61inter3));
  inv1  gate1545(.a(s_143), .O(gate61inter4));
  nand2 gate1546(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1547(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1548(.a(G21), .O(gate61inter7));
  inv1  gate1549(.a(G296), .O(gate61inter8));
  nand2 gate1550(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1551(.a(s_143), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1552(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1553(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1554(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1093(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1094(.a(gate65inter0), .b(s_78), .O(gate65inter1));
  and2  gate1095(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1096(.a(s_78), .O(gate65inter3));
  inv1  gate1097(.a(s_79), .O(gate65inter4));
  nand2 gate1098(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1099(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1100(.a(G25), .O(gate65inter7));
  inv1  gate1101(.a(G302), .O(gate65inter8));
  nand2 gate1102(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1103(.a(s_79), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1104(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1105(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1106(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1877(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1878(.a(gate67inter0), .b(s_190), .O(gate67inter1));
  and2  gate1879(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1880(.a(s_190), .O(gate67inter3));
  inv1  gate1881(.a(s_191), .O(gate67inter4));
  nand2 gate1882(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1883(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1884(.a(G27), .O(gate67inter7));
  inv1  gate1885(.a(G305), .O(gate67inter8));
  nand2 gate1886(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1887(.a(s_191), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1888(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1889(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1890(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1527(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1528(.a(gate68inter0), .b(s_140), .O(gate68inter1));
  and2  gate1529(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1530(.a(s_140), .O(gate68inter3));
  inv1  gate1531(.a(s_141), .O(gate68inter4));
  nand2 gate1532(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1533(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1534(.a(G28), .O(gate68inter7));
  inv1  gate1535(.a(G305), .O(gate68inter8));
  nand2 gate1536(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1537(.a(s_141), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1538(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1539(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1540(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1023(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1024(.a(gate75inter0), .b(s_68), .O(gate75inter1));
  and2  gate1025(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1026(.a(s_68), .O(gate75inter3));
  inv1  gate1027(.a(s_69), .O(gate75inter4));
  nand2 gate1028(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1029(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1030(.a(G9), .O(gate75inter7));
  inv1  gate1031(.a(G317), .O(gate75inter8));
  nand2 gate1032(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1033(.a(s_69), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1034(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1035(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1036(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate855(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate856(.a(gate78inter0), .b(s_44), .O(gate78inter1));
  and2  gate857(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate858(.a(s_44), .O(gate78inter3));
  inv1  gate859(.a(s_45), .O(gate78inter4));
  nand2 gate860(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate861(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate862(.a(G6), .O(gate78inter7));
  inv1  gate863(.a(G320), .O(gate78inter8));
  nand2 gate864(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate865(.a(s_45), .b(gate78inter3), .O(gate78inter10));
  nor2  gate866(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate867(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate868(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1807(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1808(.a(gate80inter0), .b(s_180), .O(gate80inter1));
  and2  gate1809(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1810(.a(s_180), .O(gate80inter3));
  inv1  gate1811(.a(s_181), .O(gate80inter4));
  nand2 gate1812(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1813(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1814(.a(G14), .O(gate80inter7));
  inv1  gate1815(.a(G323), .O(gate80inter8));
  nand2 gate1816(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1817(.a(s_181), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1818(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1819(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1820(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1723(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1724(.a(gate83inter0), .b(s_168), .O(gate83inter1));
  and2  gate1725(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1726(.a(s_168), .O(gate83inter3));
  inv1  gate1727(.a(s_169), .O(gate83inter4));
  nand2 gate1728(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1729(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1730(.a(G11), .O(gate83inter7));
  inv1  gate1731(.a(G329), .O(gate83inter8));
  nand2 gate1732(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1733(.a(s_169), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1734(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1735(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1736(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate575(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate576(.a(gate88inter0), .b(s_4), .O(gate88inter1));
  and2  gate577(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate578(.a(s_4), .O(gate88inter3));
  inv1  gate579(.a(s_5), .O(gate88inter4));
  nand2 gate580(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate581(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate582(.a(G16), .O(gate88inter7));
  inv1  gate583(.a(G335), .O(gate88inter8));
  nand2 gate584(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate585(.a(s_5), .b(gate88inter3), .O(gate88inter10));
  nor2  gate586(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate587(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate588(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate953(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate954(.a(gate106inter0), .b(s_58), .O(gate106inter1));
  and2  gate955(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate956(.a(s_58), .O(gate106inter3));
  inv1  gate957(.a(s_59), .O(gate106inter4));
  nand2 gate958(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate959(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate960(.a(G364), .O(gate106inter7));
  inv1  gate961(.a(G365), .O(gate106inter8));
  nand2 gate962(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate963(.a(s_59), .b(gate106inter3), .O(gate106inter10));
  nor2  gate964(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate965(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate966(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1737(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1738(.a(gate107inter0), .b(s_170), .O(gate107inter1));
  and2  gate1739(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1740(.a(s_170), .O(gate107inter3));
  inv1  gate1741(.a(s_171), .O(gate107inter4));
  nand2 gate1742(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1743(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1744(.a(G366), .O(gate107inter7));
  inv1  gate1745(.a(G367), .O(gate107inter8));
  nand2 gate1746(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1747(.a(s_171), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1748(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1749(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1750(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1863(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1864(.a(gate110inter0), .b(s_188), .O(gate110inter1));
  and2  gate1865(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1866(.a(s_188), .O(gate110inter3));
  inv1  gate1867(.a(s_189), .O(gate110inter4));
  nand2 gate1868(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1869(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1870(.a(G372), .O(gate110inter7));
  inv1  gate1871(.a(G373), .O(gate110inter8));
  nand2 gate1872(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1873(.a(s_189), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1874(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1875(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1876(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate561(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate562(.a(gate115inter0), .b(s_2), .O(gate115inter1));
  and2  gate563(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate564(.a(s_2), .O(gate115inter3));
  inv1  gate565(.a(s_3), .O(gate115inter4));
  nand2 gate566(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate567(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate568(.a(G382), .O(gate115inter7));
  inv1  gate569(.a(G383), .O(gate115inter8));
  nand2 gate570(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate571(.a(s_3), .b(gate115inter3), .O(gate115inter10));
  nor2  gate572(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate573(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate574(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate813(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate814(.a(gate117inter0), .b(s_38), .O(gate117inter1));
  and2  gate815(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate816(.a(s_38), .O(gate117inter3));
  inv1  gate817(.a(s_39), .O(gate117inter4));
  nand2 gate818(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate819(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate820(.a(G386), .O(gate117inter7));
  inv1  gate821(.a(G387), .O(gate117inter8));
  nand2 gate822(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate823(.a(s_39), .b(gate117inter3), .O(gate117inter10));
  nor2  gate824(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate825(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate826(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate701(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate702(.a(gate119inter0), .b(s_22), .O(gate119inter1));
  and2  gate703(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate704(.a(s_22), .O(gate119inter3));
  inv1  gate705(.a(s_23), .O(gate119inter4));
  nand2 gate706(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate707(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate708(.a(G390), .O(gate119inter7));
  inv1  gate709(.a(G391), .O(gate119inter8));
  nand2 gate710(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate711(.a(s_23), .b(gate119inter3), .O(gate119inter10));
  nor2  gate712(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate713(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate714(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate743(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate744(.a(gate124inter0), .b(s_28), .O(gate124inter1));
  and2  gate745(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate746(.a(s_28), .O(gate124inter3));
  inv1  gate747(.a(s_29), .O(gate124inter4));
  nand2 gate748(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate749(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate750(.a(G400), .O(gate124inter7));
  inv1  gate751(.a(G401), .O(gate124inter8));
  nand2 gate752(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate753(.a(s_29), .b(gate124inter3), .O(gate124inter10));
  nor2  gate754(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate755(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate756(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1947(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1948(.a(gate134inter0), .b(s_200), .O(gate134inter1));
  and2  gate1949(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1950(.a(s_200), .O(gate134inter3));
  inv1  gate1951(.a(s_201), .O(gate134inter4));
  nand2 gate1952(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1953(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1954(.a(G420), .O(gate134inter7));
  inv1  gate1955(.a(G421), .O(gate134inter8));
  nand2 gate1956(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1957(.a(s_201), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1958(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1959(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1960(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate715(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate716(.a(gate138inter0), .b(s_24), .O(gate138inter1));
  and2  gate717(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate718(.a(s_24), .O(gate138inter3));
  inv1  gate719(.a(s_25), .O(gate138inter4));
  nand2 gate720(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate721(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate722(.a(G432), .O(gate138inter7));
  inv1  gate723(.a(G435), .O(gate138inter8));
  nand2 gate724(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate725(.a(s_25), .b(gate138inter3), .O(gate138inter10));
  nor2  gate726(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate727(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate728(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1135(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1136(.a(gate141inter0), .b(s_84), .O(gate141inter1));
  and2  gate1137(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1138(.a(s_84), .O(gate141inter3));
  inv1  gate1139(.a(s_85), .O(gate141inter4));
  nand2 gate1140(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1141(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1142(.a(G450), .O(gate141inter7));
  inv1  gate1143(.a(G453), .O(gate141inter8));
  nand2 gate1144(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1145(.a(s_85), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1146(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1147(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1148(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate841(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate842(.a(gate142inter0), .b(s_42), .O(gate142inter1));
  and2  gate843(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate844(.a(s_42), .O(gate142inter3));
  inv1  gate845(.a(s_43), .O(gate142inter4));
  nand2 gate846(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate847(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate848(.a(G456), .O(gate142inter7));
  inv1  gate849(.a(G459), .O(gate142inter8));
  nand2 gate850(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate851(.a(s_43), .b(gate142inter3), .O(gate142inter10));
  nor2  gate852(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate853(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate854(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1219(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1220(.a(gate144inter0), .b(s_96), .O(gate144inter1));
  and2  gate1221(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1222(.a(s_96), .O(gate144inter3));
  inv1  gate1223(.a(s_97), .O(gate144inter4));
  nand2 gate1224(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1225(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1226(.a(G468), .O(gate144inter7));
  inv1  gate1227(.a(G471), .O(gate144inter8));
  nand2 gate1228(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1229(.a(s_97), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1230(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1231(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1232(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate981(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate982(.a(gate150inter0), .b(s_62), .O(gate150inter1));
  and2  gate983(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate984(.a(s_62), .O(gate150inter3));
  inv1  gate985(.a(s_63), .O(gate150inter4));
  nand2 gate986(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate987(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate988(.a(G504), .O(gate150inter7));
  inv1  gate989(.a(G507), .O(gate150inter8));
  nand2 gate990(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate991(.a(s_63), .b(gate150inter3), .O(gate150inter10));
  nor2  gate992(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate993(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate994(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1359(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1360(.a(gate153inter0), .b(s_116), .O(gate153inter1));
  and2  gate1361(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1362(.a(s_116), .O(gate153inter3));
  inv1  gate1363(.a(s_117), .O(gate153inter4));
  nand2 gate1364(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1365(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1366(.a(G426), .O(gate153inter7));
  inv1  gate1367(.a(G522), .O(gate153inter8));
  nand2 gate1368(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1369(.a(s_117), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1370(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1371(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1372(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1429(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1430(.a(gate155inter0), .b(s_126), .O(gate155inter1));
  and2  gate1431(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1432(.a(s_126), .O(gate155inter3));
  inv1  gate1433(.a(s_127), .O(gate155inter4));
  nand2 gate1434(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1435(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1436(.a(G432), .O(gate155inter7));
  inv1  gate1437(.a(G525), .O(gate155inter8));
  nand2 gate1438(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1439(.a(s_127), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1440(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1441(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1442(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1849(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1850(.a(gate156inter0), .b(s_186), .O(gate156inter1));
  and2  gate1851(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1852(.a(s_186), .O(gate156inter3));
  inv1  gate1853(.a(s_187), .O(gate156inter4));
  nand2 gate1854(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1855(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1856(.a(G435), .O(gate156inter7));
  inv1  gate1857(.a(G525), .O(gate156inter8));
  nand2 gate1858(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1859(.a(s_187), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1860(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1861(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1862(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate757(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate758(.a(gate159inter0), .b(s_30), .O(gate159inter1));
  and2  gate759(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate760(.a(s_30), .O(gate159inter3));
  inv1  gate761(.a(s_31), .O(gate159inter4));
  nand2 gate762(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate763(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate764(.a(G444), .O(gate159inter7));
  inv1  gate765(.a(G531), .O(gate159inter8));
  nand2 gate766(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate767(.a(s_31), .b(gate159inter3), .O(gate159inter10));
  nor2  gate768(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate769(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate770(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1709(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1710(.a(gate160inter0), .b(s_166), .O(gate160inter1));
  and2  gate1711(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1712(.a(s_166), .O(gate160inter3));
  inv1  gate1713(.a(s_167), .O(gate160inter4));
  nand2 gate1714(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1715(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1716(.a(G447), .O(gate160inter7));
  inv1  gate1717(.a(G531), .O(gate160inter8));
  nand2 gate1718(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1719(.a(s_167), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1720(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1721(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1722(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1443(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1444(.a(gate163inter0), .b(s_128), .O(gate163inter1));
  and2  gate1445(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1446(.a(s_128), .O(gate163inter3));
  inv1  gate1447(.a(s_129), .O(gate163inter4));
  nand2 gate1448(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1449(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1450(.a(G456), .O(gate163inter7));
  inv1  gate1451(.a(G537), .O(gate163inter8));
  nand2 gate1452(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1453(.a(s_129), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1454(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1455(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1456(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1835(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1836(.a(gate165inter0), .b(s_184), .O(gate165inter1));
  and2  gate1837(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1838(.a(s_184), .O(gate165inter3));
  inv1  gate1839(.a(s_185), .O(gate165inter4));
  nand2 gate1840(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1841(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1842(.a(G462), .O(gate165inter7));
  inv1  gate1843(.a(G540), .O(gate165inter8));
  nand2 gate1844(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1845(.a(s_185), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1846(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1847(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1848(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1891(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1892(.a(gate172inter0), .b(s_192), .O(gate172inter1));
  and2  gate1893(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1894(.a(s_192), .O(gate172inter3));
  inv1  gate1895(.a(s_193), .O(gate172inter4));
  nand2 gate1896(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1897(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1898(.a(G483), .O(gate172inter7));
  inv1  gate1899(.a(G549), .O(gate172inter8));
  nand2 gate1900(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1901(.a(s_193), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1902(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1903(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1904(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1611(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1612(.a(gate176inter0), .b(s_152), .O(gate176inter1));
  and2  gate1613(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1614(.a(s_152), .O(gate176inter3));
  inv1  gate1615(.a(s_153), .O(gate176inter4));
  nand2 gate1616(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1617(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1618(.a(G495), .O(gate176inter7));
  inv1  gate1619(.a(G555), .O(gate176inter8));
  nand2 gate1620(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1621(.a(s_153), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1622(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1623(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1624(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1499(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1500(.a(gate179inter0), .b(s_136), .O(gate179inter1));
  and2  gate1501(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1502(.a(s_136), .O(gate179inter3));
  inv1  gate1503(.a(s_137), .O(gate179inter4));
  nand2 gate1504(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1505(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1506(.a(G504), .O(gate179inter7));
  inv1  gate1507(.a(G561), .O(gate179inter8));
  nand2 gate1508(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1509(.a(s_137), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1510(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1511(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1512(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate659(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate660(.a(gate189inter0), .b(s_16), .O(gate189inter1));
  and2  gate661(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate662(.a(s_16), .O(gate189inter3));
  inv1  gate663(.a(s_17), .O(gate189inter4));
  nand2 gate664(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate665(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate666(.a(G578), .O(gate189inter7));
  inv1  gate667(.a(G579), .O(gate189inter8));
  nand2 gate668(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate669(.a(s_17), .b(gate189inter3), .O(gate189inter10));
  nor2  gate670(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate671(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate672(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1177(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1178(.a(gate192inter0), .b(s_90), .O(gate192inter1));
  and2  gate1179(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1180(.a(s_90), .O(gate192inter3));
  inv1  gate1181(.a(s_91), .O(gate192inter4));
  nand2 gate1182(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1183(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1184(.a(G584), .O(gate192inter7));
  inv1  gate1185(.a(G585), .O(gate192inter8));
  nand2 gate1186(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1187(.a(s_91), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1188(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1189(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1190(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate897(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate898(.a(gate195inter0), .b(s_50), .O(gate195inter1));
  and2  gate899(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate900(.a(s_50), .O(gate195inter3));
  inv1  gate901(.a(s_51), .O(gate195inter4));
  nand2 gate902(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate903(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate904(.a(G590), .O(gate195inter7));
  inv1  gate905(.a(G591), .O(gate195inter8));
  nand2 gate906(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate907(.a(s_51), .b(gate195inter3), .O(gate195inter10));
  nor2  gate908(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate909(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate910(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1107(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1108(.a(gate196inter0), .b(s_80), .O(gate196inter1));
  and2  gate1109(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1110(.a(s_80), .O(gate196inter3));
  inv1  gate1111(.a(s_81), .O(gate196inter4));
  nand2 gate1112(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1113(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1114(.a(G592), .O(gate196inter7));
  inv1  gate1115(.a(G593), .O(gate196inter8));
  nand2 gate1116(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1117(.a(s_81), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1118(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1119(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1120(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1779(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1780(.a(gate197inter0), .b(s_176), .O(gate197inter1));
  and2  gate1781(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1782(.a(s_176), .O(gate197inter3));
  inv1  gate1783(.a(s_177), .O(gate197inter4));
  nand2 gate1784(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1785(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1786(.a(G594), .O(gate197inter7));
  inv1  gate1787(.a(G595), .O(gate197inter8));
  nand2 gate1788(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1789(.a(s_177), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1790(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1791(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1792(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1079(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1080(.a(gate203inter0), .b(s_76), .O(gate203inter1));
  and2  gate1081(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1082(.a(s_76), .O(gate203inter3));
  inv1  gate1083(.a(s_77), .O(gate203inter4));
  nand2 gate1084(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1085(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1086(.a(G602), .O(gate203inter7));
  inv1  gate1087(.a(G612), .O(gate203inter8));
  nand2 gate1088(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1089(.a(s_77), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1090(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1091(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1092(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1261(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1262(.a(gate204inter0), .b(s_102), .O(gate204inter1));
  and2  gate1263(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1264(.a(s_102), .O(gate204inter3));
  inv1  gate1265(.a(s_103), .O(gate204inter4));
  nand2 gate1266(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1267(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1268(.a(G607), .O(gate204inter7));
  inv1  gate1269(.a(G617), .O(gate204inter8));
  nand2 gate1270(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1271(.a(s_103), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1272(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1273(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1274(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate995(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate996(.a(gate214inter0), .b(s_64), .O(gate214inter1));
  and2  gate997(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate998(.a(s_64), .O(gate214inter3));
  inv1  gate999(.a(s_65), .O(gate214inter4));
  nand2 gate1000(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1001(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1002(.a(G612), .O(gate214inter7));
  inv1  gate1003(.a(G672), .O(gate214inter8));
  nand2 gate1004(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1005(.a(s_65), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1006(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1007(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1008(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate617(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate618(.a(gate216inter0), .b(s_10), .O(gate216inter1));
  and2  gate619(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate620(.a(s_10), .O(gate216inter3));
  inv1  gate621(.a(s_11), .O(gate216inter4));
  nand2 gate622(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate623(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate624(.a(G617), .O(gate216inter7));
  inv1  gate625(.a(G675), .O(gate216inter8));
  nand2 gate626(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate627(.a(s_11), .b(gate216inter3), .O(gate216inter10));
  nor2  gate628(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate629(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate630(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1163(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1164(.a(gate220inter0), .b(s_88), .O(gate220inter1));
  and2  gate1165(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1166(.a(s_88), .O(gate220inter3));
  inv1  gate1167(.a(s_89), .O(gate220inter4));
  nand2 gate1168(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1169(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1170(.a(G637), .O(gate220inter7));
  inv1  gate1171(.a(G681), .O(gate220inter8));
  nand2 gate1172(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1173(.a(s_89), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1174(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1175(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1176(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1471(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1472(.a(gate223inter0), .b(s_132), .O(gate223inter1));
  and2  gate1473(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1474(.a(s_132), .O(gate223inter3));
  inv1  gate1475(.a(s_133), .O(gate223inter4));
  nand2 gate1476(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1477(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1478(.a(G627), .O(gate223inter7));
  inv1  gate1479(.a(G687), .O(gate223inter8));
  nand2 gate1480(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1481(.a(s_133), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1482(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1483(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1484(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1149(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1150(.a(gate235inter0), .b(s_86), .O(gate235inter1));
  and2  gate1151(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1152(.a(s_86), .O(gate235inter3));
  inv1  gate1153(.a(s_87), .O(gate235inter4));
  nand2 gate1154(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1155(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1156(.a(G248), .O(gate235inter7));
  inv1  gate1157(.a(G724), .O(gate235inter8));
  nand2 gate1158(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1159(.a(s_87), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1160(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1161(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1162(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate1569(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1570(.a(gate236inter0), .b(s_146), .O(gate236inter1));
  and2  gate1571(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1572(.a(s_146), .O(gate236inter3));
  inv1  gate1573(.a(s_147), .O(gate236inter4));
  nand2 gate1574(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1575(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1576(.a(G251), .O(gate236inter7));
  inv1  gate1577(.a(G727), .O(gate236inter8));
  nand2 gate1578(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1579(.a(s_147), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1580(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1581(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1582(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1513(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1514(.a(gate241inter0), .b(s_138), .O(gate241inter1));
  and2  gate1515(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1516(.a(s_138), .O(gate241inter3));
  inv1  gate1517(.a(s_139), .O(gate241inter4));
  nand2 gate1518(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1519(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1520(.a(G242), .O(gate241inter7));
  inv1  gate1521(.a(G730), .O(gate241inter8));
  nand2 gate1522(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1523(.a(s_139), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1524(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1525(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1526(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1317(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1318(.a(gate245inter0), .b(s_110), .O(gate245inter1));
  and2  gate1319(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1320(.a(s_110), .O(gate245inter3));
  inv1  gate1321(.a(s_111), .O(gate245inter4));
  nand2 gate1322(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1323(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1324(.a(G248), .O(gate245inter7));
  inv1  gate1325(.a(G736), .O(gate245inter8));
  nand2 gate1326(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1327(.a(s_111), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1328(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1329(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1330(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1653(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1654(.a(gate248inter0), .b(s_158), .O(gate248inter1));
  and2  gate1655(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1656(.a(s_158), .O(gate248inter3));
  inv1  gate1657(.a(s_159), .O(gate248inter4));
  nand2 gate1658(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1659(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1660(.a(G727), .O(gate248inter7));
  inv1  gate1661(.a(G739), .O(gate248inter8));
  nand2 gate1662(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1663(.a(s_159), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1664(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1665(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1666(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate547(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate548(.a(gate257inter0), .b(s_0), .O(gate257inter1));
  and2  gate549(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate550(.a(s_0), .O(gate257inter3));
  inv1  gate551(.a(s_1), .O(gate257inter4));
  nand2 gate552(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate553(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate554(.a(G754), .O(gate257inter7));
  inv1  gate555(.a(G755), .O(gate257inter8));
  nand2 gate556(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate557(.a(s_1), .b(gate257inter3), .O(gate257inter10));
  nor2  gate558(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate559(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate560(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1191(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1192(.a(gate261inter0), .b(s_92), .O(gate261inter1));
  and2  gate1193(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1194(.a(s_92), .O(gate261inter3));
  inv1  gate1195(.a(s_93), .O(gate261inter4));
  nand2 gate1196(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1197(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1198(.a(G762), .O(gate261inter7));
  inv1  gate1199(.a(G763), .O(gate261inter8));
  nand2 gate1200(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1201(.a(s_93), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1202(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1203(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1204(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1583(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1584(.a(gate262inter0), .b(s_148), .O(gate262inter1));
  and2  gate1585(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1586(.a(s_148), .O(gate262inter3));
  inv1  gate1587(.a(s_149), .O(gate262inter4));
  nand2 gate1588(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1589(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1590(.a(G764), .O(gate262inter7));
  inv1  gate1591(.a(G765), .O(gate262inter8));
  nand2 gate1592(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1593(.a(s_149), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1594(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1595(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1596(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1275(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1276(.a(gate265inter0), .b(s_104), .O(gate265inter1));
  and2  gate1277(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1278(.a(s_104), .O(gate265inter3));
  inv1  gate1279(.a(s_105), .O(gate265inter4));
  nand2 gate1280(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1281(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1282(.a(G642), .O(gate265inter7));
  inv1  gate1283(.a(G770), .O(gate265inter8));
  nand2 gate1284(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1285(.a(s_105), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1286(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1287(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1288(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1331(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1332(.a(gate268inter0), .b(s_112), .O(gate268inter1));
  and2  gate1333(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1334(.a(s_112), .O(gate268inter3));
  inv1  gate1335(.a(s_113), .O(gate268inter4));
  nand2 gate1336(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1337(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1338(.a(G651), .O(gate268inter7));
  inv1  gate1339(.a(G779), .O(gate268inter8));
  nand2 gate1340(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1341(.a(s_113), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1342(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1343(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1344(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1667(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1668(.a(gate270inter0), .b(s_160), .O(gate270inter1));
  and2  gate1669(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1670(.a(s_160), .O(gate270inter3));
  inv1  gate1671(.a(s_161), .O(gate270inter4));
  nand2 gate1672(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1673(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1674(.a(G657), .O(gate270inter7));
  inv1  gate1675(.a(G785), .O(gate270inter8));
  nand2 gate1676(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1677(.a(s_161), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1678(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1679(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1680(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1457(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1458(.a(gate275inter0), .b(s_130), .O(gate275inter1));
  and2  gate1459(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1460(.a(s_130), .O(gate275inter3));
  inv1  gate1461(.a(s_131), .O(gate275inter4));
  nand2 gate1462(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1463(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1464(.a(G645), .O(gate275inter7));
  inv1  gate1465(.a(G797), .O(gate275inter8));
  nand2 gate1466(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1467(.a(s_131), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1468(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1469(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1470(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1751(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1752(.a(gate277inter0), .b(s_172), .O(gate277inter1));
  and2  gate1753(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1754(.a(s_172), .O(gate277inter3));
  inv1  gate1755(.a(s_173), .O(gate277inter4));
  nand2 gate1756(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1757(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1758(.a(G648), .O(gate277inter7));
  inv1  gate1759(.a(G800), .O(gate277inter8));
  nand2 gate1760(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1761(.a(s_173), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1762(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1763(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1764(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1401(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1402(.a(gate279inter0), .b(s_122), .O(gate279inter1));
  and2  gate1403(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1404(.a(s_122), .O(gate279inter3));
  inv1  gate1405(.a(s_123), .O(gate279inter4));
  nand2 gate1406(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1407(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1408(.a(G651), .O(gate279inter7));
  inv1  gate1409(.a(G803), .O(gate279inter8));
  nand2 gate1410(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1411(.a(s_123), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1412(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1413(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1414(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1933(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1934(.a(gate292inter0), .b(s_198), .O(gate292inter1));
  and2  gate1935(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1936(.a(s_198), .O(gate292inter3));
  inv1  gate1937(.a(s_199), .O(gate292inter4));
  nand2 gate1938(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1939(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1940(.a(G824), .O(gate292inter7));
  inv1  gate1941(.a(G825), .O(gate292inter8));
  nand2 gate1942(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1943(.a(s_199), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1944(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1945(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1946(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate687(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate688(.a(gate293inter0), .b(s_20), .O(gate293inter1));
  and2  gate689(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate690(.a(s_20), .O(gate293inter3));
  inv1  gate691(.a(s_21), .O(gate293inter4));
  nand2 gate692(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate693(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate694(.a(G828), .O(gate293inter7));
  inv1  gate695(.a(G829), .O(gate293inter8));
  nand2 gate696(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate697(.a(s_21), .b(gate293inter3), .O(gate293inter10));
  nor2  gate698(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate699(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate700(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1247(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1248(.a(gate294inter0), .b(s_100), .O(gate294inter1));
  and2  gate1249(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1250(.a(s_100), .O(gate294inter3));
  inv1  gate1251(.a(s_101), .O(gate294inter4));
  nand2 gate1252(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1253(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1254(.a(G832), .O(gate294inter7));
  inv1  gate1255(.a(G833), .O(gate294inter8));
  nand2 gate1256(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1257(.a(s_101), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1258(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1259(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1260(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1345(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1346(.a(gate295inter0), .b(s_114), .O(gate295inter1));
  and2  gate1347(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1348(.a(s_114), .O(gate295inter3));
  inv1  gate1349(.a(s_115), .O(gate295inter4));
  nand2 gate1350(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1351(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1352(.a(G830), .O(gate295inter7));
  inv1  gate1353(.a(G831), .O(gate295inter8));
  nand2 gate1354(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1355(.a(s_115), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1356(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1357(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1358(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1415(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1416(.a(gate388inter0), .b(s_124), .O(gate388inter1));
  and2  gate1417(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1418(.a(s_124), .O(gate388inter3));
  inv1  gate1419(.a(s_125), .O(gate388inter4));
  nand2 gate1420(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1421(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1422(.a(G2), .O(gate388inter7));
  inv1  gate1423(.a(G1039), .O(gate388inter8));
  nand2 gate1424(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1425(.a(s_125), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1426(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1427(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1428(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1373(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1374(.a(gate390inter0), .b(s_118), .O(gate390inter1));
  and2  gate1375(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1376(.a(s_118), .O(gate390inter3));
  inv1  gate1377(.a(s_119), .O(gate390inter4));
  nand2 gate1378(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1379(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1380(.a(G4), .O(gate390inter7));
  inv1  gate1381(.a(G1045), .O(gate390inter8));
  nand2 gate1382(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1383(.a(s_119), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1384(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1385(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1386(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate925(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate926(.a(gate397inter0), .b(s_54), .O(gate397inter1));
  and2  gate927(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate928(.a(s_54), .O(gate397inter3));
  inv1  gate929(.a(s_55), .O(gate397inter4));
  nand2 gate930(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate931(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate932(.a(G11), .O(gate397inter7));
  inv1  gate933(.a(G1066), .O(gate397inter8));
  nand2 gate934(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate935(.a(s_55), .b(gate397inter3), .O(gate397inter10));
  nor2  gate936(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate937(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate938(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1065(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1066(.a(gate400inter0), .b(s_74), .O(gate400inter1));
  and2  gate1067(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1068(.a(s_74), .O(gate400inter3));
  inv1  gate1069(.a(s_75), .O(gate400inter4));
  nand2 gate1070(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1071(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1072(.a(G14), .O(gate400inter7));
  inv1  gate1073(.a(G1075), .O(gate400inter8));
  nand2 gate1074(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1075(.a(s_75), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1076(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1077(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1078(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1051(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1052(.a(gate406inter0), .b(s_72), .O(gate406inter1));
  and2  gate1053(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1054(.a(s_72), .O(gate406inter3));
  inv1  gate1055(.a(s_73), .O(gate406inter4));
  nand2 gate1056(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1057(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1058(.a(G20), .O(gate406inter7));
  inv1  gate1059(.a(G1093), .O(gate406inter8));
  nand2 gate1060(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1061(.a(s_73), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1062(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1063(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1064(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate603(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate604(.a(gate418inter0), .b(s_8), .O(gate418inter1));
  and2  gate605(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate606(.a(s_8), .O(gate418inter3));
  inv1  gate607(.a(s_9), .O(gate418inter4));
  nand2 gate608(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate609(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate610(.a(G32), .O(gate418inter7));
  inv1  gate611(.a(G1129), .O(gate418inter8));
  nand2 gate612(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate613(.a(s_9), .b(gate418inter3), .O(gate418inter10));
  nor2  gate614(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate615(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate616(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1793(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1794(.a(gate419inter0), .b(s_178), .O(gate419inter1));
  and2  gate1795(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1796(.a(s_178), .O(gate419inter3));
  inv1  gate1797(.a(s_179), .O(gate419inter4));
  nand2 gate1798(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1799(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1800(.a(G1), .O(gate419inter7));
  inv1  gate1801(.a(G1132), .O(gate419inter8));
  nand2 gate1802(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1803(.a(s_179), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1804(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1805(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1806(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1639(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1640(.a(gate421inter0), .b(s_156), .O(gate421inter1));
  and2  gate1641(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1642(.a(s_156), .O(gate421inter3));
  inv1  gate1643(.a(s_157), .O(gate421inter4));
  nand2 gate1644(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1645(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1646(.a(G2), .O(gate421inter7));
  inv1  gate1647(.a(G1135), .O(gate421inter8));
  nand2 gate1648(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1649(.a(s_157), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1650(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1651(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1652(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1555(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1556(.a(gate422inter0), .b(s_144), .O(gate422inter1));
  and2  gate1557(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1558(.a(s_144), .O(gate422inter3));
  inv1  gate1559(.a(s_145), .O(gate422inter4));
  nand2 gate1560(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1561(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1562(.a(G1039), .O(gate422inter7));
  inv1  gate1563(.a(G1135), .O(gate422inter8));
  nand2 gate1564(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1565(.a(s_145), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1566(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1567(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1568(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate827(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate828(.a(gate427inter0), .b(s_40), .O(gate427inter1));
  and2  gate829(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate830(.a(s_40), .O(gate427inter3));
  inv1  gate831(.a(s_41), .O(gate427inter4));
  nand2 gate832(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate833(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate834(.a(G5), .O(gate427inter7));
  inv1  gate835(.a(G1144), .O(gate427inter8));
  nand2 gate836(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate837(.a(s_41), .b(gate427inter3), .O(gate427inter10));
  nor2  gate838(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate839(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate840(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate883(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate884(.a(gate436inter0), .b(s_48), .O(gate436inter1));
  and2  gate885(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate886(.a(s_48), .O(gate436inter3));
  inv1  gate887(.a(s_49), .O(gate436inter4));
  nand2 gate888(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate889(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate890(.a(G1060), .O(gate436inter7));
  inv1  gate891(.a(G1156), .O(gate436inter8));
  nand2 gate892(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate893(.a(s_49), .b(gate436inter3), .O(gate436inter10));
  nor2  gate894(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate895(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate896(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate589(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate590(.a(gate437inter0), .b(s_6), .O(gate437inter1));
  and2  gate591(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate592(.a(s_6), .O(gate437inter3));
  inv1  gate593(.a(s_7), .O(gate437inter4));
  nand2 gate594(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate595(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate596(.a(G10), .O(gate437inter7));
  inv1  gate597(.a(G1159), .O(gate437inter8));
  nand2 gate598(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate599(.a(s_7), .b(gate437inter3), .O(gate437inter10));
  nor2  gate600(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate601(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate602(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate869(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate870(.a(gate438inter0), .b(s_46), .O(gate438inter1));
  and2  gate871(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate872(.a(s_46), .O(gate438inter3));
  inv1  gate873(.a(s_47), .O(gate438inter4));
  nand2 gate874(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate875(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate876(.a(G1063), .O(gate438inter7));
  inv1  gate877(.a(G1159), .O(gate438inter8));
  nand2 gate878(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate879(.a(s_47), .b(gate438inter3), .O(gate438inter10));
  nor2  gate880(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate881(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate882(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1205(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1206(.a(gate441inter0), .b(s_94), .O(gate441inter1));
  and2  gate1207(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1208(.a(s_94), .O(gate441inter3));
  inv1  gate1209(.a(s_95), .O(gate441inter4));
  nand2 gate1210(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1211(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1212(.a(G12), .O(gate441inter7));
  inv1  gate1213(.a(G1165), .O(gate441inter8));
  nand2 gate1214(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1215(.a(s_95), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1216(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1217(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1218(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1289(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1290(.a(gate442inter0), .b(s_106), .O(gate442inter1));
  and2  gate1291(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1292(.a(s_106), .O(gate442inter3));
  inv1  gate1293(.a(s_107), .O(gate442inter4));
  nand2 gate1294(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1295(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1296(.a(G1069), .O(gate442inter7));
  inv1  gate1297(.a(G1165), .O(gate442inter8));
  nand2 gate1298(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1299(.a(s_107), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1300(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1301(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1302(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1387(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1388(.a(gate452inter0), .b(s_120), .O(gate452inter1));
  and2  gate1389(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1390(.a(s_120), .O(gate452inter3));
  inv1  gate1391(.a(s_121), .O(gate452inter4));
  nand2 gate1392(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1393(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1394(.a(G1084), .O(gate452inter7));
  inv1  gate1395(.a(G1180), .O(gate452inter8));
  nand2 gate1396(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1397(.a(s_121), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1398(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1399(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1400(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate799(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate800(.a(gate453inter0), .b(s_36), .O(gate453inter1));
  and2  gate801(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate802(.a(s_36), .O(gate453inter3));
  inv1  gate803(.a(s_37), .O(gate453inter4));
  nand2 gate804(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate805(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate806(.a(G18), .O(gate453inter7));
  inv1  gate807(.a(G1183), .O(gate453inter8));
  nand2 gate808(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate809(.a(s_37), .b(gate453inter3), .O(gate453inter10));
  nor2  gate810(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate811(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate812(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate967(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate968(.a(gate460inter0), .b(s_60), .O(gate460inter1));
  and2  gate969(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate970(.a(s_60), .O(gate460inter3));
  inv1  gate971(.a(s_61), .O(gate460inter4));
  nand2 gate972(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate973(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate974(.a(G1096), .O(gate460inter7));
  inv1  gate975(.a(G1192), .O(gate460inter8));
  nand2 gate976(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate977(.a(s_61), .b(gate460inter3), .O(gate460inter10));
  nor2  gate978(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate979(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate980(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate785(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate786(.a(gate467inter0), .b(s_34), .O(gate467inter1));
  and2  gate787(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate788(.a(s_34), .O(gate467inter3));
  inv1  gate789(.a(s_35), .O(gate467inter4));
  nand2 gate790(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate791(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate792(.a(G25), .O(gate467inter7));
  inv1  gate793(.a(G1204), .O(gate467inter8));
  nand2 gate794(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate795(.a(s_35), .b(gate467inter3), .O(gate467inter10));
  nor2  gate796(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate797(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate798(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1233(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1234(.a(gate468inter0), .b(s_98), .O(gate468inter1));
  and2  gate1235(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1236(.a(s_98), .O(gate468inter3));
  inv1  gate1237(.a(s_99), .O(gate468inter4));
  nand2 gate1238(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1239(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1240(.a(G1108), .O(gate468inter7));
  inv1  gate1241(.a(G1204), .O(gate468inter8));
  nand2 gate1242(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1243(.a(s_99), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1244(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1245(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1246(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate631(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate632(.a(gate473inter0), .b(s_12), .O(gate473inter1));
  and2  gate633(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate634(.a(s_12), .O(gate473inter3));
  inv1  gate635(.a(s_13), .O(gate473inter4));
  nand2 gate636(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate637(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate638(.a(G28), .O(gate473inter7));
  inv1  gate639(.a(G1213), .O(gate473inter8));
  nand2 gate640(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate641(.a(s_13), .b(gate473inter3), .O(gate473inter10));
  nor2  gate642(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate643(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate644(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1905(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1906(.a(gate476inter0), .b(s_194), .O(gate476inter1));
  and2  gate1907(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1908(.a(s_194), .O(gate476inter3));
  inv1  gate1909(.a(s_195), .O(gate476inter4));
  nand2 gate1910(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1911(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1912(.a(G1120), .O(gate476inter7));
  inv1  gate1913(.a(G1216), .O(gate476inter8));
  nand2 gate1914(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1915(.a(s_195), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1916(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1917(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1918(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1695(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1696(.a(gate482inter0), .b(s_164), .O(gate482inter1));
  and2  gate1697(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1698(.a(s_164), .O(gate482inter3));
  inv1  gate1699(.a(s_165), .O(gate482inter4));
  nand2 gate1700(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1701(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1702(.a(G1129), .O(gate482inter7));
  inv1  gate1703(.a(G1225), .O(gate482inter8));
  nand2 gate1704(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1705(.a(s_165), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1706(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1707(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1708(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1821(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1822(.a(gate485inter0), .b(s_182), .O(gate485inter1));
  and2  gate1823(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1824(.a(s_182), .O(gate485inter3));
  inv1  gate1825(.a(s_183), .O(gate485inter4));
  nand2 gate1826(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1827(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1828(.a(G1232), .O(gate485inter7));
  inv1  gate1829(.a(G1233), .O(gate485inter8));
  nand2 gate1830(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1831(.a(s_183), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1832(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1833(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1834(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate673(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate674(.a(gate489inter0), .b(s_18), .O(gate489inter1));
  and2  gate675(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate676(.a(s_18), .O(gate489inter3));
  inv1  gate677(.a(s_19), .O(gate489inter4));
  nand2 gate678(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate679(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate680(.a(G1240), .O(gate489inter7));
  inv1  gate681(.a(G1241), .O(gate489inter8));
  nand2 gate682(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate683(.a(s_19), .b(gate489inter3), .O(gate489inter10));
  nor2  gate684(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate685(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate686(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1765(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1766(.a(gate492inter0), .b(s_174), .O(gate492inter1));
  and2  gate1767(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1768(.a(s_174), .O(gate492inter3));
  inv1  gate1769(.a(s_175), .O(gate492inter4));
  nand2 gate1770(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1771(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1772(.a(G1246), .O(gate492inter7));
  inv1  gate1773(.a(G1247), .O(gate492inter8));
  nand2 gate1774(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1775(.a(s_175), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1776(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1777(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1778(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1037(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1038(.a(gate496inter0), .b(s_70), .O(gate496inter1));
  and2  gate1039(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1040(.a(s_70), .O(gate496inter3));
  inv1  gate1041(.a(s_71), .O(gate496inter4));
  nand2 gate1042(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1043(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1044(.a(G1254), .O(gate496inter7));
  inv1  gate1045(.a(G1255), .O(gate496inter8));
  nand2 gate1046(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1047(.a(s_71), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1048(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1049(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1050(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1681(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1682(.a(gate500inter0), .b(s_162), .O(gate500inter1));
  and2  gate1683(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1684(.a(s_162), .O(gate500inter3));
  inv1  gate1685(.a(s_163), .O(gate500inter4));
  nand2 gate1686(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1687(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1688(.a(G1262), .O(gate500inter7));
  inv1  gate1689(.a(G1263), .O(gate500inter8));
  nand2 gate1690(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1691(.a(s_163), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1692(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1693(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1694(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1597(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1598(.a(gate510inter0), .b(s_150), .O(gate510inter1));
  and2  gate1599(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1600(.a(s_150), .O(gate510inter3));
  inv1  gate1601(.a(s_151), .O(gate510inter4));
  nand2 gate1602(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1603(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1604(.a(G1282), .O(gate510inter7));
  inv1  gate1605(.a(G1283), .O(gate510inter8));
  nand2 gate1606(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1607(.a(s_151), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1608(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1609(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1610(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1303(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1304(.a(gate511inter0), .b(s_108), .O(gate511inter1));
  and2  gate1305(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1306(.a(s_108), .O(gate511inter3));
  inv1  gate1307(.a(s_109), .O(gate511inter4));
  nand2 gate1308(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1309(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1310(.a(G1284), .O(gate511inter7));
  inv1  gate1311(.a(G1285), .O(gate511inter8));
  nand2 gate1312(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1313(.a(s_109), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1314(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1315(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1316(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule