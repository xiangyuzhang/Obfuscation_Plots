module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );

  xor2  gate469(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate470(.a(gate20inter0), .b(s_44), .O(gate20inter1));
  and2  gate471(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate472(.a(s_44), .O(gate20inter3));
  inv1  gate473(.a(s_45), .O(gate20inter4));
  nand2 gate474(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate475(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate476(.a(N8), .O(gate20inter7));
  inv1  gate477(.a(N119), .O(gate20inter8));
  nand2 gate478(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate479(.a(s_45), .b(gate20inter3), .O(gate20inter10));
  nor2  gate480(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate481(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate482(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate343(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate344(.a(gate27inter0), .b(s_26), .O(gate27inter1));
  and2  gate345(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate346(.a(s_26), .O(gate27inter3));
  inv1  gate347(.a(s_27), .O(gate27inter4));
  nand2 gate348(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate349(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate350(.a(N142), .O(gate27inter7));
  inv1  gate351(.a(N82), .O(gate27inter8));
  nand2 gate352(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate353(.a(s_27), .b(gate27inter3), .O(gate27inter10));
  nor2  gate354(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate355(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate356(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate175(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate176(.a(gate37inter0), .b(s_2), .O(gate37inter1));
  and2  gate177(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate178(.a(s_2), .O(gate37inter3));
  inv1  gate179(.a(s_3), .O(gate37inter4));
  nand2 gate180(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate181(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate182(.a(N66), .O(gate37inter7));
  inv1  gate183(.a(N135), .O(gate37inter8));
  nand2 gate184(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate185(.a(s_3), .b(gate37inter3), .O(gate37inter10));
  nor2  gate186(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate187(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate188(.a(gate37inter12), .b(gate37inter1), .O(N190));

  xor2  gate497(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate498(.a(gate38inter0), .b(s_48), .O(gate38inter1));
  and2  gate499(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate500(.a(s_48), .O(gate38inter3));
  inv1  gate501(.a(s_49), .O(gate38inter4));
  nand2 gate502(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate503(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate504(.a(N73), .O(gate38inter7));
  inv1  gate505(.a(N139), .O(gate38inter8));
  nand2 gate506(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate507(.a(s_49), .b(gate38inter3), .O(gate38inter10));
  nor2  gate508(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate509(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate510(.a(gate38inter12), .b(gate38inter1), .O(N191));
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate413(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate414(.a(gate62inter0), .b(s_36), .O(gate62inter1));
  and2  gate415(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate416(.a(s_36), .O(gate62inter3));
  inv1  gate417(.a(s_37), .O(gate62inter4));
  nand2 gate418(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate419(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate420(.a(N213), .O(gate62inter7));
  inv1  gate421(.a(N37), .O(gate62inter8));
  nand2 gate422(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate423(.a(s_37), .b(gate62inter3), .O(gate62inter10));
  nor2  gate424(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate425(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate426(.a(gate62inter12), .b(gate62inter1), .O(N254));

  xor2  gate455(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate456(.a(gate63inter0), .b(s_42), .O(gate63inter1));
  and2  gate457(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate458(.a(s_42), .O(gate63inter3));
  inv1  gate459(.a(s_43), .O(gate63inter4));
  nand2 gate460(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate461(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate462(.a(N213), .O(gate63inter7));
  inv1  gate463(.a(N50), .O(gate63inter8));
  nand2 gate464(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate465(.a(s_43), .b(gate63inter3), .O(gate63inter10));
  nor2  gate466(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate467(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate468(.a(gate63inter12), .b(gate63inter1), .O(N255));
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate567(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate568(.a(gate65inter0), .b(s_58), .O(gate65inter1));
  and2  gate569(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate570(.a(s_58), .O(gate65inter3));
  inv1  gate571(.a(s_59), .O(gate65inter4));
  nand2 gate572(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate573(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate574(.a(N213), .O(gate65inter7));
  inv1  gate575(.a(N76), .O(gate65inter8));
  nand2 gate576(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate577(.a(s_59), .b(gate65inter3), .O(gate65inter10));
  nor2  gate578(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate579(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate580(.a(gate65inter12), .b(gate65inter1), .O(N257));
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );

  xor2  gate511(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate512(.a(gate69inter0), .b(s_50), .O(gate69inter1));
  and2  gate513(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate514(.a(s_50), .O(gate69inter3));
  inv1  gate515(.a(s_51), .O(gate69inter4));
  nand2 gate516(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate517(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate518(.a(N224), .O(gate69inter7));
  inv1  gate519(.a(N158), .O(gate69inter8));
  nand2 gate520(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate521(.a(s_51), .b(gate69inter3), .O(gate69inter10));
  nor2  gate522(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate523(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate524(.a(gate69inter12), .b(gate69inter1), .O(N263));
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate315(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate316(.a(gate71inter0), .b(s_22), .O(gate71inter1));
  and2  gate317(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate318(.a(s_22), .O(gate71inter3));
  inv1  gate319(.a(s_23), .O(gate71inter4));
  nand2 gate320(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate321(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate322(.a(N230), .O(gate71inter7));
  inv1  gate323(.a(N185), .O(gate71inter8));
  nand2 gate324(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate325(.a(s_23), .b(gate71inter3), .O(gate71inter10));
  nor2  gate326(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate327(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate328(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate329(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate330(.a(gate73inter0), .b(s_24), .O(gate73inter1));
  and2  gate331(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate332(.a(s_24), .O(gate73inter3));
  inv1  gate333(.a(s_25), .O(gate73inter4));
  nand2 gate334(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate335(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate336(.a(N236), .O(gate73inter7));
  inv1  gate337(.a(N189), .O(gate73inter8));
  nand2 gate338(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate339(.a(s_25), .b(gate73inter3), .O(gate73inter10));
  nor2  gate340(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate341(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate342(.a(gate73inter12), .b(gate73inter1), .O(N273));

  xor2  gate371(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate372(.a(gate74inter0), .b(s_30), .O(gate74inter1));
  and2  gate373(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate374(.a(s_30), .O(gate74inter3));
  inv1  gate375(.a(s_31), .O(gate74inter4));
  nand2 gate376(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate377(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate378(.a(N239), .O(gate74inter7));
  inv1  gate379(.a(N191), .O(gate74inter8));
  nand2 gate380(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate381(.a(s_31), .b(gate74inter3), .O(gate74inter10));
  nor2  gate382(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate383(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate384(.a(gate74inter12), .b(gate74inter1), .O(N276));

  xor2  gate231(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate232(.a(gate75inter0), .b(s_10), .O(gate75inter1));
  and2  gate233(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate234(.a(s_10), .O(gate75inter3));
  inv1  gate235(.a(s_11), .O(gate75inter4));
  nand2 gate236(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate237(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate238(.a(N243), .O(gate75inter7));
  inv1  gate239(.a(N193), .O(gate75inter8));
  nand2 gate240(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate241(.a(s_11), .b(gate75inter3), .O(gate75inter10));
  nor2  gate242(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate243(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate244(.a(gate75inter12), .b(gate75inter1), .O(N279));

  xor2  gate441(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate442(.a(gate76inter0), .b(s_40), .O(gate76inter1));
  and2  gate443(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate444(.a(s_40), .O(gate76inter3));
  inv1  gate445(.a(s_41), .O(gate76inter4));
  nand2 gate446(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate447(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate448(.a(N247), .O(gate76inter7));
  inv1  gate449(.a(N195), .O(gate76inter8));
  nand2 gate450(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate451(.a(s_41), .b(gate76inter3), .O(gate76inter10));
  nor2  gate452(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate453(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate454(.a(gate76inter12), .b(gate76inter1), .O(N282));

  xor2  gate539(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate540(.a(gate77inter0), .b(s_54), .O(gate77inter1));
  and2  gate541(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate542(.a(s_54), .O(gate77inter3));
  inv1  gate543(.a(s_55), .O(gate77inter4));
  nand2 gate544(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate545(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate546(.a(N251), .O(gate77inter7));
  inv1  gate547(.a(N197), .O(gate77inter8));
  nand2 gate548(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate549(.a(s_55), .b(gate77inter3), .O(gate77inter10));
  nor2  gate550(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate551(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate552(.a(gate77inter12), .b(gate77inter1), .O(N285));

  xor2  gate399(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate400(.a(gate78inter0), .b(s_34), .O(gate78inter1));
  and2  gate401(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate402(.a(s_34), .O(gate78inter3));
  inv1  gate403(.a(s_35), .O(gate78inter4));
  nand2 gate404(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate405(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate406(.a(N227), .O(gate78inter7));
  inv1  gate407(.a(N184), .O(gate78inter8));
  nand2 gate408(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate409(.a(s_35), .b(gate78inter3), .O(gate78inter10));
  nor2  gate410(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate411(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate412(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );

  xor2  gate189(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate190(.a(gate81inter0), .b(s_4), .O(gate81inter1));
  and2  gate191(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate192(.a(s_4), .O(gate81inter3));
  inv1  gate193(.a(s_5), .O(gate81inter4));
  nand2 gate194(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate195(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate196(.a(N236), .O(gate81inter7));
  inv1  gate197(.a(N190), .O(gate81inter8));
  nand2 gate198(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate199(.a(s_5), .b(gate81inter3), .O(gate81inter10));
  nor2  gate200(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate201(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate202(.a(gate81inter12), .b(gate81inter1), .O(N291));

  xor2  gate483(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate484(.a(gate82inter0), .b(s_46), .O(gate82inter1));
  and2  gate485(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate486(.a(s_46), .O(gate82inter3));
  inv1  gate487(.a(s_47), .O(gate82inter4));
  nand2 gate488(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate489(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate490(.a(N239), .O(gate82inter7));
  inv1  gate491(.a(N192), .O(gate82inter8));
  nand2 gate492(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate493(.a(s_47), .b(gate82inter3), .O(gate82inter10));
  nor2  gate494(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate495(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate496(.a(gate82inter12), .b(gate82inter1), .O(N292));

  xor2  gate259(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate260(.a(gate83inter0), .b(s_14), .O(gate83inter1));
  and2  gate261(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate262(.a(s_14), .O(gate83inter3));
  inv1  gate263(.a(s_15), .O(gate83inter4));
  nand2 gate264(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate265(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate266(.a(N243), .O(gate83inter7));
  inv1  gate267(.a(N194), .O(gate83inter8));
  nand2 gate268(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate269(.a(s_15), .b(gate83inter3), .O(gate83inter10));
  nor2  gate270(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate271(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate272(.a(gate83inter12), .b(gate83inter1), .O(N293));

  xor2  gate385(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate386(.a(gate84inter0), .b(s_32), .O(gate84inter1));
  and2  gate387(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate388(.a(s_32), .O(gate84inter3));
  inv1  gate389(.a(s_33), .O(gate84inter4));
  nand2 gate390(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate391(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate392(.a(N247), .O(gate84inter7));
  inv1  gate393(.a(N196), .O(gate84inter8));
  nand2 gate394(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate395(.a(s_33), .b(gate84inter3), .O(gate84inter10));
  nor2  gate396(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate397(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate398(.a(gate84inter12), .b(gate84inter1), .O(N294));

  xor2  gate203(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate204(.a(gate85inter0), .b(s_6), .O(gate85inter1));
  and2  gate205(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate206(.a(s_6), .O(gate85inter3));
  inv1  gate207(.a(s_7), .O(gate85inter4));
  nand2 gate208(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate209(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate210(.a(N251), .O(gate85inter7));
  inv1  gate211(.a(N198), .O(gate85inter8));
  nand2 gate212(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate213(.a(s_7), .b(gate85inter3), .O(gate85inter10));
  nor2  gate214(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate215(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate216(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );

  xor2  gate301(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate302(.a(gate100inter0), .b(s_20), .O(gate100inter1));
  and2  gate303(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate304(.a(s_20), .O(gate100inter3));
  inv1  gate305(.a(s_21), .O(gate100inter4));
  nand2 gate306(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate307(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate308(.a(N309), .O(gate100inter7));
  inv1  gate309(.a(N264), .O(gate100inter8));
  nand2 gate310(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate311(.a(s_21), .b(gate100inter3), .O(gate100inter10));
  nor2  gate312(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate313(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate314(.a(gate100inter12), .b(gate100inter1), .O(N331));
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );

  xor2  gate553(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate554(.a(gate104inter0), .b(s_56), .O(gate104inter1));
  and2  gate555(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate556(.a(s_56), .O(gate104inter3));
  inv1  gate557(.a(s_57), .O(gate104inter4));
  nand2 gate558(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate559(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate560(.a(N309), .O(gate104inter7));
  inv1  gate561(.a(N273), .O(gate104inter8));
  nand2 gate562(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate563(.a(s_57), .b(gate104inter3), .O(gate104inter10));
  nor2  gate564(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate565(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate566(.a(gate104inter12), .b(gate104inter1), .O(N335));

  xor2  gate245(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate246(.a(gate105inter0), .b(s_12), .O(gate105inter1));
  and2  gate247(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate248(.a(s_12), .O(gate105inter3));
  inv1  gate249(.a(s_13), .O(gate105inter4));
  nand2 gate250(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate251(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate252(.a(N319), .O(gate105inter7));
  inv1  gate253(.a(N21), .O(gate105inter8));
  nand2 gate254(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate255(.a(s_13), .b(gate105inter3), .O(gate105inter10));
  nor2  gate256(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate257(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate258(.a(gate105inter12), .b(gate105inter1), .O(N336));

  xor2  gate427(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate428(.a(gate106inter0), .b(s_38), .O(gate106inter1));
  and2  gate429(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate430(.a(s_38), .O(gate106inter3));
  inv1  gate431(.a(s_39), .O(gate106inter4));
  nand2 gate432(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate433(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate434(.a(N309), .O(gate106inter7));
  inv1  gate435(.a(N276), .O(gate106inter8));
  nand2 gate436(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate437(.a(s_39), .b(gate106inter3), .O(gate106inter10));
  nor2  gate438(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate439(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate440(.a(gate106inter12), .b(gate106inter1), .O(N337));
nand2 gate107( .a(N319), .b(N34), .O(N338) );

  xor2  gate287(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate288(.a(gate108inter0), .b(s_18), .O(gate108inter1));
  and2  gate289(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate290(.a(s_18), .O(gate108inter3));
  inv1  gate291(.a(s_19), .O(gate108inter4));
  nand2 gate292(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate293(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate294(.a(N309), .O(gate108inter7));
  inv1  gate295(.a(N279), .O(gate108inter8));
  nand2 gate296(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate297(.a(s_19), .b(gate108inter3), .O(gate108inter10));
  nor2  gate298(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate299(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate300(.a(gate108inter12), .b(gate108inter1), .O(N339));
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate525(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate526(.a(gate111inter0), .b(s_52), .O(gate111inter1));
  and2  gate527(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate528(.a(s_52), .O(gate111inter3));
  inv1  gate529(.a(s_53), .O(gate111inter4));
  nand2 gate530(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate531(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate532(.a(N319), .O(gate111inter7));
  inv1  gate533(.a(N60), .O(gate111inter8));
  nand2 gate534(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate535(.a(s_53), .b(gate111inter3), .O(gate111inter10));
  nor2  gate536(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate537(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate538(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );

  xor2  gate161(.a(N86), .b(N319), .O(gate114inter0));
  nand2 gate162(.a(gate114inter0), .b(s_0), .O(gate114inter1));
  and2  gate163(.a(N86), .b(N319), .O(gate114inter2));
  inv1  gate164(.a(s_0), .O(gate114inter3));
  inv1  gate165(.a(s_1), .O(gate114inter4));
  nand2 gate166(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate167(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate168(.a(N319), .O(gate114inter7));
  inv1  gate169(.a(N86), .O(gate114inter8));
  nand2 gate170(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate171(.a(s_1), .b(gate114inter3), .O(gate114inter10));
  nor2  gate172(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate173(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate174(.a(gate114inter12), .b(gate114inter1), .O(N345));
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate581(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate582(.a(gate118inter0), .b(s_60), .O(gate118inter1));
  and2  gate583(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate584(.a(s_60), .O(gate118inter3));
  inv1  gate585(.a(s_61), .O(gate118inter4));
  nand2 gate586(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate587(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate588(.a(N331), .O(gate118inter7));
  inv1  gate589(.a(N301), .O(gate118inter8));
  nand2 gate590(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate591(.a(s_61), .b(gate118inter3), .O(gate118inter10));
  nor2  gate592(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate593(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate594(.a(gate118inter12), .b(gate118inter1), .O(N349));
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );

  xor2  gate217(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate218(.a(gate125inter0), .b(s_8), .O(gate125inter1));
  and2  gate219(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate220(.a(s_8), .O(gate125inter3));
  inv1  gate221(.a(s_9), .O(gate125inter4));
  nand2 gate222(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate223(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate224(.a(N343), .O(gate125inter7));
  inv1  gate225(.a(N308), .O(gate125inter8));
  nand2 gate226(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate227(.a(s_9), .b(gate125inter3), .O(gate125inter10));
  nor2  gate228(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate229(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate230(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate357(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate358(.a(gate131inter0), .b(s_28), .O(gate131inter1));
  and2  gate359(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate360(.a(s_28), .O(gate131inter3));
  inv1  gate361(.a(s_29), .O(gate131inter4));
  nand2 gate362(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate363(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate364(.a(N360), .O(gate131inter7));
  inv1  gate365(.a(N40), .O(gate131inter8));
  nand2 gate366(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate367(.a(s_29), .b(gate131inter3), .O(gate131inter10));
  nor2  gate368(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate369(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate370(.a(gate131inter12), .b(gate131inter1), .O(N373));
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate273(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate274(.a(gate136inter0), .b(s_16), .O(gate136inter1));
  and2  gate275(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate276(.a(s_16), .O(gate136inter3));
  inv1  gate277(.a(s_17), .O(gate136inter4));
  nand2 gate278(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate279(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate280(.a(N360), .O(gate136inter7));
  inv1  gate281(.a(N105), .O(gate136inter8));
  nand2 gate282(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate283(.a(s_17), .b(gate136inter3), .O(gate136inter10));
  nor2  gate284(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate285(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate286(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule