module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1443(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1444(.a(gate9inter0), .b(s_128), .O(gate9inter1));
  and2  gate1445(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1446(.a(s_128), .O(gate9inter3));
  inv1  gate1447(.a(s_129), .O(gate9inter4));
  nand2 gate1448(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1449(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1450(.a(G1), .O(gate9inter7));
  inv1  gate1451(.a(G2), .O(gate9inter8));
  nand2 gate1452(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1453(.a(s_129), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1454(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1455(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1456(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate673(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate674(.a(gate10inter0), .b(s_18), .O(gate10inter1));
  and2  gate675(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate676(.a(s_18), .O(gate10inter3));
  inv1  gate677(.a(s_19), .O(gate10inter4));
  nand2 gate678(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate679(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate680(.a(G3), .O(gate10inter7));
  inv1  gate681(.a(G4), .O(gate10inter8));
  nand2 gate682(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate683(.a(s_19), .b(gate10inter3), .O(gate10inter10));
  nor2  gate684(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate685(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate686(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate1765(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1766(.a(gate11inter0), .b(s_174), .O(gate11inter1));
  and2  gate1767(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1768(.a(s_174), .O(gate11inter3));
  inv1  gate1769(.a(s_175), .O(gate11inter4));
  nand2 gate1770(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1771(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1772(.a(G5), .O(gate11inter7));
  inv1  gate1773(.a(G6), .O(gate11inter8));
  nand2 gate1774(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1775(.a(s_175), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1776(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1777(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1778(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2087(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2088(.a(gate12inter0), .b(s_220), .O(gate12inter1));
  and2  gate2089(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2090(.a(s_220), .O(gate12inter3));
  inv1  gate2091(.a(s_221), .O(gate12inter4));
  nand2 gate2092(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2093(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2094(.a(G7), .O(gate12inter7));
  inv1  gate2095(.a(G8), .O(gate12inter8));
  nand2 gate2096(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2097(.a(s_221), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2098(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2099(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2100(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1625(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1626(.a(gate13inter0), .b(s_154), .O(gate13inter1));
  and2  gate1627(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1628(.a(s_154), .O(gate13inter3));
  inv1  gate1629(.a(s_155), .O(gate13inter4));
  nand2 gate1630(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1631(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1632(.a(G9), .O(gate13inter7));
  inv1  gate1633(.a(G10), .O(gate13inter8));
  nand2 gate1634(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1635(.a(s_155), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1636(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1637(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1638(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate967(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate968(.a(gate15inter0), .b(s_60), .O(gate15inter1));
  and2  gate969(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate970(.a(s_60), .O(gate15inter3));
  inv1  gate971(.a(s_61), .O(gate15inter4));
  nand2 gate972(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate973(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate974(.a(G13), .O(gate15inter7));
  inv1  gate975(.a(G14), .O(gate15inter8));
  nand2 gate976(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate977(.a(s_61), .b(gate15inter3), .O(gate15inter10));
  nor2  gate978(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate979(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate980(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1863(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1864(.a(gate17inter0), .b(s_188), .O(gate17inter1));
  and2  gate1865(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1866(.a(s_188), .O(gate17inter3));
  inv1  gate1867(.a(s_189), .O(gate17inter4));
  nand2 gate1868(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1869(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1870(.a(G17), .O(gate17inter7));
  inv1  gate1871(.a(G18), .O(gate17inter8));
  nand2 gate1872(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1873(.a(s_189), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1874(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1875(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1876(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1849(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1850(.a(gate19inter0), .b(s_186), .O(gate19inter1));
  and2  gate1851(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1852(.a(s_186), .O(gate19inter3));
  inv1  gate1853(.a(s_187), .O(gate19inter4));
  nand2 gate1854(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1855(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1856(.a(G21), .O(gate19inter7));
  inv1  gate1857(.a(G22), .O(gate19inter8));
  nand2 gate1858(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1859(.a(s_187), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1860(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1861(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1862(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1989(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1990(.a(gate22inter0), .b(s_206), .O(gate22inter1));
  and2  gate1991(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1992(.a(s_206), .O(gate22inter3));
  inv1  gate1993(.a(s_207), .O(gate22inter4));
  nand2 gate1994(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1995(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1996(.a(G27), .O(gate22inter7));
  inv1  gate1997(.a(G28), .O(gate22inter8));
  nand2 gate1998(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1999(.a(s_207), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2000(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2001(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2002(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate589(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate590(.a(gate23inter0), .b(s_6), .O(gate23inter1));
  and2  gate591(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate592(.a(s_6), .O(gate23inter3));
  inv1  gate593(.a(s_7), .O(gate23inter4));
  nand2 gate594(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate595(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate596(.a(G29), .O(gate23inter7));
  inv1  gate597(.a(G30), .O(gate23inter8));
  nand2 gate598(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate599(.a(s_7), .b(gate23inter3), .O(gate23inter10));
  nor2  gate600(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate601(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate602(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1975(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1976(.a(gate24inter0), .b(s_204), .O(gate24inter1));
  and2  gate1977(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1978(.a(s_204), .O(gate24inter3));
  inv1  gate1979(.a(s_205), .O(gate24inter4));
  nand2 gate1980(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1981(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1982(.a(G31), .O(gate24inter7));
  inv1  gate1983(.a(G32), .O(gate24inter8));
  nand2 gate1984(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1985(.a(s_205), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1986(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1987(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1988(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2549(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2550(.a(gate27inter0), .b(s_286), .O(gate27inter1));
  and2  gate2551(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2552(.a(s_286), .O(gate27inter3));
  inv1  gate2553(.a(s_287), .O(gate27inter4));
  nand2 gate2554(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2555(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2556(.a(G2), .O(gate27inter7));
  inv1  gate2557(.a(G6), .O(gate27inter8));
  nand2 gate2558(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2559(.a(s_287), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2560(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2561(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2562(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1485(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1486(.a(gate28inter0), .b(s_134), .O(gate28inter1));
  and2  gate1487(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1488(.a(s_134), .O(gate28inter3));
  inv1  gate1489(.a(s_135), .O(gate28inter4));
  nand2 gate1490(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1491(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1492(.a(G10), .O(gate28inter7));
  inv1  gate1493(.a(G14), .O(gate28inter8));
  nand2 gate1494(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1495(.a(s_135), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1496(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1497(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1498(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1527(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1528(.a(gate48inter0), .b(s_140), .O(gate48inter1));
  and2  gate1529(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1530(.a(s_140), .O(gate48inter3));
  inv1  gate1531(.a(s_141), .O(gate48inter4));
  nand2 gate1532(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1533(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1534(.a(G8), .O(gate48inter7));
  inv1  gate1535(.a(G275), .O(gate48inter8));
  nand2 gate1536(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1537(.a(s_141), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1538(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1539(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1540(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate701(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate702(.a(gate52inter0), .b(s_22), .O(gate52inter1));
  and2  gate703(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate704(.a(s_22), .O(gate52inter3));
  inv1  gate705(.a(s_23), .O(gate52inter4));
  nand2 gate706(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate707(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate708(.a(G12), .O(gate52inter7));
  inv1  gate709(.a(G281), .O(gate52inter8));
  nand2 gate710(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate711(.a(s_23), .b(gate52inter3), .O(gate52inter10));
  nor2  gate712(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate713(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate714(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate883(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate884(.a(gate53inter0), .b(s_48), .O(gate53inter1));
  and2  gate885(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate886(.a(s_48), .O(gate53inter3));
  inv1  gate887(.a(s_49), .O(gate53inter4));
  nand2 gate888(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate889(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate890(.a(G13), .O(gate53inter7));
  inv1  gate891(.a(G284), .O(gate53inter8));
  nand2 gate892(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate893(.a(s_49), .b(gate53inter3), .O(gate53inter10));
  nor2  gate894(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate895(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate896(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2227(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2228(.a(gate56inter0), .b(s_240), .O(gate56inter1));
  and2  gate2229(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2230(.a(s_240), .O(gate56inter3));
  inv1  gate2231(.a(s_241), .O(gate56inter4));
  nand2 gate2232(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2233(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2234(.a(G16), .O(gate56inter7));
  inv1  gate2235(.a(G287), .O(gate56inter8));
  nand2 gate2236(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2237(.a(s_241), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2238(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2239(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2240(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate2059(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2060(.a(gate57inter0), .b(s_216), .O(gate57inter1));
  and2  gate2061(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2062(.a(s_216), .O(gate57inter3));
  inv1  gate2063(.a(s_217), .O(gate57inter4));
  nand2 gate2064(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2065(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2066(.a(G17), .O(gate57inter7));
  inv1  gate2067(.a(G290), .O(gate57inter8));
  nand2 gate2068(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2069(.a(s_217), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2070(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2071(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2072(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate827(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate828(.a(gate58inter0), .b(s_40), .O(gate58inter1));
  and2  gate829(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate830(.a(s_40), .O(gate58inter3));
  inv1  gate831(.a(s_41), .O(gate58inter4));
  nand2 gate832(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate833(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate834(.a(G18), .O(gate58inter7));
  inv1  gate835(.a(G290), .O(gate58inter8));
  nand2 gate836(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate837(.a(s_41), .b(gate58inter3), .O(gate58inter10));
  nor2  gate838(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate839(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate840(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate2605(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2606(.a(gate59inter0), .b(s_294), .O(gate59inter1));
  and2  gate2607(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2608(.a(s_294), .O(gate59inter3));
  inv1  gate2609(.a(s_295), .O(gate59inter4));
  nand2 gate2610(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2611(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2612(.a(G19), .O(gate59inter7));
  inv1  gate2613(.a(G293), .O(gate59inter8));
  nand2 gate2614(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2615(.a(s_295), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2616(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2617(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2618(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1681(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1682(.a(gate61inter0), .b(s_162), .O(gate61inter1));
  and2  gate1683(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1684(.a(s_162), .O(gate61inter3));
  inv1  gate1685(.a(s_163), .O(gate61inter4));
  nand2 gate1686(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1687(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1688(.a(G21), .O(gate61inter7));
  inv1  gate1689(.a(G296), .O(gate61inter8));
  nand2 gate1690(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1691(.a(s_163), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1692(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1693(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1694(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2073(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2074(.a(gate68inter0), .b(s_218), .O(gate68inter1));
  and2  gate2075(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2076(.a(s_218), .O(gate68inter3));
  inv1  gate2077(.a(s_219), .O(gate68inter4));
  nand2 gate2078(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2079(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2080(.a(G28), .O(gate68inter7));
  inv1  gate2081(.a(G305), .O(gate68inter8));
  nand2 gate2082(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2083(.a(s_219), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2084(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2085(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2086(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1961(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1962(.a(gate72inter0), .b(s_202), .O(gate72inter1));
  and2  gate1963(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1964(.a(s_202), .O(gate72inter3));
  inv1  gate1965(.a(s_203), .O(gate72inter4));
  nand2 gate1966(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1967(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1968(.a(G32), .O(gate72inter7));
  inv1  gate1969(.a(G311), .O(gate72inter8));
  nand2 gate1970(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1971(.a(s_203), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1972(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1973(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1974(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate645(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate646(.a(gate73inter0), .b(s_14), .O(gate73inter1));
  and2  gate647(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate648(.a(s_14), .O(gate73inter3));
  inv1  gate649(.a(s_15), .O(gate73inter4));
  nand2 gate650(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate651(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate652(.a(G1), .O(gate73inter7));
  inv1  gate653(.a(G314), .O(gate73inter8));
  nand2 gate654(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate655(.a(s_15), .b(gate73inter3), .O(gate73inter10));
  nor2  gate656(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate657(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate658(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1429(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1430(.a(gate81inter0), .b(s_126), .O(gate81inter1));
  and2  gate1431(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1432(.a(s_126), .O(gate81inter3));
  inv1  gate1433(.a(s_127), .O(gate81inter4));
  nand2 gate1434(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1435(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1436(.a(G3), .O(gate81inter7));
  inv1  gate1437(.a(G326), .O(gate81inter8));
  nand2 gate1438(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1439(.a(s_127), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1440(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1441(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1442(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1709(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1710(.a(gate82inter0), .b(s_166), .O(gate82inter1));
  and2  gate1711(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1712(.a(s_166), .O(gate82inter3));
  inv1  gate1713(.a(s_167), .O(gate82inter4));
  nand2 gate1714(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1715(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1716(.a(G7), .O(gate82inter7));
  inv1  gate1717(.a(G326), .O(gate82inter8));
  nand2 gate1718(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1719(.a(s_167), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1720(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1721(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1722(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2381(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2382(.a(gate83inter0), .b(s_262), .O(gate83inter1));
  and2  gate2383(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2384(.a(s_262), .O(gate83inter3));
  inv1  gate2385(.a(s_263), .O(gate83inter4));
  nand2 gate2386(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2387(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2388(.a(G11), .O(gate83inter7));
  inv1  gate2389(.a(G329), .O(gate83inter8));
  nand2 gate2390(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2391(.a(s_263), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2392(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2393(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2394(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2213(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2214(.a(gate86inter0), .b(s_238), .O(gate86inter1));
  and2  gate2215(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2216(.a(s_238), .O(gate86inter3));
  inv1  gate2217(.a(s_239), .O(gate86inter4));
  nand2 gate2218(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2219(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2220(.a(G8), .O(gate86inter7));
  inv1  gate2221(.a(G332), .O(gate86inter8));
  nand2 gate2222(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2223(.a(s_239), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2224(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2225(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2226(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1821(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1822(.a(gate89inter0), .b(s_182), .O(gate89inter1));
  and2  gate1823(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1824(.a(s_182), .O(gate89inter3));
  inv1  gate1825(.a(s_183), .O(gate89inter4));
  nand2 gate1826(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1827(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1828(.a(G17), .O(gate89inter7));
  inv1  gate1829(.a(G338), .O(gate89inter8));
  nand2 gate1830(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1831(.a(s_183), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1832(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1833(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1834(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1737(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1738(.a(gate97inter0), .b(s_170), .O(gate97inter1));
  and2  gate1739(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1740(.a(s_170), .O(gate97inter3));
  inv1  gate1741(.a(s_171), .O(gate97inter4));
  nand2 gate1742(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1743(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1744(.a(G19), .O(gate97inter7));
  inv1  gate1745(.a(G350), .O(gate97inter8));
  nand2 gate1746(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1747(.a(s_171), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1748(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1749(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1750(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1877(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1878(.a(gate98inter0), .b(s_190), .O(gate98inter1));
  and2  gate1879(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1880(.a(s_190), .O(gate98inter3));
  inv1  gate1881(.a(s_191), .O(gate98inter4));
  nand2 gate1882(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1883(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1884(.a(G23), .O(gate98inter7));
  inv1  gate1885(.a(G350), .O(gate98inter8));
  nand2 gate1886(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1887(.a(s_191), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1888(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1889(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1890(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1317(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1318(.a(gate101inter0), .b(s_110), .O(gate101inter1));
  and2  gate1319(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1320(.a(s_110), .O(gate101inter3));
  inv1  gate1321(.a(s_111), .O(gate101inter4));
  nand2 gate1322(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1323(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1324(.a(G20), .O(gate101inter7));
  inv1  gate1325(.a(G356), .O(gate101inter8));
  nand2 gate1326(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1327(.a(s_111), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1328(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1329(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1330(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate2465(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2466(.a(gate102inter0), .b(s_274), .O(gate102inter1));
  and2  gate2467(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2468(.a(s_274), .O(gate102inter3));
  inv1  gate2469(.a(s_275), .O(gate102inter4));
  nand2 gate2470(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2471(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2472(.a(G24), .O(gate102inter7));
  inv1  gate2473(.a(G356), .O(gate102inter8));
  nand2 gate2474(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2475(.a(s_275), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2476(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2477(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2478(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2269(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2270(.a(gate104inter0), .b(s_246), .O(gate104inter1));
  and2  gate2271(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2272(.a(s_246), .O(gate104inter3));
  inv1  gate2273(.a(s_247), .O(gate104inter4));
  nand2 gate2274(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2275(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2276(.a(G32), .O(gate104inter7));
  inv1  gate2277(.a(G359), .O(gate104inter8));
  nand2 gate2278(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2279(.a(s_247), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2280(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2281(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2282(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate2143(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2144(.a(gate105inter0), .b(s_228), .O(gate105inter1));
  and2  gate2145(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2146(.a(s_228), .O(gate105inter3));
  inv1  gate2147(.a(s_229), .O(gate105inter4));
  nand2 gate2148(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2149(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2150(.a(G362), .O(gate105inter7));
  inv1  gate2151(.a(G363), .O(gate105inter8));
  nand2 gate2152(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2153(.a(s_229), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2154(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2155(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2156(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate631(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate632(.a(gate106inter0), .b(s_12), .O(gate106inter1));
  and2  gate633(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate634(.a(s_12), .O(gate106inter3));
  inv1  gate635(.a(s_13), .O(gate106inter4));
  nand2 gate636(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate637(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate638(.a(G364), .O(gate106inter7));
  inv1  gate639(.a(G365), .O(gate106inter8));
  nand2 gate640(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate641(.a(s_13), .b(gate106inter3), .O(gate106inter10));
  nor2  gate642(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate643(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate644(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2437(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2438(.a(gate114inter0), .b(s_270), .O(gate114inter1));
  and2  gate2439(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2440(.a(s_270), .O(gate114inter3));
  inv1  gate2441(.a(s_271), .O(gate114inter4));
  nand2 gate2442(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2443(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2444(.a(G380), .O(gate114inter7));
  inv1  gate2445(.a(G381), .O(gate114inter8));
  nand2 gate2446(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2447(.a(s_271), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2448(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2449(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2450(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1219(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1220(.a(gate118inter0), .b(s_96), .O(gate118inter1));
  and2  gate1221(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1222(.a(s_96), .O(gate118inter3));
  inv1  gate1223(.a(s_97), .O(gate118inter4));
  nand2 gate1224(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1225(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1226(.a(G388), .O(gate118inter7));
  inv1  gate1227(.a(G389), .O(gate118inter8));
  nand2 gate1228(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1229(.a(s_97), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1230(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1231(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1232(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1513(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1514(.a(gate124inter0), .b(s_138), .O(gate124inter1));
  and2  gate1515(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1516(.a(s_138), .O(gate124inter3));
  inv1  gate1517(.a(s_139), .O(gate124inter4));
  nand2 gate1518(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1519(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1520(.a(G400), .O(gate124inter7));
  inv1  gate1521(.a(G401), .O(gate124inter8));
  nand2 gate1522(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1523(.a(s_139), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1524(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1525(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1526(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate2493(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2494(.a(gate125inter0), .b(s_278), .O(gate125inter1));
  and2  gate2495(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2496(.a(s_278), .O(gate125inter3));
  inv1  gate2497(.a(s_279), .O(gate125inter4));
  nand2 gate2498(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2499(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2500(.a(G402), .O(gate125inter7));
  inv1  gate2501(.a(G403), .O(gate125inter8));
  nand2 gate2502(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2503(.a(s_279), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2504(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2505(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2506(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate953(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate954(.a(gate126inter0), .b(s_58), .O(gate126inter1));
  and2  gate955(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate956(.a(s_58), .O(gate126inter3));
  inv1  gate957(.a(s_59), .O(gate126inter4));
  nand2 gate958(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate959(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate960(.a(G404), .O(gate126inter7));
  inv1  gate961(.a(G405), .O(gate126inter8));
  nand2 gate962(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate963(.a(s_59), .b(gate126inter3), .O(gate126inter10));
  nor2  gate964(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate965(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate966(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate659(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate660(.a(gate127inter0), .b(s_16), .O(gate127inter1));
  and2  gate661(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate662(.a(s_16), .O(gate127inter3));
  inv1  gate663(.a(s_17), .O(gate127inter4));
  nand2 gate664(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate665(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate666(.a(G406), .O(gate127inter7));
  inv1  gate667(.a(G407), .O(gate127inter8));
  nand2 gate668(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate669(.a(s_17), .b(gate127inter3), .O(gate127inter10));
  nor2  gate670(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate671(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate672(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1261(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1262(.a(gate130inter0), .b(s_102), .O(gate130inter1));
  and2  gate1263(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1264(.a(s_102), .O(gate130inter3));
  inv1  gate1265(.a(s_103), .O(gate130inter4));
  nand2 gate1266(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1267(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1268(.a(G412), .O(gate130inter7));
  inv1  gate1269(.a(G413), .O(gate130inter8));
  nand2 gate1270(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1271(.a(s_103), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1272(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1273(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1274(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2521(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2522(.a(gate134inter0), .b(s_282), .O(gate134inter1));
  and2  gate2523(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2524(.a(s_282), .O(gate134inter3));
  inv1  gate2525(.a(s_283), .O(gate134inter4));
  nand2 gate2526(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2527(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2528(.a(G420), .O(gate134inter7));
  inv1  gate2529(.a(G421), .O(gate134inter8));
  nand2 gate2530(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2531(.a(s_283), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2532(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2533(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2534(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1163(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1164(.a(gate137inter0), .b(s_88), .O(gate137inter1));
  and2  gate1165(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1166(.a(s_88), .O(gate137inter3));
  inv1  gate1167(.a(s_89), .O(gate137inter4));
  nand2 gate1168(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1169(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1170(.a(G426), .O(gate137inter7));
  inv1  gate1171(.a(G429), .O(gate137inter8));
  nand2 gate1172(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1173(.a(s_89), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1174(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1175(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1176(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate939(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate940(.a(gate139inter0), .b(s_56), .O(gate139inter1));
  and2  gate941(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate942(.a(s_56), .O(gate139inter3));
  inv1  gate943(.a(s_57), .O(gate139inter4));
  nand2 gate944(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate945(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate946(.a(G438), .O(gate139inter7));
  inv1  gate947(.a(G441), .O(gate139inter8));
  nand2 gate948(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate949(.a(s_57), .b(gate139inter3), .O(gate139inter10));
  nor2  gate950(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate951(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate952(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1093(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1094(.a(gate140inter0), .b(s_78), .O(gate140inter1));
  and2  gate1095(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1096(.a(s_78), .O(gate140inter3));
  inv1  gate1097(.a(s_79), .O(gate140inter4));
  nand2 gate1098(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1099(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1100(.a(G444), .O(gate140inter7));
  inv1  gate1101(.a(G447), .O(gate140inter8));
  nand2 gate1102(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1103(.a(s_79), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1104(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1105(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1106(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2395(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2396(.a(gate142inter0), .b(s_264), .O(gate142inter1));
  and2  gate2397(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2398(.a(s_264), .O(gate142inter3));
  inv1  gate2399(.a(s_265), .O(gate142inter4));
  nand2 gate2400(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2401(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2402(.a(G456), .O(gate142inter7));
  inv1  gate2403(.a(G459), .O(gate142inter8));
  nand2 gate2404(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2405(.a(s_265), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2406(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2407(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2408(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2283(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2284(.a(gate148inter0), .b(s_248), .O(gate148inter1));
  and2  gate2285(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2286(.a(s_248), .O(gate148inter3));
  inv1  gate2287(.a(s_249), .O(gate148inter4));
  nand2 gate2288(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2289(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2290(.a(G492), .O(gate148inter7));
  inv1  gate2291(.a(G495), .O(gate148inter8));
  nand2 gate2292(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2293(.a(s_249), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2294(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2295(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2296(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2297(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2298(.a(gate150inter0), .b(s_250), .O(gate150inter1));
  and2  gate2299(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2300(.a(s_250), .O(gate150inter3));
  inv1  gate2301(.a(s_251), .O(gate150inter4));
  nand2 gate2302(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2303(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2304(.a(G504), .O(gate150inter7));
  inv1  gate2305(.a(G507), .O(gate150inter8));
  nand2 gate2306(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2307(.a(s_251), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2308(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2309(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2310(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1121(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1122(.a(gate152inter0), .b(s_82), .O(gate152inter1));
  and2  gate1123(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1124(.a(s_82), .O(gate152inter3));
  inv1  gate1125(.a(s_83), .O(gate152inter4));
  nand2 gate1126(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1127(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1128(.a(G516), .O(gate152inter7));
  inv1  gate1129(.a(G519), .O(gate152inter8));
  nand2 gate1130(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1131(.a(s_83), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1132(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1133(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1134(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2591(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2592(.a(gate156inter0), .b(s_292), .O(gate156inter1));
  and2  gate2593(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2594(.a(s_292), .O(gate156inter3));
  inv1  gate2595(.a(s_293), .O(gate156inter4));
  nand2 gate2596(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2597(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2598(.a(G435), .O(gate156inter7));
  inv1  gate2599(.a(G525), .O(gate156inter8));
  nand2 gate2600(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2601(.a(s_293), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2602(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2603(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2604(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2367(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2368(.a(gate162inter0), .b(s_260), .O(gate162inter1));
  and2  gate2369(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2370(.a(s_260), .O(gate162inter3));
  inv1  gate2371(.a(s_261), .O(gate162inter4));
  nand2 gate2372(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2373(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2374(.a(G453), .O(gate162inter7));
  inv1  gate2375(.a(G534), .O(gate162inter8));
  nand2 gate2376(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2377(.a(s_261), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2378(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2379(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2380(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate911(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate912(.a(gate163inter0), .b(s_52), .O(gate163inter1));
  and2  gate913(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate914(.a(s_52), .O(gate163inter3));
  inv1  gate915(.a(s_53), .O(gate163inter4));
  nand2 gate916(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate917(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate918(.a(G456), .O(gate163inter7));
  inv1  gate919(.a(G537), .O(gate163inter8));
  nand2 gate920(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate921(.a(s_53), .b(gate163inter3), .O(gate163inter10));
  nor2  gate922(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate923(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate924(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2563(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2564(.a(gate164inter0), .b(s_288), .O(gate164inter1));
  and2  gate2565(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2566(.a(s_288), .O(gate164inter3));
  inv1  gate2567(.a(s_289), .O(gate164inter4));
  nand2 gate2568(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2569(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2570(.a(G459), .O(gate164inter7));
  inv1  gate2571(.a(G537), .O(gate164inter8));
  nand2 gate2572(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2573(.a(s_289), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2574(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2575(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2576(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate869(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate870(.a(gate167inter0), .b(s_46), .O(gate167inter1));
  and2  gate871(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate872(.a(s_46), .O(gate167inter3));
  inv1  gate873(.a(s_47), .O(gate167inter4));
  nand2 gate874(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate875(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate876(.a(G468), .O(gate167inter7));
  inv1  gate877(.a(G543), .O(gate167inter8));
  nand2 gate878(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate879(.a(s_47), .b(gate167inter3), .O(gate167inter10));
  nor2  gate880(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate881(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate882(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2045(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2046(.a(gate170inter0), .b(s_214), .O(gate170inter1));
  and2  gate2047(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2048(.a(s_214), .O(gate170inter3));
  inv1  gate2049(.a(s_215), .O(gate170inter4));
  nand2 gate2050(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2051(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2052(.a(G477), .O(gate170inter7));
  inv1  gate2053(.a(G546), .O(gate170inter8));
  nand2 gate2054(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2055(.a(s_215), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2056(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2057(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2058(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1051(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1052(.a(gate172inter0), .b(s_72), .O(gate172inter1));
  and2  gate1053(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1054(.a(s_72), .O(gate172inter3));
  inv1  gate1055(.a(s_73), .O(gate172inter4));
  nand2 gate1056(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1057(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1058(.a(G483), .O(gate172inter7));
  inv1  gate1059(.a(G549), .O(gate172inter8));
  nand2 gate1060(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1061(.a(s_73), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1062(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1063(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1064(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1331(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1332(.a(gate178inter0), .b(s_112), .O(gate178inter1));
  and2  gate1333(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1334(.a(s_112), .O(gate178inter3));
  inv1  gate1335(.a(s_113), .O(gate178inter4));
  nand2 gate1336(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1337(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1338(.a(G501), .O(gate178inter7));
  inv1  gate1339(.a(G558), .O(gate178inter8));
  nand2 gate1340(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1341(.a(s_113), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1342(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1343(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1344(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate925(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate926(.a(gate180inter0), .b(s_54), .O(gate180inter1));
  and2  gate927(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate928(.a(s_54), .O(gate180inter3));
  inv1  gate929(.a(s_55), .O(gate180inter4));
  nand2 gate930(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate931(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate932(.a(G507), .O(gate180inter7));
  inv1  gate933(.a(G561), .O(gate180inter8));
  nand2 gate934(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate935(.a(s_55), .b(gate180inter3), .O(gate180inter10));
  nor2  gate936(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate937(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate938(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate2409(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2410(.a(gate181inter0), .b(s_266), .O(gate181inter1));
  and2  gate2411(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2412(.a(s_266), .O(gate181inter3));
  inv1  gate2413(.a(s_267), .O(gate181inter4));
  nand2 gate2414(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2415(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2416(.a(G510), .O(gate181inter7));
  inv1  gate2417(.a(G564), .O(gate181inter8));
  nand2 gate2418(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2419(.a(s_267), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2420(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2421(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2422(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1457(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1458(.a(gate185inter0), .b(s_130), .O(gate185inter1));
  and2  gate1459(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1460(.a(s_130), .O(gate185inter3));
  inv1  gate1461(.a(s_131), .O(gate185inter4));
  nand2 gate1462(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1463(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1464(.a(G570), .O(gate185inter7));
  inv1  gate1465(.a(G571), .O(gate185inter8));
  nand2 gate1466(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1467(.a(s_131), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1468(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1469(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1470(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate715(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate716(.a(gate186inter0), .b(s_24), .O(gate186inter1));
  and2  gate717(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate718(.a(s_24), .O(gate186inter3));
  inv1  gate719(.a(s_25), .O(gate186inter4));
  nand2 gate720(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate721(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate722(.a(G572), .O(gate186inter7));
  inv1  gate723(.a(G573), .O(gate186inter8));
  nand2 gate724(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate725(.a(s_25), .b(gate186inter3), .O(gate186inter10));
  nor2  gate726(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate727(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate728(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2647(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2648(.a(gate188inter0), .b(s_300), .O(gate188inter1));
  and2  gate2649(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2650(.a(s_300), .O(gate188inter3));
  inv1  gate2651(.a(s_301), .O(gate188inter4));
  nand2 gate2652(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2653(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2654(.a(G576), .O(gate188inter7));
  inv1  gate2655(.a(G577), .O(gate188inter8));
  nand2 gate2656(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2657(.a(s_301), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2658(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2659(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2660(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2115(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2116(.a(gate189inter0), .b(s_224), .O(gate189inter1));
  and2  gate2117(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2118(.a(s_224), .O(gate189inter3));
  inv1  gate2119(.a(s_225), .O(gate189inter4));
  nand2 gate2120(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2121(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2122(.a(G578), .O(gate189inter7));
  inv1  gate2123(.a(G579), .O(gate189inter8));
  nand2 gate2124(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2125(.a(s_225), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2126(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2127(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2128(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate799(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate800(.a(gate190inter0), .b(s_36), .O(gate190inter1));
  and2  gate801(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate802(.a(s_36), .O(gate190inter3));
  inv1  gate803(.a(s_37), .O(gate190inter4));
  nand2 gate804(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate805(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate806(.a(G580), .O(gate190inter7));
  inv1  gate807(.a(G581), .O(gate190inter8));
  nand2 gate808(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate809(.a(s_37), .b(gate190inter3), .O(gate190inter10));
  nor2  gate810(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate811(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate812(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate743(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate744(.a(gate194inter0), .b(s_28), .O(gate194inter1));
  and2  gate745(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate746(.a(s_28), .O(gate194inter3));
  inv1  gate747(.a(s_29), .O(gate194inter4));
  nand2 gate748(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate749(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate750(.a(G588), .O(gate194inter7));
  inv1  gate751(.a(G589), .O(gate194inter8));
  nand2 gate752(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate753(.a(s_29), .b(gate194inter3), .O(gate194inter10));
  nor2  gate754(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate755(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate756(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1191(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1192(.a(gate197inter0), .b(s_92), .O(gate197inter1));
  and2  gate1193(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1194(.a(s_92), .O(gate197inter3));
  inv1  gate1195(.a(s_93), .O(gate197inter4));
  nand2 gate1196(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1197(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1198(.a(G594), .O(gate197inter7));
  inv1  gate1199(.a(G595), .O(gate197inter8));
  nand2 gate1200(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1201(.a(s_93), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1202(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1203(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1204(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1079(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1080(.a(gate198inter0), .b(s_76), .O(gate198inter1));
  and2  gate1081(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1082(.a(s_76), .O(gate198inter3));
  inv1  gate1083(.a(s_77), .O(gate198inter4));
  nand2 gate1084(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1085(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1086(.a(G596), .O(gate198inter7));
  inv1  gate1087(.a(G597), .O(gate198inter8));
  nand2 gate1088(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1089(.a(s_77), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1090(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1091(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1092(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate2325(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate2326(.a(gate201inter0), .b(s_254), .O(gate201inter1));
  and2  gate2327(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate2328(.a(s_254), .O(gate201inter3));
  inv1  gate2329(.a(s_255), .O(gate201inter4));
  nand2 gate2330(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2331(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2332(.a(G602), .O(gate201inter7));
  inv1  gate2333(.a(G607), .O(gate201inter8));
  nand2 gate2334(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2335(.a(s_255), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2336(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2337(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2338(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate2507(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2508(.a(gate202inter0), .b(s_280), .O(gate202inter1));
  and2  gate2509(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2510(.a(s_280), .O(gate202inter3));
  inv1  gate2511(.a(s_281), .O(gate202inter4));
  nand2 gate2512(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2513(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2514(.a(G612), .O(gate202inter7));
  inv1  gate2515(.a(G617), .O(gate202inter8));
  nand2 gate2516(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2517(.a(s_281), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2518(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2519(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2520(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2199(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2200(.a(gate205inter0), .b(s_236), .O(gate205inter1));
  and2  gate2201(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2202(.a(s_236), .O(gate205inter3));
  inv1  gate2203(.a(s_237), .O(gate205inter4));
  nand2 gate2204(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2205(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2206(.a(G622), .O(gate205inter7));
  inv1  gate2207(.a(G627), .O(gate205inter8));
  nand2 gate2208(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2209(.a(s_237), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2210(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2211(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2212(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate729(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate730(.a(gate208inter0), .b(s_26), .O(gate208inter1));
  and2  gate731(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate732(.a(s_26), .O(gate208inter3));
  inv1  gate733(.a(s_27), .O(gate208inter4));
  nand2 gate734(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate735(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate736(.a(G627), .O(gate208inter7));
  inv1  gate737(.a(G637), .O(gate208inter8));
  nand2 gate738(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate739(.a(s_27), .b(gate208inter3), .O(gate208inter10));
  nor2  gate740(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate741(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate742(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate2003(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2004(.a(gate209inter0), .b(s_208), .O(gate209inter1));
  and2  gate2005(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2006(.a(s_208), .O(gate209inter3));
  inv1  gate2007(.a(s_209), .O(gate209inter4));
  nand2 gate2008(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2009(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2010(.a(G602), .O(gate209inter7));
  inv1  gate2011(.a(G666), .O(gate209inter8));
  nand2 gate2012(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2013(.a(s_209), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2014(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2015(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2016(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1905(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1906(.a(gate210inter0), .b(s_194), .O(gate210inter1));
  and2  gate1907(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1908(.a(s_194), .O(gate210inter3));
  inv1  gate1909(.a(s_195), .O(gate210inter4));
  nand2 gate1910(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1911(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1912(.a(G607), .O(gate210inter7));
  inv1  gate1913(.a(G666), .O(gate210inter8));
  nand2 gate1914(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1915(.a(s_195), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1916(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1917(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1918(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2311(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2312(.a(gate212inter0), .b(s_252), .O(gate212inter1));
  and2  gate2313(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2314(.a(s_252), .O(gate212inter3));
  inv1  gate2315(.a(s_253), .O(gate212inter4));
  nand2 gate2316(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2317(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2318(.a(G617), .O(gate212inter7));
  inv1  gate2319(.a(G669), .O(gate212inter8));
  nand2 gate2320(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2321(.a(s_253), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2322(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2323(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2324(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate2185(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2186(.a(gate213inter0), .b(s_234), .O(gate213inter1));
  and2  gate2187(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2188(.a(s_234), .O(gate213inter3));
  inv1  gate2189(.a(s_235), .O(gate213inter4));
  nand2 gate2190(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2191(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2192(.a(G602), .O(gate213inter7));
  inv1  gate2193(.a(G672), .O(gate213inter8));
  nand2 gate2194(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2195(.a(s_235), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2196(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2197(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2198(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate603(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate604(.a(gate220inter0), .b(s_8), .O(gate220inter1));
  and2  gate605(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate606(.a(s_8), .O(gate220inter3));
  inv1  gate607(.a(s_9), .O(gate220inter4));
  nand2 gate608(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate609(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate610(.a(G637), .O(gate220inter7));
  inv1  gate611(.a(G681), .O(gate220inter8));
  nand2 gate612(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate613(.a(s_9), .b(gate220inter3), .O(gate220inter10));
  nor2  gate614(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate615(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate616(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1597(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1598(.a(gate222inter0), .b(s_150), .O(gate222inter1));
  and2  gate1599(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1600(.a(s_150), .O(gate222inter3));
  inv1  gate1601(.a(s_151), .O(gate222inter4));
  nand2 gate1602(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1603(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1604(.a(G632), .O(gate222inter7));
  inv1  gate1605(.a(G684), .O(gate222inter8));
  nand2 gate1606(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1607(.a(s_151), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1608(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1609(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1610(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1009(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1010(.a(gate223inter0), .b(s_66), .O(gate223inter1));
  and2  gate1011(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1012(.a(s_66), .O(gate223inter3));
  inv1  gate1013(.a(s_67), .O(gate223inter4));
  nand2 gate1014(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1015(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1016(.a(G627), .O(gate223inter7));
  inv1  gate1017(.a(G687), .O(gate223inter8));
  nand2 gate1018(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1019(.a(s_67), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1020(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1021(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1022(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate981(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate982(.a(gate224inter0), .b(s_62), .O(gate224inter1));
  and2  gate983(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate984(.a(s_62), .O(gate224inter3));
  inv1  gate985(.a(s_63), .O(gate224inter4));
  nand2 gate986(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate987(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate988(.a(G637), .O(gate224inter7));
  inv1  gate989(.a(G687), .O(gate224inter8));
  nand2 gate990(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate991(.a(s_63), .b(gate224inter3), .O(gate224inter10));
  nor2  gate992(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate993(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate994(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1107(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1108(.a(gate226inter0), .b(s_80), .O(gate226inter1));
  and2  gate1109(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1110(.a(s_80), .O(gate226inter3));
  inv1  gate1111(.a(s_81), .O(gate226inter4));
  nand2 gate1112(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1113(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1114(.a(G692), .O(gate226inter7));
  inv1  gate1115(.a(G693), .O(gate226inter8));
  nand2 gate1116(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1117(.a(s_81), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1118(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1119(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1120(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1037(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1038(.a(gate228inter0), .b(s_70), .O(gate228inter1));
  and2  gate1039(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1040(.a(s_70), .O(gate228inter3));
  inv1  gate1041(.a(s_71), .O(gate228inter4));
  nand2 gate1042(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1043(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1044(.a(G696), .O(gate228inter7));
  inv1  gate1045(.a(G697), .O(gate228inter8));
  nand2 gate1046(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1047(.a(s_71), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1048(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1049(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1050(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2171(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2172(.a(gate229inter0), .b(s_232), .O(gate229inter1));
  and2  gate2173(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2174(.a(s_232), .O(gate229inter3));
  inv1  gate2175(.a(s_233), .O(gate229inter4));
  nand2 gate2176(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2177(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2178(.a(G698), .O(gate229inter7));
  inv1  gate2179(.a(G699), .O(gate229inter8));
  nand2 gate2180(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2181(.a(s_233), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2182(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2183(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2184(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate2423(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2424(.a(gate232inter0), .b(s_268), .O(gate232inter1));
  and2  gate2425(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2426(.a(s_268), .O(gate232inter3));
  inv1  gate2427(.a(s_269), .O(gate232inter4));
  nand2 gate2428(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2429(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2430(.a(G704), .O(gate232inter7));
  inv1  gate2431(.a(G705), .O(gate232inter8));
  nand2 gate2432(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2433(.a(s_269), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2434(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2435(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2436(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1653(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1654(.a(gate233inter0), .b(s_158), .O(gate233inter1));
  and2  gate1655(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1656(.a(s_158), .O(gate233inter3));
  inv1  gate1657(.a(s_159), .O(gate233inter4));
  nand2 gate1658(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1659(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1660(.a(G242), .O(gate233inter7));
  inv1  gate1661(.a(G718), .O(gate233inter8));
  nand2 gate1662(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1663(.a(s_159), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1664(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1665(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1666(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate897(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate898(.a(gate235inter0), .b(s_50), .O(gate235inter1));
  and2  gate899(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate900(.a(s_50), .O(gate235inter3));
  inv1  gate901(.a(s_51), .O(gate235inter4));
  nand2 gate902(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate903(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate904(.a(G248), .O(gate235inter7));
  inv1  gate905(.a(G724), .O(gate235inter8));
  nand2 gate906(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate907(.a(s_51), .b(gate235inter3), .O(gate235inter10));
  nor2  gate908(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate909(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate910(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2339(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2340(.a(gate236inter0), .b(s_256), .O(gate236inter1));
  and2  gate2341(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2342(.a(s_256), .O(gate236inter3));
  inv1  gate2343(.a(s_257), .O(gate236inter4));
  nand2 gate2344(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2345(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2346(.a(G251), .O(gate236inter7));
  inv1  gate2347(.a(G727), .O(gate236inter8));
  nand2 gate2348(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2349(.a(s_257), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2350(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2351(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2352(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1667(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1668(.a(gate238inter0), .b(s_160), .O(gate238inter1));
  and2  gate1669(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1670(.a(s_160), .O(gate238inter3));
  inv1  gate1671(.a(s_161), .O(gate238inter4));
  nand2 gate1672(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1673(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1674(.a(G257), .O(gate238inter7));
  inv1  gate1675(.a(G709), .O(gate238inter8));
  nand2 gate1676(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1677(.a(s_161), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1678(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1679(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1680(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1205(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1206(.a(gate240inter0), .b(s_94), .O(gate240inter1));
  and2  gate1207(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1208(.a(s_94), .O(gate240inter3));
  inv1  gate1209(.a(s_95), .O(gate240inter4));
  nand2 gate1210(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1211(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1212(.a(G263), .O(gate240inter7));
  inv1  gate1213(.a(G715), .O(gate240inter8));
  nand2 gate1214(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1215(.a(s_95), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1216(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1217(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1218(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate575(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate576(.a(gate244inter0), .b(s_4), .O(gate244inter1));
  and2  gate577(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate578(.a(s_4), .O(gate244inter3));
  inv1  gate579(.a(s_5), .O(gate244inter4));
  nand2 gate580(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate581(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate582(.a(G721), .O(gate244inter7));
  inv1  gate583(.a(G733), .O(gate244inter8));
  nand2 gate584(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate585(.a(s_5), .b(gate244inter3), .O(gate244inter10));
  nor2  gate586(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate587(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate588(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1289(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1290(.a(gate246inter0), .b(s_106), .O(gate246inter1));
  and2  gate1291(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1292(.a(s_106), .O(gate246inter3));
  inv1  gate1293(.a(s_107), .O(gate246inter4));
  nand2 gate1294(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1295(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1296(.a(G724), .O(gate246inter7));
  inv1  gate1297(.a(G736), .O(gate246inter8));
  nand2 gate1298(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1299(.a(s_107), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1300(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1301(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1302(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate2017(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2018(.a(gate247inter0), .b(s_210), .O(gate247inter1));
  and2  gate2019(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2020(.a(s_210), .O(gate247inter3));
  inv1  gate2021(.a(s_211), .O(gate247inter4));
  nand2 gate2022(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2023(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2024(.a(G251), .O(gate247inter7));
  inv1  gate2025(.a(G739), .O(gate247inter8));
  nand2 gate2026(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2027(.a(s_211), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2028(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2029(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2030(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate687(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate688(.a(gate248inter0), .b(s_20), .O(gate248inter1));
  and2  gate689(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate690(.a(s_20), .O(gate248inter3));
  inv1  gate691(.a(s_21), .O(gate248inter4));
  nand2 gate692(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate693(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate694(.a(G727), .O(gate248inter7));
  inv1  gate695(.a(G739), .O(gate248inter8));
  nand2 gate696(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate697(.a(s_21), .b(gate248inter3), .O(gate248inter10));
  nor2  gate698(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate699(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate700(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2577(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2578(.a(gate249inter0), .b(s_290), .O(gate249inter1));
  and2  gate2579(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2580(.a(s_290), .O(gate249inter3));
  inv1  gate2581(.a(s_291), .O(gate249inter4));
  nand2 gate2582(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2583(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2584(.a(G254), .O(gate249inter7));
  inv1  gate2585(.a(G742), .O(gate249inter8));
  nand2 gate2586(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2587(.a(s_291), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2588(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2589(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2590(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1373(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1374(.a(gate252inter0), .b(s_118), .O(gate252inter1));
  and2  gate1375(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1376(.a(s_118), .O(gate252inter3));
  inv1  gate1377(.a(s_119), .O(gate252inter4));
  nand2 gate1378(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1379(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1380(.a(G709), .O(gate252inter7));
  inv1  gate1381(.a(G745), .O(gate252inter8));
  nand2 gate1382(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1383(.a(s_119), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1384(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1385(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1386(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate617(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate618(.a(gate256inter0), .b(s_10), .O(gate256inter1));
  and2  gate619(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate620(.a(s_10), .O(gate256inter3));
  inv1  gate621(.a(s_11), .O(gate256inter4));
  nand2 gate622(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate623(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate624(.a(G715), .O(gate256inter7));
  inv1  gate625(.a(G751), .O(gate256inter8));
  nand2 gate626(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate627(.a(s_11), .b(gate256inter3), .O(gate256inter10));
  nor2  gate628(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate629(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate630(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1723(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1724(.a(gate260inter0), .b(s_168), .O(gate260inter1));
  and2  gate1725(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1726(.a(s_168), .O(gate260inter3));
  inv1  gate1727(.a(s_169), .O(gate260inter4));
  nand2 gate1728(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1729(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1730(.a(G760), .O(gate260inter7));
  inv1  gate1731(.a(G761), .O(gate260inter8));
  nand2 gate1732(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1733(.a(s_169), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1734(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1735(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1736(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1387(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1388(.a(gate261inter0), .b(s_120), .O(gate261inter1));
  and2  gate1389(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1390(.a(s_120), .O(gate261inter3));
  inv1  gate1391(.a(s_121), .O(gate261inter4));
  nand2 gate1392(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1393(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1394(.a(G762), .O(gate261inter7));
  inv1  gate1395(.a(G763), .O(gate261inter8));
  nand2 gate1396(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1397(.a(s_121), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1398(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1399(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1400(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate813(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate814(.a(gate262inter0), .b(s_38), .O(gate262inter1));
  and2  gate815(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate816(.a(s_38), .O(gate262inter3));
  inv1  gate817(.a(s_39), .O(gate262inter4));
  nand2 gate818(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate819(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate820(.a(G764), .O(gate262inter7));
  inv1  gate821(.a(G765), .O(gate262inter8));
  nand2 gate822(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate823(.a(s_39), .b(gate262inter3), .O(gate262inter10));
  nor2  gate824(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate825(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate826(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1611(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1612(.a(gate264inter0), .b(s_152), .O(gate264inter1));
  and2  gate1613(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1614(.a(s_152), .O(gate264inter3));
  inv1  gate1615(.a(s_153), .O(gate264inter4));
  nand2 gate1616(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1617(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1618(.a(G768), .O(gate264inter7));
  inv1  gate1619(.a(G769), .O(gate264inter8));
  nand2 gate1620(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1621(.a(s_153), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1622(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1623(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1624(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate771(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate772(.a(gate268inter0), .b(s_32), .O(gate268inter1));
  and2  gate773(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate774(.a(s_32), .O(gate268inter3));
  inv1  gate775(.a(s_33), .O(gate268inter4));
  nand2 gate776(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate777(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate778(.a(G651), .O(gate268inter7));
  inv1  gate779(.a(G779), .O(gate268inter8));
  nand2 gate780(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate781(.a(s_33), .b(gate268inter3), .O(gate268inter10));
  nor2  gate782(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate783(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate784(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1779(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1780(.a(gate270inter0), .b(s_176), .O(gate270inter1));
  and2  gate1781(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1782(.a(s_176), .O(gate270inter3));
  inv1  gate1783(.a(s_177), .O(gate270inter4));
  nand2 gate1784(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1785(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1786(.a(G657), .O(gate270inter7));
  inv1  gate1787(.a(G785), .O(gate270inter8));
  nand2 gate1788(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1789(.a(s_177), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1790(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1791(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1792(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1499(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1500(.a(gate271inter0), .b(s_136), .O(gate271inter1));
  and2  gate1501(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1502(.a(s_136), .O(gate271inter3));
  inv1  gate1503(.a(s_137), .O(gate271inter4));
  nand2 gate1504(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1505(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1506(.a(G660), .O(gate271inter7));
  inv1  gate1507(.a(G788), .O(gate271inter8));
  nand2 gate1508(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1509(.a(s_137), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1510(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1511(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1512(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate841(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate842(.a(gate273inter0), .b(s_42), .O(gate273inter1));
  and2  gate843(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate844(.a(s_42), .O(gate273inter3));
  inv1  gate845(.a(s_43), .O(gate273inter4));
  nand2 gate846(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate847(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate848(.a(G642), .O(gate273inter7));
  inv1  gate849(.a(G794), .O(gate273inter8));
  nand2 gate850(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate851(.a(s_43), .b(gate273inter3), .O(gate273inter10));
  nor2  gate852(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate853(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate854(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1415(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1416(.a(gate275inter0), .b(s_124), .O(gate275inter1));
  and2  gate1417(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1418(.a(s_124), .O(gate275inter3));
  inv1  gate1419(.a(s_125), .O(gate275inter4));
  nand2 gate1420(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1421(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1422(.a(G645), .O(gate275inter7));
  inv1  gate1423(.a(G797), .O(gate275inter8));
  nand2 gate1424(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1425(.a(s_125), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1426(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1427(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1428(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1807(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1808(.a(gate282inter0), .b(s_180), .O(gate282inter1));
  and2  gate1809(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1810(.a(s_180), .O(gate282inter3));
  inv1  gate1811(.a(s_181), .O(gate282inter4));
  nand2 gate1812(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1813(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1814(.a(G782), .O(gate282inter7));
  inv1  gate1815(.a(G806), .O(gate282inter8));
  nand2 gate1816(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1817(.a(s_181), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1818(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1819(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1820(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2101(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2102(.a(gate283inter0), .b(s_222), .O(gate283inter1));
  and2  gate2103(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2104(.a(s_222), .O(gate283inter3));
  inv1  gate2105(.a(s_223), .O(gate283inter4));
  nand2 gate2106(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2107(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2108(.a(G657), .O(gate283inter7));
  inv1  gate2109(.a(G809), .O(gate283inter8));
  nand2 gate2110(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2111(.a(s_223), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2112(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2113(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2114(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate757(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate758(.a(gate286inter0), .b(s_30), .O(gate286inter1));
  and2  gate759(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate760(.a(s_30), .O(gate286inter3));
  inv1  gate761(.a(s_31), .O(gate286inter4));
  nand2 gate762(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate763(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate764(.a(G788), .O(gate286inter7));
  inv1  gate765(.a(G812), .O(gate286inter8));
  nand2 gate766(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate767(.a(s_31), .b(gate286inter3), .O(gate286inter10));
  nor2  gate768(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate769(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate770(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2031(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2032(.a(gate288inter0), .b(s_212), .O(gate288inter1));
  and2  gate2033(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2034(.a(s_212), .O(gate288inter3));
  inv1  gate2035(.a(s_213), .O(gate288inter4));
  nand2 gate2036(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2037(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2038(.a(G791), .O(gate288inter7));
  inv1  gate2039(.a(G815), .O(gate288inter8));
  nand2 gate2040(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2041(.a(s_213), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2042(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2043(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2044(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1793(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1794(.a(gate290inter0), .b(s_178), .O(gate290inter1));
  and2  gate1795(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1796(.a(s_178), .O(gate290inter3));
  inv1  gate1797(.a(s_179), .O(gate290inter4));
  nand2 gate1798(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1799(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1800(.a(G820), .O(gate290inter7));
  inv1  gate1801(.a(G821), .O(gate290inter8));
  nand2 gate1802(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1803(.a(s_179), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1804(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1805(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1806(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1135(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1136(.a(gate294inter0), .b(s_84), .O(gate294inter1));
  and2  gate1137(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1138(.a(s_84), .O(gate294inter3));
  inv1  gate1139(.a(s_85), .O(gate294inter4));
  nand2 gate1140(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1141(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1142(.a(G832), .O(gate294inter7));
  inv1  gate1143(.a(G833), .O(gate294inter8));
  nand2 gate1144(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1145(.a(s_85), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1146(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1147(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1148(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1065(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1066(.a(gate389inter0), .b(s_74), .O(gate389inter1));
  and2  gate1067(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1068(.a(s_74), .O(gate389inter3));
  inv1  gate1069(.a(s_75), .O(gate389inter4));
  nand2 gate1070(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1071(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1072(.a(G3), .O(gate389inter7));
  inv1  gate1073(.a(G1042), .O(gate389inter8));
  nand2 gate1074(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1075(.a(s_75), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1076(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1077(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1078(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1149(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1150(.a(gate399inter0), .b(s_86), .O(gate399inter1));
  and2  gate1151(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1152(.a(s_86), .O(gate399inter3));
  inv1  gate1153(.a(s_87), .O(gate399inter4));
  nand2 gate1154(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1155(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1156(.a(G13), .O(gate399inter7));
  inv1  gate1157(.a(G1072), .O(gate399inter8));
  nand2 gate1158(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1159(.a(s_87), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1160(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1161(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1162(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate855(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate856(.a(gate402inter0), .b(s_44), .O(gate402inter1));
  and2  gate857(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate858(.a(s_44), .O(gate402inter3));
  inv1  gate859(.a(s_45), .O(gate402inter4));
  nand2 gate860(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate861(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate862(.a(G16), .O(gate402inter7));
  inv1  gate863(.a(G1081), .O(gate402inter8));
  nand2 gate864(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate865(.a(s_45), .b(gate402inter3), .O(gate402inter10));
  nor2  gate866(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate867(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate868(.a(gate402inter12), .b(gate402inter1), .O(G1177));

  xor2  gate1401(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1402(.a(gate403inter0), .b(s_122), .O(gate403inter1));
  and2  gate1403(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1404(.a(s_122), .O(gate403inter3));
  inv1  gate1405(.a(s_123), .O(gate403inter4));
  nand2 gate1406(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1407(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1408(.a(G17), .O(gate403inter7));
  inv1  gate1409(.a(G1084), .O(gate403inter8));
  nand2 gate1410(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1411(.a(s_123), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1412(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1413(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1414(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate1471(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1472(.a(gate404inter0), .b(s_132), .O(gate404inter1));
  and2  gate1473(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1474(.a(s_132), .O(gate404inter3));
  inv1  gate1475(.a(s_133), .O(gate404inter4));
  nand2 gate1476(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1477(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1478(.a(G18), .O(gate404inter7));
  inv1  gate1479(.a(G1087), .O(gate404inter8));
  nand2 gate1480(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1481(.a(s_133), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1482(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1483(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1484(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1751(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1752(.a(gate406inter0), .b(s_172), .O(gate406inter1));
  and2  gate1753(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1754(.a(s_172), .O(gate406inter3));
  inv1  gate1755(.a(s_173), .O(gate406inter4));
  nand2 gate1756(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1757(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1758(.a(G20), .O(gate406inter7));
  inv1  gate1759(.a(G1093), .O(gate406inter8));
  nand2 gate1760(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1761(.a(s_173), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1762(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1763(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1764(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1891(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1892(.a(gate407inter0), .b(s_192), .O(gate407inter1));
  and2  gate1893(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1894(.a(s_192), .O(gate407inter3));
  inv1  gate1895(.a(s_193), .O(gate407inter4));
  nand2 gate1896(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1897(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1898(.a(G21), .O(gate407inter7));
  inv1  gate1899(.a(G1096), .O(gate407inter8));
  nand2 gate1900(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1901(.a(s_193), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1902(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1903(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1904(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1359(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1360(.a(gate410inter0), .b(s_116), .O(gate410inter1));
  and2  gate1361(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1362(.a(s_116), .O(gate410inter3));
  inv1  gate1363(.a(s_117), .O(gate410inter4));
  nand2 gate1364(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1365(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1366(.a(G24), .O(gate410inter7));
  inv1  gate1367(.a(G1105), .O(gate410inter8));
  nand2 gate1368(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1369(.a(s_117), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1370(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1371(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1372(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1345(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1346(.a(gate412inter0), .b(s_114), .O(gate412inter1));
  and2  gate1347(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1348(.a(s_114), .O(gate412inter3));
  inv1  gate1349(.a(s_115), .O(gate412inter4));
  nand2 gate1350(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1351(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1352(.a(G26), .O(gate412inter7));
  inv1  gate1353(.a(G1111), .O(gate412inter8));
  nand2 gate1354(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1355(.a(s_115), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1356(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1357(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1358(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1555(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1556(.a(gate419inter0), .b(s_144), .O(gate419inter1));
  and2  gate1557(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1558(.a(s_144), .O(gate419inter3));
  inv1  gate1559(.a(s_145), .O(gate419inter4));
  nand2 gate1560(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1561(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1562(.a(G1), .O(gate419inter7));
  inv1  gate1563(.a(G1132), .O(gate419inter8));
  nand2 gate1564(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1565(.a(s_145), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1566(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1567(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1568(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1583(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1584(.a(gate420inter0), .b(s_148), .O(gate420inter1));
  and2  gate1585(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1586(.a(s_148), .O(gate420inter3));
  inv1  gate1587(.a(s_149), .O(gate420inter4));
  nand2 gate1588(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1589(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1590(.a(G1036), .O(gate420inter7));
  inv1  gate1591(.a(G1132), .O(gate420inter8));
  nand2 gate1592(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1593(.a(s_149), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1594(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1595(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1596(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2129(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2130(.a(gate421inter0), .b(s_226), .O(gate421inter1));
  and2  gate2131(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2132(.a(s_226), .O(gate421inter3));
  inv1  gate2133(.a(s_227), .O(gate421inter4));
  nand2 gate2134(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2135(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2136(.a(G2), .O(gate421inter7));
  inv1  gate2137(.a(G1135), .O(gate421inter8));
  nand2 gate2138(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2139(.a(s_227), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2140(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2141(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2142(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate785(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate786(.a(gate422inter0), .b(s_34), .O(gate422inter1));
  and2  gate787(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate788(.a(s_34), .O(gate422inter3));
  inv1  gate789(.a(s_35), .O(gate422inter4));
  nand2 gate790(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate791(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate792(.a(G1039), .O(gate422inter7));
  inv1  gate793(.a(G1135), .O(gate422inter8));
  nand2 gate794(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate795(.a(s_35), .b(gate422inter3), .O(gate422inter10));
  nor2  gate796(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate797(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate798(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate547(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate548(.a(gate423inter0), .b(s_0), .O(gate423inter1));
  and2  gate549(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate550(.a(s_0), .O(gate423inter3));
  inv1  gate551(.a(s_1), .O(gate423inter4));
  nand2 gate552(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate553(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate554(.a(G3), .O(gate423inter7));
  inv1  gate555(.a(G1138), .O(gate423inter8));
  nand2 gate556(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate557(.a(s_1), .b(gate423inter3), .O(gate423inter10));
  nor2  gate558(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate559(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate560(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1303(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1304(.a(gate424inter0), .b(s_108), .O(gate424inter1));
  and2  gate1305(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1306(.a(s_108), .O(gate424inter3));
  inv1  gate1307(.a(s_109), .O(gate424inter4));
  nand2 gate1308(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1309(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1310(.a(G1042), .O(gate424inter7));
  inv1  gate1311(.a(G1138), .O(gate424inter8));
  nand2 gate1312(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1313(.a(s_109), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1314(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1315(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1316(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1569(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1570(.a(gate435inter0), .b(s_146), .O(gate435inter1));
  and2  gate1571(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1572(.a(s_146), .O(gate435inter3));
  inv1  gate1573(.a(s_147), .O(gate435inter4));
  nand2 gate1574(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1575(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1576(.a(G9), .O(gate435inter7));
  inv1  gate1577(.a(G1156), .O(gate435inter8));
  nand2 gate1578(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1579(.a(s_147), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1580(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1581(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1582(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate1947(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1948(.a(gate436inter0), .b(s_200), .O(gate436inter1));
  and2  gate1949(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1950(.a(s_200), .O(gate436inter3));
  inv1  gate1951(.a(s_201), .O(gate436inter4));
  nand2 gate1952(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1953(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1954(.a(G1060), .O(gate436inter7));
  inv1  gate1955(.a(G1156), .O(gate436inter8));
  nand2 gate1956(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1957(.a(s_201), .b(gate436inter3), .O(gate436inter10));
  nor2  gate1958(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate1959(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate1960(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate995(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate996(.a(gate439inter0), .b(s_64), .O(gate439inter1));
  and2  gate997(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate998(.a(s_64), .O(gate439inter3));
  inv1  gate999(.a(s_65), .O(gate439inter4));
  nand2 gate1000(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1001(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1002(.a(G11), .O(gate439inter7));
  inv1  gate1003(.a(G1162), .O(gate439inter8));
  nand2 gate1004(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1005(.a(s_65), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1006(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1007(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1008(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate1023(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1024(.a(gate440inter0), .b(s_68), .O(gate440inter1));
  and2  gate1025(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1026(.a(s_68), .O(gate440inter3));
  inv1  gate1027(.a(s_69), .O(gate440inter4));
  nand2 gate1028(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1029(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1030(.a(G1066), .O(gate440inter7));
  inv1  gate1031(.a(G1162), .O(gate440inter8));
  nand2 gate1032(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1033(.a(s_69), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1034(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1035(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1036(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1639(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1640(.a(gate441inter0), .b(s_156), .O(gate441inter1));
  and2  gate1641(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1642(.a(s_156), .O(gate441inter3));
  inv1  gate1643(.a(s_157), .O(gate441inter4));
  nand2 gate1644(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1645(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1646(.a(G12), .O(gate441inter7));
  inv1  gate1647(.a(G1165), .O(gate441inter8));
  nand2 gate1648(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1649(.a(s_157), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1650(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1651(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1652(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate2157(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate2158(.a(gate453inter0), .b(s_230), .O(gate453inter1));
  and2  gate2159(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate2160(.a(s_230), .O(gate453inter3));
  inv1  gate2161(.a(s_231), .O(gate453inter4));
  nand2 gate2162(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate2163(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate2164(.a(G18), .O(gate453inter7));
  inv1  gate2165(.a(G1183), .O(gate453inter8));
  nand2 gate2166(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate2167(.a(s_231), .b(gate453inter3), .O(gate453inter10));
  nor2  gate2168(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate2169(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate2170(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2479(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2480(.a(gate458inter0), .b(s_276), .O(gate458inter1));
  and2  gate2481(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2482(.a(s_276), .O(gate458inter3));
  inv1  gate2483(.a(s_277), .O(gate458inter4));
  nand2 gate2484(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2485(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2486(.a(G1093), .O(gate458inter7));
  inv1  gate2487(.a(G1189), .O(gate458inter8));
  nand2 gate2488(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2489(.a(s_277), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2490(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2491(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2492(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1177(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1178(.a(gate463inter0), .b(s_90), .O(gate463inter1));
  and2  gate1179(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1180(.a(s_90), .O(gate463inter3));
  inv1  gate1181(.a(s_91), .O(gate463inter4));
  nand2 gate1182(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1183(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1184(.a(G23), .O(gate463inter7));
  inv1  gate1185(.a(G1198), .O(gate463inter8));
  nand2 gate1186(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1187(.a(s_91), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1188(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1189(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1190(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate2535(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2536(.a(gate473inter0), .b(s_284), .O(gate473inter1));
  and2  gate2537(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2538(.a(s_284), .O(gate473inter3));
  inv1  gate2539(.a(s_285), .O(gate473inter4));
  nand2 gate2540(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2541(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2542(.a(G28), .O(gate473inter7));
  inv1  gate2543(.a(G1213), .O(gate473inter8));
  nand2 gate2544(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2545(.a(s_285), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2546(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2547(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2548(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate2633(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2634(.a(gate474inter0), .b(s_298), .O(gate474inter1));
  and2  gate2635(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2636(.a(s_298), .O(gate474inter3));
  inv1  gate2637(.a(s_299), .O(gate474inter4));
  nand2 gate2638(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2639(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2640(.a(G1117), .O(gate474inter7));
  inv1  gate2641(.a(G1213), .O(gate474inter8));
  nand2 gate2642(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2643(.a(s_299), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2644(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2645(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2646(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1247(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1248(.a(gate478inter0), .b(s_100), .O(gate478inter1));
  and2  gate1249(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1250(.a(s_100), .O(gate478inter3));
  inv1  gate1251(.a(s_101), .O(gate478inter4));
  nand2 gate1252(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1253(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1254(.a(G1123), .O(gate478inter7));
  inv1  gate1255(.a(G1219), .O(gate478inter8));
  nand2 gate1256(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1257(.a(s_101), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1258(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1259(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1260(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate2353(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2354(.a(gate481inter0), .b(s_258), .O(gate481inter1));
  and2  gate2355(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2356(.a(s_258), .O(gate481inter3));
  inv1  gate2357(.a(s_259), .O(gate481inter4));
  nand2 gate2358(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2359(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2360(.a(G32), .O(gate481inter7));
  inv1  gate2361(.a(G1225), .O(gate481inter8));
  nand2 gate2362(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2363(.a(s_259), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2364(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2365(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2366(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1835(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1836(.a(gate483inter0), .b(s_184), .O(gate483inter1));
  and2  gate1837(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1838(.a(s_184), .O(gate483inter3));
  inv1  gate1839(.a(s_185), .O(gate483inter4));
  nand2 gate1840(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1841(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1842(.a(G1228), .O(gate483inter7));
  inv1  gate1843(.a(G1229), .O(gate483inter8));
  nand2 gate1844(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1845(.a(s_185), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1846(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1847(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1848(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2451(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2452(.a(gate492inter0), .b(s_272), .O(gate492inter1));
  and2  gate2453(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2454(.a(s_272), .O(gate492inter3));
  inv1  gate2455(.a(s_273), .O(gate492inter4));
  nand2 gate2456(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2457(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2458(.a(G1246), .O(gate492inter7));
  inv1  gate2459(.a(G1247), .O(gate492inter8));
  nand2 gate2460(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2461(.a(s_273), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2462(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2463(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2464(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate561(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate562(.a(gate494inter0), .b(s_2), .O(gate494inter1));
  and2  gate563(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate564(.a(s_2), .O(gate494inter3));
  inv1  gate565(.a(s_3), .O(gate494inter4));
  nand2 gate566(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate567(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate568(.a(G1250), .O(gate494inter7));
  inv1  gate569(.a(G1251), .O(gate494inter8));
  nand2 gate570(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate571(.a(s_3), .b(gate494inter3), .O(gate494inter10));
  nor2  gate572(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate573(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate574(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2241(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2242(.a(gate497inter0), .b(s_242), .O(gate497inter1));
  and2  gate2243(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2244(.a(s_242), .O(gate497inter3));
  inv1  gate2245(.a(s_243), .O(gate497inter4));
  nand2 gate2246(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2247(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2248(.a(G1256), .O(gate497inter7));
  inv1  gate2249(.a(G1257), .O(gate497inter8));
  nand2 gate2250(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2251(.a(s_243), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2252(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2253(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2254(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1919(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1920(.a(gate502inter0), .b(s_196), .O(gate502inter1));
  and2  gate1921(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1922(.a(s_196), .O(gate502inter3));
  inv1  gate1923(.a(s_197), .O(gate502inter4));
  nand2 gate1924(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1925(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1926(.a(G1266), .O(gate502inter7));
  inv1  gate1927(.a(G1267), .O(gate502inter8));
  nand2 gate1928(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1929(.a(s_197), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1930(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1931(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1932(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1933(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1934(.a(gate504inter0), .b(s_198), .O(gate504inter1));
  and2  gate1935(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1936(.a(s_198), .O(gate504inter3));
  inv1  gate1937(.a(s_199), .O(gate504inter4));
  nand2 gate1938(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1939(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1940(.a(G1270), .O(gate504inter7));
  inv1  gate1941(.a(G1271), .O(gate504inter8));
  nand2 gate1942(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1943(.a(s_199), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1944(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1945(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1946(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate2255(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2256(.a(gate505inter0), .b(s_244), .O(gate505inter1));
  and2  gate2257(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2258(.a(s_244), .O(gate505inter3));
  inv1  gate2259(.a(s_245), .O(gate505inter4));
  nand2 gate2260(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2261(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2262(.a(G1272), .O(gate505inter7));
  inv1  gate2263(.a(G1273), .O(gate505inter8));
  nand2 gate2264(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2265(.a(s_245), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2266(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2267(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2268(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1275(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1276(.a(gate506inter0), .b(s_104), .O(gate506inter1));
  and2  gate1277(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1278(.a(s_104), .O(gate506inter3));
  inv1  gate1279(.a(s_105), .O(gate506inter4));
  nand2 gate1280(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1281(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1282(.a(G1274), .O(gate506inter7));
  inv1  gate1283(.a(G1275), .O(gate506inter8));
  nand2 gate1284(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1285(.a(s_105), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1286(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1287(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1288(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2619(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2620(.a(gate510inter0), .b(s_296), .O(gate510inter1));
  and2  gate2621(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2622(.a(s_296), .O(gate510inter3));
  inv1  gate2623(.a(s_297), .O(gate510inter4));
  nand2 gate2624(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2625(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2626(.a(G1282), .O(gate510inter7));
  inv1  gate2627(.a(G1283), .O(gate510inter8));
  nand2 gate2628(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2629(.a(s_297), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2630(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2631(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2632(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1541(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1542(.a(gate511inter0), .b(s_142), .O(gate511inter1));
  and2  gate1543(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1544(.a(s_142), .O(gate511inter3));
  inv1  gate1545(.a(s_143), .O(gate511inter4));
  nand2 gate1546(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1547(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1548(.a(G1284), .O(gate511inter7));
  inv1  gate1549(.a(G1285), .O(gate511inter8));
  nand2 gate1550(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1551(.a(s_143), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1552(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1553(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1554(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1695(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1696(.a(gate513inter0), .b(s_164), .O(gate513inter1));
  and2  gate1697(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1698(.a(s_164), .O(gate513inter3));
  inv1  gate1699(.a(s_165), .O(gate513inter4));
  nand2 gate1700(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1701(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1702(.a(G1288), .O(gate513inter7));
  inv1  gate1703(.a(G1289), .O(gate513inter8));
  nand2 gate1704(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1705(.a(s_165), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1706(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1707(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1708(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1233(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1234(.a(gate514inter0), .b(s_98), .O(gate514inter1));
  and2  gate1235(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1236(.a(s_98), .O(gate514inter3));
  inv1  gate1237(.a(s_99), .O(gate514inter4));
  nand2 gate1238(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1239(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1240(.a(G1290), .O(gate514inter7));
  inv1  gate1241(.a(G1291), .O(gate514inter8));
  nand2 gate1242(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1243(.a(s_99), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1244(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1245(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1246(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule