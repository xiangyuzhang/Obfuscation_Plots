module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate617(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate618(.a(gate11inter0), .b(s_10), .O(gate11inter1));
  and2  gate619(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate620(.a(s_10), .O(gate11inter3));
  inv1  gate621(.a(s_11), .O(gate11inter4));
  nand2 gate622(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate623(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate624(.a(G5), .O(gate11inter7));
  inv1  gate625(.a(G6), .O(gate11inter8));
  nand2 gate626(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate627(.a(s_11), .b(gate11inter3), .O(gate11inter10));
  nor2  gate628(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate629(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate630(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1793(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1794(.a(gate14inter0), .b(s_178), .O(gate14inter1));
  and2  gate1795(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1796(.a(s_178), .O(gate14inter3));
  inv1  gate1797(.a(s_179), .O(gate14inter4));
  nand2 gate1798(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1799(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1800(.a(G11), .O(gate14inter7));
  inv1  gate1801(.a(G12), .O(gate14inter8));
  nand2 gate1802(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1803(.a(s_179), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1804(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1805(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1806(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate897(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate898(.a(gate16inter0), .b(s_50), .O(gate16inter1));
  and2  gate899(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate900(.a(s_50), .O(gate16inter3));
  inv1  gate901(.a(s_51), .O(gate16inter4));
  nand2 gate902(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate903(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate904(.a(G15), .O(gate16inter7));
  inv1  gate905(.a(G16), .O(gate16inter8));
  nand2 gate906(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate907(.a(s_51), .b(gate16inter3), .O(gate16inter10));
  nor2  gate908(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate909(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate910(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2479(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2480(.a(gate20inter0), .b(s_276), .O(gate20inter1));
  and2  gate2481(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2482(.a(s_276), .O(gate20inter3));
  inv1  gate2483(.a(s_277), .O(gate20inter4));
  nand2 gate2484(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2485(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2486(.a(G23), .O(gate20inter7));
  inv1  gate2487(.a(G24), .O(gate20inter8));
  nand2 gate2488(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2489(.a(s_277), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2490(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2491(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2492(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate687(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate688(.a(gate22inter0), .b(s_20), .O(gate22inter1));
  and2  gate689(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate690(.a(s_20), .O(gate22inter3));
  inv1  gate691(.a(s_21), .O(gate22inter4));
  nand2 gate692(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate693(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate694(.a(G27), .O(gate22inter7));
  inv1  gate695(.a(G28), .O(gate22inter8));
  nand2 gate696(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate697(.a(s_21), .b(gate22inter3), .O(gate22inter10));
  nor2  gate698(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate699(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate700(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2073(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2074(.a(gate23inter0), .b(s_218), .O(gate23inter1));
  and2  gate2075(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2076(.a(s_218), .O(gate23inter3));
  inv1  gate2077(.a(s_219), .O(gate23inter4));
  nand2 gate2078(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2079(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2080(.a(G29), .O(gate23inter7));
  inv1  gate2081(.a(G30), .O(gate23inter8));
  nand2 gate2082(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2083(.a(s_219), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2084(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2085(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2086(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate743(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate744(.a(gate27inter0), .b(s_28), .O(gate27inter1));
  and2  gate745(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate746(.a(s_28), .O(gate27inter3));
  inv1  gate747(.a(s_29), .O(gate27inter4));
  nand2 gate748(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate749(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate750(.a(G2), .O(gate27inter7));
  inv1  gate751(.a(G6), .O(gate27inter8));
  nand2 gate752(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate753(.a(s_29), .b(gate27inter3), .O(gate27inter10));
  nor2  gate754(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate755(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate756(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1317(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1318(.a(gate28inter0), .b(s_110), .O(gate28inter1));
  and2  gate1319(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1320(.a(s_110), .O(gate28inter3));
  inv1  gate1321(.a(s_111), .O(gate28inter4));
  nand2 gate1322(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1323(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1324(.a(G10), .O(gate28inter7));
  inv1  gate1325(.a(G14), .O(gate28inter8));
  nand2 gate1326(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1327(.a(s_111), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1328(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1329(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1330(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate757(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate758(.a(gate33inter0), .b(s_30), .O(gate33inter1));
  and2  gate759(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate760(.a(s_30), .O(gate33inter3));
  inv1  gate761(.a(s_31), .O(gate33inter4));
  nand2 gate762(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate763(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate764(.a(G17), .O(gate33inter7));
  inv1  gate765(.a(G21), .O(gate33inter8));
  nand2 gate766(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate767(.a(s_31), .b(gate33inter3), .O(gate33inter10));
  nor2  gate768(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate769(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate770(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1429(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1430(.a(gate35inter0), .b(s_126), .O(gate35inter1));
  and2  gate1431(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1432(.a(s_126), .O(gate35inter3));
  inv1  gate1433(.a(s_127), .O(gate35inter4));
  nand2 gate1434(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1435(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1436(.a(G18), .O(gate35inter7));
  inv1  gate1437(.a(G22), .O(gate35inter8));
  nand2 gate1438(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1439(.a(s_127), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1440(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1441(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1442(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1681(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1682(.a(gate38inter0), .b(s_162), .O(gate38inter1));
  and2  gate1683(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1684(.a(s_162), .O(gate38inter3));
  inv1  gate1685(.a(s_163), .O(gate38inter4));
  nand2 gate1686(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1687(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1688(.a(G27), .O(gate38inter7));
  inv1  gate1689(.a(G31), .O(gate38inter8));
  nand2 gate1690(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1691(.a(s_163), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1692(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1693(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1694(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2045(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2046(.a(gate44inter0), .b(s_214), .O(gate44inter1));
  and2  gate2047(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2048(.a(s_214), .O(gate44inter3));
  inv1  gate2049(.a(s_215), .O(gate44inter4));
  nand2 gate2050(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2051(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2052(.a(G4), .O(gate44inter7));
  inv1  gate2053(.a(G269), .O(gate44inter8));
  nand2 gate2054(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2055(.a(s_215), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2056(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2057(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2058(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1849(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1850(.a(gate46inter0), .b(s_186), .O(gate46inter1));
  and2  gate1851(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1852(.a(s_186), .O(gate46inter3));
  inv1  gate1853(.a(s_187), .O(gate46inter4));
  nand2 gate1854(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1855(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1856(.a(G6), .O(gate46inter7));
  inv1  gate1857(.a(G272), .O(gate46inter8));
  nand2 gate1858(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1859(.a(s_187), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1860(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1861(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1862(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2017(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2018(.a(gate48inter0), .b(s_210), .O(gate48inter1));
  and2  gate2019(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2020(.a(s_210), .O(gate48inter3));
  inv1  gate2021(.a(s_211), .O(gate48inter4));
  nand2 gate2022(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2023(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2024(.a(G8), .O(gate48inter7));
  inv1  gate2025(.a(G275), .O(gate48inter8));
  nand2 gate2026(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2027(.a(s_211), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2028(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2029(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2030(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate2493(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2494(.a(gate49inter0), .b(s_278), .O(gate49inter1));
  and2  gate2495(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2496(.a(s_278), .O(gate49inter3));
  inv1  gate2497(.a(s_279), .O(gate49inter4));
  nand2 gate2498(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2499(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2500(.a(G9), .O(gate49inter7));
  inv1  gate2501(.a(G278), .O(gate49inter8));
  nand2 gate2502(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2503(.a(s_279), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2504(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2505(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2506(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1653(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1654(.a(gate51inter0), .b(s_158), .O(gate51inter1));
  and2  gate1655(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1656(.a(s_158), .O(gate51inter3));
  inv1  gate1657(.a(s_159), .O(gate51inter4));
  nand2 gate1658(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1659(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1660(.a(G11), .O(gate51inter7));
  inv1  gate1661(.a(G281), .O(gate51inter8));
  nand2 gate1662(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1663(.a(s_159), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1664(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1665(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1666(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate981(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate982(.a(gate54inter0), .b(s_62), .O(gate54inter1));
  and2  gate983(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate984(.a(s_62), .O(gate54inter3));
  inv1  gate985(.a(s_63), .O(gate54inter4));
  nand2 gate986(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate987(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate988(.a(G14), .O(gate54inter7));
  inv1  gate989(.a(G284), .O(gate54inter8));
  nand2 gate990(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate991(.a(s_63), .b(gate54inter3), .O(gate54inter10));
  nor2  gate992(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate993(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate994(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1359(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1360(.a(gate57inter0), .b(s_116), .O(gate57inter1));
  and2  gate1361(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1362(.a(s_116), .O(gate57inter3));
  inv1  gate1363(.a(s_117), .O(gate57inter4));
  nand2 gate1364(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1365(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1366(.a(G17), .O(gate57inter7));
  inv1  gate1367(.a(G290), .O(gate57inter8));
  nand2 gate1368(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1369(.a(s_117), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1370(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1371(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1372(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1289(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1290(.a(gate62inter0), .b(s_106), .O(gate62inter1));
  and2  gate1291(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1292(.a(s_106), .O(gate62inter3));
  inv1  gate1293(.a(s_107), .O(gate62inter4));
  nand2 gate1294(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1295(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1296(.a(G22), .O(gate62inter7));
  inv1  gate1297(.a(G296), .O(gate62inter8));
  nand2 gate1298(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1299(.a(s_107), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1300(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1301(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1302(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate883(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate884(.a(gate65inter0), .b(s_48), .O(gate65inter1));
  and2  gate885(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate886(.a(s_48), .O(gate65inter3));
  inv1  gate887(.a(s_49), .O(gate65inter4));
  nand2 gate888(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate889(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate890(.a(G25), .O(gate65inter7));
  inv1  gate891(.a(G302), .O(gate65inter8));
  nand2 gate892(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate893(.a(s_49), .b(gate65inter3), .O(gate65inter10));
  nor2  gate894(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate895(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate896(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1751(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1752(.a(gate69inter0), .b(s_172), .O(gate69inter1));
  and2  gate1753(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1754(.a(s_172), .O(gate69inter3));
  inv1  gate1755(.a(s_173), .O(gate69inter4));
  nand2 gate1756(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1757(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1758(.a(G29), .O(gate69inter7));
  inv1  gate1759(.a(G308), .O(gate69inter8));
  nand2 gate1760(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1761(.a(s_173), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1762(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1763(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1764(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate1695(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1696(.a(gate78inter0), .b(s_164), .O(gate78inter1));
  and2  gate1697(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1698(.a(s_164), .O(gate78inter3));
  inv1  gate1699(.a(s_165), .O(gate78inter4));
  nand2 gate1700(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1701(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1702(.a(G6), .O(gate78inter7));
  inv1  gate1703(.a(G320), .O(gate78inter8));
  nand2 gate1704(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1705(.a(s_165), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1706(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1707(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1708(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2031(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2032(.a(gate81inter0), .b(s_212), .O(gate81inter1));
  and2  gate2033(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2034(.a(s_212), .O(gate81inter3));
  inv1  gate2035(.a(s_213), .O(gate81inter4));
  nand2 gate2036(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2037(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2038(.a(G3), .O(gate81inter7));
  inv1  gate2039(.a(G326), .O(gate81inter8));
  nand2 gate2040(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2041(.a(s_213), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2042(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2043(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2044(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate561(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate562(.a(gate86inter0), .b(s_2), .O(gate86inter1));
  and2  gate563(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate564(.a(s_2), .O(gate86inter3));
  inv1  gate565(.a(s_3), .O(gate86inter4));
  nand2 gate566(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate567(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate568(.a(G8), .O(gate86inter7));
  inv1  gate569(.a(G332), .O(gate86inter8));
  nand2 gate570(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate571(.a(s_3), .b(gate86inter3), .O(gate86inter10));
  nor2  gate572(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate573(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate574(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1947(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1948(.a(gate87inter0), .b(s_200), .O(gate87inter1));
  and2  gate1949(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1950(.a(s_200), .O(gate87inter3));
  inv1  gate1951(.a(s_201), .O(gate87inter4));
  nand2 gate1952(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1953(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1954(.a(G12), .O(gate87inter7));
  inv1  gate1955(.a(G335), .O(gate87inter8));
  nand2 gate1956(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1957(.a(s_201), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1958(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1959(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1960(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate603(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate604(.a(gate88inter0), .b(s_8), .O(gate88inter1));
  and2  gate605(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate606(.a(s_8), .O(gate88inter3));
  inv1  gate607(.a(s_9), .O(gate88inter4));
  nand2 gate608(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate609(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate610(.a(G16), .O(gate88inter7));
  inv1  gate611(.a(G335), .O(gate88inter8));
  nand2 gate612(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate613(.a(s_9), .b(gate88inter3), .O(gate88inter10));
  nor2  gate614(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate615(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate616(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1821(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1822(.a(gate90inter0), .b(s_182), .O(gate90inter1));
  and2  gate1823(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1824(.a(s_182), .O(gate90inter3));
  inv1  gate1825(.a(s_183), .O(gate90inter4));
  nand2 gate1826(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1827(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1828(.a(G21), .O(gate90inter7));
  inv1  gate1829(.a(G338), .O(gate90inter8));
  nand2 gate1830(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1831(.a(s_183), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1832(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1833(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1834(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2521(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2522(.a(gate95inter0), .b(s_282), .O(gate95inter1));
  and2  gate2523(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2524(.a(s_282), .O(gate95inter3));
  inv1  gate2525(.a(s_283), .O(gate95inter4));
  nand2 gate2526(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2527(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2528(.a(G26), .O(gate95inter7));
  inv1  gate2529(.a(G347), .O(gate95inter8));
  nand2 gate2530(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2531(.a(s_283), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2532(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2533(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2534(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1233(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1234(.a(gate98inter0), .b(s_98), .O(gate98inter1));
  and2  gate1235(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1236(.a(s_98), .O(gate98inter3));
  inv1  gate1237(.a(s_99), .O(gate98inter4));
  nand2 gate1238(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1239(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1240(.a(G23), .O(gate98inter7));
  inv1  gate1241(.a(G350), .O(gate98inter8));
  nand2 gate1242(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1243(.a(s_99), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1244(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1245(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1246(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2087(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2088(.a(gate99inter0), .b(s_220), .O(gate99inter1));
  and2  gate2089(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2090(.a(s_220), .O(gate99inter3));
  inv1  gate2091(.a(s_221), .O(gate99inter4));
  nand2 gate2092(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2093(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2094(.a(G27), .O(gate99inter7));
  inv1  gate2095(.a(G353), .O(gate99inter8));
  nand2 gate2096(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2097(.a(s_221), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2098(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2099(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2100(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1345(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1346(.a(gate100inter0), .b(s_114), .O(gate100inter1));
  and2  gate1347(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1348(.a(s_114), .O(gate100inter3));
  inv1  gate1349(.a(s_115), .O(gate100inter4));
  nand2 gate1350(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1351(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1352(.a(G31), .O(gate100inter7));
  inv1  gate1353(.a(G353), .O(gate100inter8));
  nand2 gate1354(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1355(.a(s_115), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1356(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1357(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1358(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2003(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2004(.a(gate106inter0), .b(s_208), .O(gate106inter1));
  and2  gate2005(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2006(.a(s_208), .O(gate106inter3));
  inv1  gate2007(.a(s_209), .O(gate106inter4));
  nand2 gate2008(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2009(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2010(.a(G364), .O(gate106inter7));
  inv1  gate2011(.a(G365), .O(gate106inter8));
  nand2 gate2012(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2013(.a(s_209), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2014(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2015(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2016(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1555(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1556(.a(gate108inter0), .b(s_144), .O(gate108inter1));
  and2  gate1557(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1558(.a(s_144), .O(gate108inter3));
  inv1  gate1559(.a(s_145), .O(gate108inter4));
  nand2 gate1560(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1561(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1562(.a(G368), .O(gate108inter7));
  inv1  gate1563(.a(G369), .O(gate108inter8));
  nand2 gate1564(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1565(.a(s_145), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1566(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1567(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1568(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate631(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate632(.a(gate109inter0), .b(s_12), .O(gate109inter1));
  and2  gate633(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate634(.a(s_12), .O(gate109inter3));
  inv1  gate635(.a(s_13), .O(gate109inter4));
  nand2 gate636(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate637(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate638(.a(G370), .O(gate109inter7));
  inv1  gate639(.a(G371), .O(gate109inter8));
  nand2 gate640(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate641(.a(s_13), .b(gate109inter3), .O(gate109inter10));
  nor2  gate642(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate643(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate644(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate995(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate996(.a(gate112inter0), .b(s_64), .O(gate112inter1));
  and2  gate997(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate998(.a(s_64), .O(gate112inter3));
  inv1  gate999(.a(s_65), .O(gate112inter4));
  nand2 gate1000(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1001(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1002(.a(G376), .O(gate112inter7));
  inv1  gate1003(.a(G377), .O(gate112inter8));
  nand2 gate1004(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1005(.a(s_65), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1006(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1007(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1008(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate2507(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2508(.a(gate113inter0), .b(s_280), .O(gate113inter1));
  and2  gate2509(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2510(.a(s_280), .O(gate113inter3));
  inv1  gate2511(.a(s_281), .O(gate113inter4));
  nand2 gate2512(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2513(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2514(.a(G378), .O(gate113inter7));
  inv1  gate2515(.a(G379), .O(gate113inter8));
  nand2 gate2516(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2517(.a(s_281), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2518(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2519(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2520(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1065(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1066(.a(gate116inter0), .b(s_74), .O(gate116inter1));
  and2  gate1067(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1068(.a(s_74), .O(gate116inter3));
  inv1  gate1069(.a(s_75), .O(gate116inter4));
  nand2 gate1070(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1071(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1072(.a(G384), .O(gate116inter7));
  inv1  gate1073(.a(G385), .O(gate116inter8));
  nand2 gate1074(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1075(.a(s_75), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1076(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1077(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1078(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate2353(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2354(.a(gate117inter0), .b(s_258), .O(gate117inter1));
  and2  gate2355(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2356(.a(s_258), .O(gate117inter3));
  inv1  gate2357(.a(s_259), .O(gate117inter4));
  nand2 gate2358(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2359(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2360(.a(G386), .O(gate117inter7));
  inv1  gate2361(.a(G387), .O(gate117inter8));
  nand2 gate2362(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2363(.a(s_259), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2364(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2365(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2366(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1163(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1164(.a(gate120inter0), .b(s_88), .O(gate120inter1));
  and2  gate1165(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1166(.a(s_88), .O(gate120inter3));
  inv1  gate1167(.a(s_89), .O(gate120inter4));
  nand2 gate1168(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1169(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1170(.a(G392), .O(gate120inter7));
  inv1  gate1171(.a(G393), .O(gate120inter8));
  nand2 gate1172(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1173(.a(s_89), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1174(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1175(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1176(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2367(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2368(.a(gate122inter0), .b(s_260), .O(gate122inter1));
  and2  gate2369(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2370(.a(s_260), .O(gate122inter3));
  inv1  gate2371(.a(s_261), .O(gate122inter4));
  nand2 gate2372(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2373(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2374(.a(G396), .O(gate122inter7));
  inv1  gate2375(.a(G397), .O(gate122inter8));
  nand2 gate2376(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2377(.a(s_261), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2378(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2379(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2380(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate925(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate926(.a(gate123inter0), .b(s_54), .O(gate123inter1));
  and2  gate927(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate928(.a(s_54), .O(gate123inter3));
  inv1  gate929(.a(s_55), .O(gate123inter4));
  nand2 gate930(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate931(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate932(.a(G398), .O(gate123inter7));
  inv1  gate933(.a(G399), .O(gate123inter8));
  nand2 gate934(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate935(.a(s_55), .b(gate123inter3), .O(gate123inter10));
  nor2  gate936(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate937(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate938(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2409(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2410(.a(gate129inter0), .b(s_266), .O(gate129inter1));
  and2  gate2411(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2412(.a(s_266), .O(gate129inter3));
  inv1  gate2413(.a(s_267), .O(gate129inter4));
  nand2 gate2414(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2415(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2416(.a(G410), .O(gate129inter7));
  inv1  gate2417(.a(G411), .O(gate129inter8));
  nand2 gate2418(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2419(.a(s_267), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2420(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2421(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2422(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate2297(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2298(.a(gate130inter0), .b(s_250), .O(gate130inter1));
  and2  gate2299(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2300(.a(s_250), .O(gate130inter3));
  inv1  gate2301(.a(s_251), .O(gate130inter4));
  nand2 gate2302(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2303(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2304(.a(G412), .O(gate130inter7));
  inv1  gate2305(.a(G413), .O(gate130inter8));
  nand2 gate2306(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2307(.a(s_251), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2308(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2309(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2310(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1989(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1990(.a(gate132inter0), .b(s_206), .O(gate132inter1));
  and2  gate1991(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1992(.a(s_206), .O(gate132inter3));
  inv1  gate1993(.a(s_207), .O(gate132inter4));
  nand2 gate1994(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1995(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1996(.a(G416), .O(gate132inter7));
  inv1  gate1997(.a(G417), .O(gate132inter8));
  nand2 gate1998(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1999(.a(s_207), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2000(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2001(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2002(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1933(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1934(.a(gate135inter0), .b(s_198), .O(gate135inter1));
  and2  gate1935(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1936(.a(s_198), .O(gate135inter3));
  inv1  gate1937(.a(s_199), .O(gate135inter4));
  nand2 gate1938(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1939(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1940(.a(G422), .O(gate135inter7));
  inv1  gate1941(.a(G423), .O(gate135inter8));
  nand2 gate1942(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1943(.a(s_199), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1944(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1945(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1946(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate729(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate730(.a(gate136inter0), .b(s_26), .O(gate136inter1));
  and2  gate731(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate732(.a(s_26), .O(gate136inter3));
  inv1  gate733(.a(s_27), .O(gate136inter4));
  nand2 gate734(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate735(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate736(.a(G424), .O(gate136inter7));
  inv1  gate737(.a(G425), .O(gate136inter8));
  nand2 gate738(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate739(.a(s_27), .b(gate136inter3), .O(gate136inter10));
  nor2  gate740(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate741(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate742(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1191(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1192(.a(gate145inter0), .b(s_92), .O(gate145inter1));
  and2  gate1193(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1194(.a(s_92), .O(gate145inter3));
  inv1  gate1195(.a(s_93), .O(gate145inter4));
  nand2 gate1196(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1197(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1198(.a(G474), .O(gate145inter7));
  inv1  gate1199(.a(G477), .O(gate145inter8));
  nand2 gate1200(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1201(.a(s_93), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1202(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1203(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1204(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate2157(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2158(.a(gate146inter0), .b(s_230), .O(gate146inter1));
  and2  gate2159(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2160(.a(s_230), .O(gate146inter3));
  inv1  gate2161(.a(s_231), .O(gate146inter4));
  nand2 gate2162(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2163(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2164(.a(G480), .O(gate146inter7));
  inv1  gate2165(.a(G483), .O(gate146inter8));
  nand2 gate2166(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2167(.a(s_231), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2168(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2169(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2170(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1723(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1724(.a(gate149inter0), .b(s_168), .O(gate149inter1));
  and2  gate1725(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1726(.a(s_168), .O(gate149inter3));
  inv1  gate1727(.a(s_169), .O(gate149inter4));
  nand2 gate1728(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1729(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1730(.a(G498), .O(gate149inter7));
  inv1  gate1731(.a(G501), .O(gate149inter8));
  nand2 gate1732(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1733(.a(s_169), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1734(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1735(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1736(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate771(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate772(.a(gate152inter0), .b(s_32), .O(gate152inter1));
  and2  gate773(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate774(.a(s_32), .O(gate152inter3));
  inv1  gate775(.a(s_33), .O(gate152inter4));
  nand2 gate776(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate777(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate778(.a(G516), .O(gate152inter7));
  inv1  gate779(.a(G519), .O(gate152inter8));
  nand2 gate780(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate781(.a(s_33), .b(gate152inter3), .O(gate152inter10));
  nor2  gate782(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate783(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate784(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2395(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2396(.a(gate156inter0), .b(s_264), .O(gate156inter1));
  and2  gate2397(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2398(.a(s_264), .O(gate156inter3));
  inv1  gate2399(.a(s_265), .O(gate156inter4));
  nand2 gate2400(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2401(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2402(.a(G435), .O(gate156inter7));
  inv1  gate2403(.a(G525), .O(gate156inter8));
  nand2 gate2404(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2405(.a(s_265), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2406(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2407(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2408(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2213(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2214(.a(gate165inter0), .b(s_238), .O(gate165inter1));
  and2  gate2215(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2216(.a(s_238), .O(gate165inter3));
  inv1  gate2217(.a(s_239), .O(gate165inter4));
  nand2 gate2218(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2219(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2220(.a(G462), .O(gate165inter7));
  inv1  gate2221(.a(G540), .O(gate165inter8));
  nand2 gate2222(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2223(.a(s_239), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2224(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2225(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2226(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1625(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1626(.a(gate168inter0), .b(s_154), .O(gate168inter1));
  and2  gate1627(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1628(.a(s_154), .O(gate168inter3));
  inv1  gate1629(.a(s_155), .O(gate168inter4));
  nand2 gate1630(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1631(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1632(.a(G471), .O(gate168inter7));
  inv1  gate1633(.a(G543), .O(gate168inter8));
  nand2 gate1634(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1635(.a(s_155), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1636(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1637(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1638(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1093(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1094(.a(gate169inter0), .b(s_78), .O(gate169inter1));
  and2  gate1095(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1096(.a(s_78), .O(gate169inter3));
  inv1  gate1097(.a(s_79), .O(gate169inter4));
  nand2 gate1098(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1099(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1100(.a(G474), .O(gate169inter7));
  inv1  gate1101(.a(G546), .O(gate169inter8));
  nand2 gate1102(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1103(.a(s_79), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1104(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1105(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1106(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1373(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1374(.a(gate174inter0), .b(s_118), .O(gate174inter1));
  and2  gate1375(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1376(.a(s_118), .O(gate174inter3));
  inv1  gate1377(.a(s_119), .O(gate174inter4));
  nand2 gate1378(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1379(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1380(.a(G489), .O(gate174inter7));
  inv1  gate1381(.a(G552), .O(gate174inter8));
  nand2 gate1382(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1383(.a(s_119), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1384(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1385(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1386(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1051(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1052(.a(gate176inter0), .b(s_72), .O(gate176inter1));
  and2  gate1053(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1054(.a(s_72), .O(gate176inter3));
  inv1  gate1055(.a(s_73), .O(gate176inter4));
  nand2 gate1056(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1057(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1058(.a(G495), .O(gate176inter7));
  inv1  gate1059(.a(G555), .O(gate176inter8));
  nand2 gate1060(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1061(.a(s_73), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1062(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1063(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1064(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1401(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1402(.a(gate178inter0), .b(s_122), .O(gate178inter1));
  and2  gate1403(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1404(.a(s_122), .O(gate178inter3));
  inv1  gate1405(.a(s_123), .O(gate178inter4));
  nand2 gate1406(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1407(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1408(.a(G501), .O(gate178inter7));
  inv1  gate1409(.a(G558), .O(gate178inter8));
  nand2 gate1410(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1411(.a(s_123), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1412(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1413(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1414(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate589(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate590(.a(gate184inter0), .b(s_6), .O(gate184inter1));
  and2  gate591(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate592(.a(s_6), .O(gate184inter3));
  inv1  gate593(.a(s_7), .O(gate184inter4));
  nand2 gate594(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate595(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate596(.a(G519), .O(gate184inter7));
  inv1  gate597(.a(G567), .O(gate184inter8));
  nand2 gate598(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate599(.a(s_7), .b(gate184inter3), .O(gate184inter10));
  nor2  gate600(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate601(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate602(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1247(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1248(.a(gate186inter0), .b(s_100), .O(gate186inter1));
  and2  gate1249(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1250(.a(s_100), .O(gate186inter3));
  inv1  gate1251(.a(s_101), .O(gate186inter4));
  nand2 gate1252(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1253(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1254(.a(G572), .O(gate186inter7));
  inv1  gate1255(.a(G573), .O(gate186inter8));
  nand2 gate1256(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1257(.a(s_101), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1258(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1259(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1260(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate911(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate912(.a(gate191inter0), .b(s_52), .O(gate191inter1));
  and2  gate913(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate914(.a(s_52), .O(gate191inter3));
  inv1  gate915(.a(s_53), .O(gate191inter4));
  nand2 gate916(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate917(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate918(.a(G582), .O(gate191inter7));
  inv1  gate919(.a(G583), .O(gate191inter8));
  nand2 gate920(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate921(.a(s_53), .b(gate191inter3), .O(gate191inter10));
  nor2  gate922(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate923(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate924(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1541(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1542(.a(gate194inter0), .b(s_142), .O(gate194inter1));
  and2  gate1543(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1544(.a(s_142), .O(gate194inter3));
  inv1  gate1545(.a(s_143), .O(gate194inter4));
  nand2 gate1546(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1547(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1548(.a(G588), .O(gate194inter7));
  inv1  gate1549(.a(G589), .O(gate194inter8));
  nand2 gate1550(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1551(.a(s_143), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1552(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1553(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1554(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate2115(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2116(.a(gate195inter0), .b(s_224), .O(gate195inter1));
  and2  gate2117(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2118(.a(s_224), .O(gate195inter3));
  inv1  gate2119(.a(s_225), .O(gate195inter4));
  nand2 gate2120(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2121(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2122(.a(G590), .O(gate195inter7));
  inv1  gate2123(.a(G591), .O(gate195inter8));
  nand2 gate2124(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2125(.a(s_225), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2126(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2127(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2128(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1331(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1332(.a(gate196inter0), .b(s_112), .O(gate196inter1));
  and2  gate1333(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1334(.a(s_112), .O(gate196inter3));
  inv1  gate1335(.a(s_113), .O(gate196inter4));
  nand2 gate1336(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1337(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1338(.a(G592), .O(gate196inter7));
  inv1  gate1339(.a(G593), .O(gate196inter8));
  nand2 gate1340(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1341(.a(s_113), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1342(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1343(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1344(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2423(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2424(.a(gate200inter0), .b(s_268), .O(gate200inter1));
  and2  gate2425(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2426(.a(s_268), .O(gate200inter3));
  inv1  gate2427(.a(s_269), .O(gate200inter4));
  nand2 gate2428(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2429(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2430(.a(G600), .O(gate200inter7));
  inv1  gate2431(.a(G601), .O(gate200inter8));
  nand2 gate2432(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2433(.a(s_269), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2434(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2435(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2436(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2059(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2060(.a(gate207inter0), .b(s_216), .O(gate207inter1));
  and2  gate2061(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2062(.a(s_216), .O(gate207inter3));
  inv1  gate2063(.a(s_217), .O(gate207inter4));
  nand2 gate2064(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2065(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2066(.a(G622), .O(gate207inter7));
  inv1  gate2067(.a(G632), .O(gate207inter8));
  nand2 gate2068(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2069(.a(s_217), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2070(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2071(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2072(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2381(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2382(.a(gate209inter0), .b(s_262), .O(gate209inter1));
  and2  gate2383(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2384(.a(s_262), .O(gate209inter3));
  inv1  gate2385(.a(s_263), .O(gate209inter4));
  nand2 gate2386(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2387(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2388(.a(G602), .O(gate209inter7));
  inv1  gate2389(.a(G666), .O(gate209inter8));
  nand2 gate2390(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2391(.a(s_263), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2392(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2393(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2394(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate2549(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2550(.a(gate210inter0), .b(s_286), .O(gate210inter1));
  and2  gate2551(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2552(.a(s_286), .O(gate210inter3));
  inv1  gate2553(.a(s_287), .O(gate210inter4));
  nand2 gate2554(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2555(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2556(.a(G607), .O(gate210inter7));
  inv1  gate2557(.a(G666), .O(gate210inter8));
  nand2 gate2558(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2559(.a(s_287), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2560(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2561(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2562(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate2535(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2536(.a(gate211inter0), .b(s_284), .O(gate211inter1));
  and2  gate2537(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2538(.a(s_284), .O(gate211inter3));
  inv1  gate2539(.a(s_285), .O(gate211inter4));
  nand2 gate2540(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2541(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2542(.a(G612), .O(gate211inter7));
  inv1  gate2543(.a(G669), .O(gate211inter8));
  nand2 gate2544(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2545(.a(s_285), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2546(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2547(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2548(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate547(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate548(.a(gate213inter0), .b(s_0), .O(gate213inter1));
  and2  gate549(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate550(.a(s_0), .O(gate213inter3));
  inv1  gate551(.a(s_1), .O(gate213inter4));
  nand2 gate552(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate553(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate554(.a(G602), .O(gate213inter7));
  inv1  gate555(.a(G672), .O(gate213inter8));
  nand2 gate556(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate557(.a(s_1), .b(gate213inter3), .O(gate213inter10));
  nor2  gate558(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate559(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate560(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1877(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1878(.a(gate215inter0), .b(s_190), .O(gate215inter1));
  and2  gate1879(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1880(.a(s_190), .O(gate215inter3));
  inv1  gate1881(.a(s_191), .O(gate215inter4));
  nand2 gate1882(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1883(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1884(.a(G607), .O(gate215inter7));
  inv1  gate1885(.a(G675), .O(gate215inter8));
  nand2 gate1886(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1887(.a(s_191), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1888(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1889(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1890(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1779(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1780(.a(gate216inter0), .b(s_176), .O(gate216inter1));
  and2  gate1781(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1782(.a(s_176), .O(gate216inter3));
  inv1  gate1783(.a(s_177), .O(gate216inter4));
  nand2 gate1784(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1785(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1786(.a(G617), .O(gate216inter7));
  inv1  gate1787(.a(G675), .O(gate216inter8));
  nand2 gate1788(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1789(.a(s_177), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1790(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1791(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1792(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate785(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate786(.a(gate219inter0), .b(s_34), .O(gate219inter1));
  and2  gate787(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate788(.a(s_34), .O(gate219inter3));
  inv1  gate789(.a(s_35), .O(gate219inter4));
  nand2 gate790(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate791(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate792(.a(G632), .O(gate219inter7));
  inv1  gate793(.a(G681), .O(gate219inter8));
  nand2 gate794(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate795(.a(s_35), .b(gate219inter3), .O(gate219inter10));
  nor2  gate796(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate797(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate798(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2241(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2242(.a(gate223inter0), .b(s_242), .O(gate223inter1));
  and2  gate2243(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2244(.a(s_242), .O(gate223inter3));
  inv1  gate2245(.a(s_243), .O(gate223inter4));
  nand2 gate2246(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2247(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2248(.a(G627), .O(gate223inter7));
  inv1  gate2249(.a(G687), .O(gate223inter8));
  nand2 gate2250(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2251(.a(s_243), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2252(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2253(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2254(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2143(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2144(.a(gate227inter0), .b(s_228), .O(gate227inter1));
  and2  gate2145(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2146(.a(s_228), .O(gate227inter3));
  inv1  gate2147(.a(s_229), .O(gate227inter4));
  nand2 gate2148(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2149(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2150(.a(G694), .O(gate227inter7));
  inv1  gate2151(.a(G695), .O(gate227inter8));
  nand2 gate2152(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2153(.a(s_229), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2154(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2155(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2156(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1387(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1388(.a(gate228inter0), .b(s_120), .O(gate228inter1));
  and2  gate1389(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1390(.a(s_120), .O(gate228inter3));
  inv1  gate1391(.a(s_121), .O(gate228inter4));
  nand2 gate1392(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1393(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1394(.a(G696), .O(gate228inter7));
  inv1  gate1395(.a(G697), .O(gate228inter8));
  nand2 gate1396(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1397(.a(s_121), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1398(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1399(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1400(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate855(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate856(.a(gate229inter0), .b(s_44), .O(gate229inter1));
  and2  gate857(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate858(.a(s_44), .O(gate229inter3));
  inv1  gate859(.a(s_45), .O(gate229inter4));
  nand2 gate860(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate861(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate862(.a(G698), .O(gate229inter7));
  inv1  gate863(.a(G699), .O(gate229inter8));
  nand2 gate864(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate865(.a(s_45), .b(gate229inter3), .O(gate229inter10));
  nor2  gate866(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate867(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate868(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1037(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1038(.a(gate235inter0), .b(s_70), .O(gate235inter1));
  and2  gate1039(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1040(.a(s_70), .O(gate235inter3));
  inv1  gate1041(.a(s_71), .O(gate235inter4));
  nand2 gate1042(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1043(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1044(.a(G248), .O(gate235inter7));
  inv1  gate1045(.a(G724), .O(gate235inter8));
  nand2 gate1046(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1047(.a(s_71), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1048(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1049(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1050(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1527(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1528(.a(gate242inter0), .b(s_140), .O(gate242inter1));
  and2  gate1529(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1530(.a(s_140), .O(gate242inter3));
  inv1  gate1531(.a(s_141), .O(gate242inter4));
  nand2 gate1532(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1533(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1534(.a(G718), .O(gate242inter7));
  inv1  gate1535(.a(G730), .O(gate242inter8));
  nand2 gate1536(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1537(.a(s_141), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1538(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1539(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1540(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1457(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1458(.a(gate244inter0), .b(s_130), .O(gate244inter1));
  and2  gate1459(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1460(.a(s_130), .O(gate244inter3));
  inv1  gate1461(.a(s_131), .O(gate244inter4));
  nand2 gate1462(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1463(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1464(.a(G721), .O(gate244inter7));
  inv1  gate1465(.a(G733), .O(gate244inter8));
  nand2 gate1466(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1467(.a(s_131), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1468(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1469(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1470(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1443(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1444(.a(gate246inter0), .b(s_128), .O(gate246inter1));
  and2  gate1445(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1446(.a(s_128), .O(gate246inter3));
  inv1  gate1447(.a(s_129), .O(gate246inter4));
  nand2 gate1448(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1449(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1450(.a(G724), .O(gate246inter7));
  inv1  gate1451(.a(G736), .O(gate246inter8));
  nand2 gate1452(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1453(.a(s_129), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1454(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1455(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1456(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1807(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1808(.a(gate249inter0), .b(s_180), .O(gate249inter1));
  and2  gate1809(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1810(.a(s_180), .O(gate249inter3));
  inv1  gate1811(.a(s_181), .O(gate249inter4));
  nand2 gate1812(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1813(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1814(.a(G254), .O(gate249inter7));
  inv1  gate1815(.a(G742), .O(gate249inter8));
  nand2 gate1816(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1817(.a(s_181), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1818(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1819(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1820(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1583(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1584(.a(gate250inter0), .b(s_148), .O(gate250inter1));
  and2  gate1585(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1586(.a(s_148), .O(gate250inter3));
  inv1  gate1587(.a(s_149), .O(gate250inter4));
  nand2 gate1588(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1589(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1590(.a(G706), .O(gate250inter7));
  inv1  gate1591(.a(G742), .O(gate250inter8));
  nand2 gate1592(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1593(.a(s_149), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1594(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1595(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1596(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1107(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1108(.a(gate251inter0), .b(s_80), .O(gate251inter1));
  and2  gate1109(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1110(.a(s_80), .O(gate251inter3));
  inv1  gate1111(.a(s_81), .O(gate251inter4));
  nand2 gate1112(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1113(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1114(.a(G257), .O(gate251inter7));
  inv1  gate1115(.a(G745), .O(gate251inter8));
  nand2 gate1116(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1117(.a(s_81), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1118(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1119(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1120(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate701(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate702(.a(gate252inter0), .b(s_22), .O(gate252inter1));
  and2  gate703(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate704(.a(s_22), .O(gate252inter3));
  inv1  gate705(.a(s_23), .O(gate252inter4));
  nand2 gate706(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate707(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate708(.a(G709), .O(gate252inter7));
  inv1  gate709(.a(G745), .O(gate252inter8));
  nand2 gate710(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate711(.a(s_23), .b(gate252inter3), .O(gate252inter10));
  nor2  gate712(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate713(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate714(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate939(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate940(.a(gate253inter0), .b(s_56), .O(gate253inter1));
  and2  gate941(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate942(.a(s_56), .O(gate253inter3));
  inv1  gate943(.a(s_57), .O(gate253inter4));
  nand2 gate944(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate945(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate946(.a(G260), .O(gate253inter7));
  inv1  gate947(.a(G748), .O(gate253inter8));
  nand2 gate948(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate949(.a(s_57), .b(gate253inter3), .O(gate253inter10));
  nor2  gate950(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate951(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate952(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1863(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1864(.a(gate255inter0), .b(s_188), .O(gate255inter1));
  and2  gate1865(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1866(.a(s_188), .O(gate255inter3));
  inv1  gate1867(.a(s_189), .O(gate255inter4));
  nand2 gate1868(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1869(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1870(.a(G263), .O(gate255inter7));
  inv1  gate1871(.a(G751), .O(gate255inter8));
  nand2 gate1872(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1873(.a(s_189), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1874(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1875(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1876(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate827(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate828(.a(gate258inter0), .b(s_40), .O(gate258inter1));
  and2  gate829(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate830(.a(s_40), .O(gate258inter3));
  inv1  gate831(.a(s_41), .O(gate258inter4));
  nand2 gate832(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate833(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate834(.a(G756), .O(gate258inter7));
  inv1  gate835(.a(G757), .O(gate258inter8));
  nand2 gate836(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate837(.a(s_41), .b(gate258inter3), .O(gate258inter10));
  nor2  gate838(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate839(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate840(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1975(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1976(.a(gate261inter0), .b(s_204), .O(gate261inter1));
  and2  gate1977(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1978(.a(s_204), .O(gate261inter3));
  inv1  gate1979(.a(s_205), .O(gate261inter4));
  nand2 gate1980(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1981(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1982(.a(G762), .O(gate261inter7));
  inv1  gate1983(.a(G763), .O(gate261inter8));
  nand2 gate1984(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1985(.a(s_205), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1986(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1987(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1988(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2325(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2326(.a(gate264inter0), .b(s_254), .O(gate264inter1));
  and2  gate2327(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2328(.a(s_254), .O(gate264inter3));
  inv1  gate2329(.a(s_255), .O(gate264inter4));
  nand2 gate2330(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2331(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2332(.a(G768), .O(gate264inter7));
  inv1  gate2333(.a(G769), .O(gate264inter8));
  nand2 gate2334(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2335(.a(s_255), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2336(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2337(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2338(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1569(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1570(.a(gate268inter0), .b(s_146), .O(gate268inter1));
  and2  gate1571(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1572(.a(s_146), .O(gate268inter3));
  inv1  gate1573(.a(s_147), .O(gate268inter4));
  nand2 gate1574(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1575(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1576(.a(G651), .O(gate268inter7));
  inv1  gate1577(.a(G779), .O(gate268inter8));
  nand2 gate1578(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1579(.a(s_147), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1580(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1581(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1582(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate2199(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate2200(.a(gate273inter0), .b(s_236), .O(gate273inter1));
  and2  gate2201(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate2202(.a(s_236), .O(gate273inter3));
  inv1  gate2203(.a(s_237), .O(gate273inter4));
  nand2 gate2204(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate2205(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate2206(.a(G642), .O(gate273inter7));
  inv1  gate2207(.a(G794), .O(gate273inter8));
  nand2 gate2208(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate2209(.a(s_237), .b(gate273inter3), .O(gate273inter10));
  nor2  gate2210(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate2211(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate2212(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate2437(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2438(.a(gate276inter0), .b(s_270), .O(gate276inter1));
  and2  gate2439(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2440(.a(s_270), .O(gate276inter3));
  inv1  gate2441(.a(s_271), .O(gate276inter4));
  nand2 gate2442(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2443(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2444(.a(G773), .O(gate276inter7));
  inv1  gate2445(.a(G797), .O(gate276inter8));
  nand2 gate2446(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2447(.a(s_271), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2448(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2449(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2450(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate2563(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2564(.a(gate280inter0), .b(s_288), .O(gate280inter1));
  and2  gate2565(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2566(.a(s_288), .O(gate280inter3));
  inv1  gate2567(.a(s_289), .O(gate280inter4));
  nand2 gate2568(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2569(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2570(.a(G779), .O(gate280inter7));
  inv1  gate2571(.a(G803), .O(gate280inter8));
  nand2 gate2572(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2573(.a(s_289), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2574(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2575(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2576(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1639(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1640(.a(gate289inter0), .b(s_156), .O(gate289inter1));
  and2  gate1641(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1642(.a(s_156), .O(gate289inter3));
  inv1  gate1643(.a(s_157), .O(gate289inter4));
  nand2 gate1644(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1645(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1646(.a(G818), .O(gate289inter7));
  inv1  gate1647(.a(G819), .O(gate289inter8));
  nand2 gate1648(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1649(.a(s_157), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1650(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1651(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1652(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2101(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2102(.a(gate291inter0), .b(s_222), .O(gate291inter1));
  and2  gate2103(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2104(.a(s_222), .O(gate291inter3));
  inv1  gate2105(.a(s_223), .O(gate291inter4));
  nand2 gate2106(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2107(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2108(.a(G822), .O(gate291inter7));
  inv1  gate2109(.a(G823), .O(gate291inter8));
  nand2 gate2110(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2111(.a(s_223), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2112(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2113(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2114(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate673(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate674(.a(gate292inter0), .b(s_18), .O(gate292inter1));
  and2  gate675(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate676(.a(s_18), .O(gate292inter3));
  inv1  gate677(.a(s_19), .O(gate292inter4));
  nand2 gate678(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate679(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate680(.a(G824), .O(gate292inter7));
  inv1  gate681(.a(G825), .O(gate292inter8));
  nand2 gate682(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate683(.a(s_19), .b(gate292inter3), .O(gate292inter10));
  nor2  gate684(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate685(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate686(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1597(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1598(.a(gate293inter0), .b(s_150), .O(gate293inter1));
  and2  gate1599(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1600(.a(s_150), .O(gate293inter3));
  inv1  gate1601(.a(s_151), .O(gate293inter4));
  nand2 gate1602(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1603(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1604(.a(G828), .O(gate293inter7));
  inv1  gate1605(.a(G829), .O(gate293inter8));
  nand2 gate1606(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1607(.a(s_151), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1608(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1609(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1610(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1009(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1010(.a(gate390inter0), .b(s_66), .O(gate390inter1));
  and2  gate1011(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1012(.a(s_66), .O(gate390inter3));
  inv1  gate1013(.a(s_67), .O(gate390inter4));
  nand2 gate1014(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1015(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1016(.a(G4), .O(gate390inter7));
  inv1  gate1017(.a(G1045), .O(gate390inter8));
  nand2 gate1018(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1019(.a(s_67), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1020(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1021(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1022(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1121(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1122(.a(gate393inter0), .b(s_82), .O(gate393inter1));
  and2  gate1123(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1124(.a(s_82), .O(gate393inter3));
  inv1  gate1125(.a(s_83), .O(gate393inter4));
  nand2 gate1126(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1127(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1128(.a(G7), .O(gate393inter7));
  inv1  gate1129(.a(G1054), .O(gate393inter8));
  nand2 gate1130(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1131(.a(s_83), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1132(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1133(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1134(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate2171(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2172(.a(gate394inter0), .b(s_232), .O(gate394inter1));
  and2  gate2173(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2174(.a(s_232), .O(gate394inter3));
  inv1  gate2175(.a(s_233), .O(gate394inter4));
  nand2 gate2176(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2177(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2178(.a(G8), .O(gate394inter7));
  inv1  gate2179(.a(G1057), .O(gate394inter8));
  nand2 gate2180(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2181(.a(s_233), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2182(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2183(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2184(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate813(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate814(.a(gate395inter0), .b(s_38), .O(gate395inter1));
  and2  gate815(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate816(.a(s_38), .O(gate395inter3));
  inv1  gate817(.a(s_39), .O(gate395inter4));
  nand2 gate818(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate819(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate820(.a(G9), .O(gate395inter7));
  inv1  gate821(.a(G1060), .O(gate395inter8));
  nand2 gate822(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate823(.a(s_39), .b(gate395inter3), .O(gate395inter10));
  nor2  gate824(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate825(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate826(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2311(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2312(.a(gate396inter0), .b(s_252), .O(gate396inter1));
  and2  gate2313(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2314(.a(s_252), .O(gate396inter3));
  inv1  gate2315(.a(s_253), .O(gate396inter4));
  nand2 gate2316(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2317(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2318(.a(G10), .O(gate396inter7));
  inv1  gate2319(.a(G1063), .O(gate396inter8));
  nand2 gate2320(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2321(.a(s_253), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2322(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2323(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2324(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1205(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1206(.a(gate399inter0), .b(s_94), .O(gate399inter1));
  and2  gate1207(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1208(.a(s_94), .O(gate399inter3));
  inv1  gate1209(.a(s_95), .O(gate399inter4));
  nand2 gate1210(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1211(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1212(.a(G13), .O(gate399inter7));
  inv1  gate1213(.a(G1072), .O(gate399inter8));
  nand2 gate1214(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1215(.a(s_95), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1216(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1217(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1218(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate715(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate716(.a(gate403inter0), .b(s_24), .O(gate403inter1));
  and2  gate717(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate718(.a(s_24), .O(gate403inter3));
  inv1  gate719(.a(s_25), .O(gate403inter4));
  nand2 gate720(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate721(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate722(.a(G17), .O(gate403inter7));
  inv1  gate723(.a(G1084), .O(gate403inter8));
  nand2 gate724(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate725(.a(s_25), .b(gate403inter3), .O(gate403inter10));
  nor2  gate726(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate727(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate728(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1079(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1080(.a(gate405inter0), .b(s_76), .O(gate405inter1));
  and2  gate1081(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1082(.a(s_76), .O(gate405inter3));
  inv1  gate1083(.a(s_77), .O(gate405inter4));
  nand2 gate1084(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1085(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1086(.a(G19), .O(gate405inter7));
  inv1  gate1087(.a(G1090), .O(gate405inter8));
  nand2 gate1088(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1089(.a(s_77), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1090(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1091(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1092(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate659(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate660(.a(gate406inter0), .b(s_16), .O(gate406inter1));
  and2  gate661(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate662(.a(s_16), .O(gate406inter3));
  inv1  gate663(.a(s_17), .O(gate406inter4));
  nand2 gate664(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate665(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate666(.a(G20), .O(gate406inter7));
  inv1  gate667(.a(G1093), .O(gate406inter8));
  nand2 gate668(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate669(.a(s_17), .b(gate406inter3), .O(gate406inter10));
  nor2  gate670(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate671(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate672(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1471(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1472(.a(gate407inter0), .b(s_132), .O(gate407inter1));
  and2  gate1473(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1474(.a(s_132), .O(gate407inter3));
  inv1  gate1475(.a(s_133), .O(gate407inter4));
  nand2 gate1476(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1477(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1478(.a(G21), .O(gate407inter7));
  inv1  gate1479(.a(G1096), .O(gate407inter8));
  nand2 gate1480(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1481(.a(s_133), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1482(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1483(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1484(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1737(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1738(.a(gate411inter0), .b(s_170), .O(gate411inter1));
  and2  gate1739(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1740(.a(s_170), .O(gate411inter3));
  inv1  gate1741(.a(s_171), .O(gate411inter4));
  nand2 gate1742(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1743(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1744(.a(G25), .O(gate411inter7));
  inv1  gate1745(.a(G1108), .O(gate411inter8));
  nand2 gate1746(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1747(.a(s_171), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1748(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1749(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1750(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2269(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2270(.a(gate412inter0), .b(s_246), .O(gate412inter1));
  and2  gate2271(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2272(.a(s_246), .O(gate412inter3));
  inv1  gate2273(.a(s_247), .O(gate412inter4));
  nand2 gate2274(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2275(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2276(.a(G26), .O(gate412inter7));
  inv1  gate2277(.a(G1111), .O(gate412inter8));
  nand2 gate2278(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2279(.a(s_247), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2280(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2281(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2282(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate645(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate646(.a(gate416inter0), .b(s_14), .O(gate416inter1));
  and2  gate647(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate648(.a(s_14), .O(gate416inter3));
  inv1  gate649(.a(s_15), .O(gate416inter4));
  nand2 gate650(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate651(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate652(.a(G30), .O(gate416inter7));
  inv1  gate653(.a(G1123), .O(gate416inter8));
  nand2 gate654(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate655(.a(s_15), .b(gate416inter3), .O(gate416inter10));
  nor2  gate656(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate657(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate658(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1261(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1262(.a(gate421inter0), .b(s_102), .O(gate421inter1));
  and2  gate1263(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1264(.a(s_102), .O(gate421inter3));
  inv1  gate1265(.a(s_103), .O(gate421inter4));
  nand2 gate1266(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1267(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1268(.a(G2), .O(gate421inter7));
  inv1  gate1269(.a(G1135), .O(gate421inter8));
  nand2 gate1270(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1271(.a(s_103), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1272(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1273(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1274(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1485(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1486(.a(gate423inter0), .b(s_134), .O(gate423inter1));
  and2  gate1487(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1488(.a(s_134), .O(gate423inter3));
  inv1  gate1489(.a(s_135), .O(gate423inter4));
  nand2 gate1490(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1491(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1492(.a(G3), .O(gate423inter7));
  inv1  gate1493(.a(G1138), .O(gate423inter8));
  nand2 gate1494(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1495(.a(s_135), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1496(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1497(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1498(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1835(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1836(.a(gate429inter0), .b(s_184), .O(gate429inter1));
  and2  gate1837(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1838(.a(s_184), .O(gate429inter3));
  inv1  gate1839(.a(s_185), .O(gate429inter4));
  nand2 gate1840(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1841(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1842(.a(G6), .O(gate429inter7));
  inv1  gate1843(.a(G1147), .O(gate429inter8));
  nand2 gate1844(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1845(.a(s_185), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1846(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1847(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1848(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate2129(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2130(.a(gate430inter0), .b(s_226), .O(gate430inter1));
  and2  gate2131(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2132(.a(s_226), .O(gate430inter3));
  inv1  gate2133(.a(s_227), .O(gate430inter4));
  nand2 gate2134(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2135(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2136(.a(G1051), .O(gate430inter7));
  inv1  gate2137(.a(G1147), .O(gate430inter8));
  nand2 gate2138(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2139(.a(s_227), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2140(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2141(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2142(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1961(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1962(.a(gate431inter0), .b(s_202), .O(gate431inter1));
  and2  gate1963(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1964(.a(s_202), .O(gate431inter3));
  inv1  gate1965(.a(s_203), .O(gate431inter4));
  nand2 gate1966(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1967(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1968(.a(G7), .O(gate431inter7));
  inv1  gate1969(.a(G1150), .O(gate431inter8));
  nand2 gate1970(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1971(.a(s_203), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1972(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1973(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1974(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1275(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1276(.a(gate433inter0), .b(s_104), .O(gate433inter1));
  and2  gate1277(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1278(.a(s_104), .O(gate433inter3));
  inv1  gate1279(.a(s_105), .O(gate433inter4));
  nand2 gate1280(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1281(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1282(.a(G8), .O(gate433inter7));
  inv1  gate1283(.a(G1153), .O(gate433inter8));
  nand2 gate1284(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1285(.a(s_105), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1286(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1287(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1288(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate2451(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2452(.a(gate436inter0), .b(s_272), .O(gate436inter1));
  and2  gate2453(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2454(.a(s_272), .O(gate436inter3));
  inv1  gate2455(.a(s_273), .O(gate436inter4));
  nand2 gate2456(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2457(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2458(.a(G1060), .O(gate436inter7));
  inv1  gate2459(.a(G1156), .O(gate436inter8));
  nand2 gate2460(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2461(.a(s_273), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2462(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2463(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2464(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate953(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate954(.a(gate440inter0), .b(s_58), .O(gate440inter1));
  and2  gate955(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate956(.a(s_58), .O(gate440inter3));
  inv1  gate957(.a(s_59), .O(gate440inter4));
  nand2 gate958(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate959(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate960(.a(G1066), .O(gate440inter7));
  inv1  gate961(.a(G1162), .O(gate440inter8));
  nand2 gate962(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate963(.a(s_59), .b(gate440inter3), .O(gate440inter10));
  nor2  gate964(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate965(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate966(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1919(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1920(.a(gate441inter0), .b(s_196), .O(gate441inter1));
  and2  gate1921(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1922(.a(s_196), .O(gate441inter3));
  inv1  gate1923(.a(s_197), .O(gate441inter4));
  nand2 gate1924(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1925(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1926(.a(G12), .O(gate441inter7));
  inv1  gate1927(.a(G1165), .O(gate441inter8));
  nand2 gate1928(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1929(.a(s_197), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1930(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1931(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1932(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1709(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1710(.a(gate445inter0), .b(s_166), .O(gate445inter1));
  and2  gate1711(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1712(.a(s_166), .O(gate445inter3));
  inv1  gate1713(.a(s_167), .O(gate445inter4));
  nand2 gate1714(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1715(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1716(.a(G14), .O(gate445inter7));
  inv1  gate1717(.a(G1171), .O(gate445inter8));
  nand2 gate1718(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1719(.a(s_167), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1720(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1721(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1722(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1499(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1500(.a(gate450inter0), .b(s_136), .O(gate450inter1));
  and2  gate1501(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1502(.a(s_136), .O(gate450inter3));
  inv1  gate1503(.a(s_137), .O(gate450inter4));
  nand2 gate1504(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1505(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1506(.a(G1081), .O(gate450inter7));
  inv1  gate1507(.a(G1177), .O(gate450inter8));
  nand2 gate1508(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1509(.a(s_137), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1510(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1511(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1512(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2283(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2284(.a(gate451inter0), .b(s_248), .O(gate451inter1));
  and2  gate2285(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2286(.a(s_248), .O(gate451inter3));
  inv1  gate2287(.a(s_249), .O(gate451inter4));
  nand2 gate2288(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2289(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2290(.a(G17), .O(gate451inter7));
  inv1  gate2291(.a(G1180), .O(gate451inter8));
  nand2 gate2292(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2293(.a(s_249), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2294(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2295(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2296(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1891(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1892(.a(gate452inter0), .b(s_192), .O(gate452inter1));
  and2  gate1893(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1894(.a(s_192), .O(gate452inter3));
  inv1  gate1895(.a(s_193), .O(gate452inter4));
  nand2 gate1896(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1897(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1898(.a(G1084), .O(gate452inter7));
  inv1  gate1899(.a(G1180), .O(gate452inter8));
  nand2 gate1900(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1901(.a(s_193), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1902(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1903(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1904(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate841(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate842(.a(gate453inter0), .b(s_42), .O(gate453inter1));
  and2  gate843(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate844(.a(s_42), .O(gate453inter3));
  inv1  gate845(.a(s_43), .O(gate453inter4));
  nand2 gate846(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate847(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate848(.a(G18), .O(gate453inter7));
  inv1  gate849(.a(G1183), .O(gate453inter8));
  nand2 gate850(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate851(.a(s_43), .b(gate453inter3), .O(gate453inter10));
  nor2  gate852(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate853(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate854(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate869(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate870(.a(gate455inter0), .b(s_46), .O(gate455inter1));
  and2  gate871(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate872(.a(s_46), .O(gate455inter3));
  inv1  gate873(.a(s_47), .O(gate455inter4));
  nand2 gate874(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate875(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate876(.a(G19), .O(gate455inter7));
  inv1  gate877(.a(G1186), .O(gate455inter8));
  nand2 gate878(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate879(.a(s_47), .b(gate455inter3), .O(gate455inter10));
  nor2  gate880(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate881(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate882(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate2339(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2340(.a(gate456inter0), .b(s_256), .O(gate456inter1));
  and2  gate2341(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2342(.a(s_256), .O(gate456inter3));
  inv1  gate2343(.a(s_257), .O(gate456inter4));
  nand2 gate2344(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2345(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2346(.a(G1090), .O(gate456inter7));
  inv1  gate2347(.a(G1186), .O(gate456inter8));
  nand2 gate2348(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2349(.a(s_257), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2350(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2351(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2352(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1765(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1766(.a(gate458inter0), .b(s_174), .O(gate458inter1));
  and2  gate1767(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1768(.a(s_174), .O(gate458inter3));
  inv1  gate1769(.a(s_175), .O(gate458inter4));
  nand2 gate1770(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1771(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1772(.a(G1093), .O(gate458inter7));
  inv1  gate1773(.a(G1189), .O(gate458inter8));
  nand2 gate1774(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1775(.a(s_175), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1776(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1777(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1778(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate2465(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2466(.a(gate465inter0), .b(s_274), .O(gate465inter1));
  and2  gate2467(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2468(.a(s_274), .O(gate465inter3));
  inv1  gate2469(.a(s_275), .O(gate465inter4));
  nand2 gate2470(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2471(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2472(.a(G24), .O(gate465inter7));
  inv1  gate2473(.a(G1201), .O(gate465inter8));
  nand2 gate2474(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2475(.a(s_275), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2476(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2477(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2478(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2185(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2186(.a(gate470inter0), .b(s_234), .O(gate470inter1));
  and2  gate2187(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2188(.a(s_234), .O(gate470inter3));
  inv1  gate2189(.a(s_235), .O(gate470inter4));
  nand2 gate2190(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2191(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2192(.a(G1111), .O(gate470inter7));
  inv1  gate2193(.a(G1207), .O(gate470inter8));
  nand2 gate2194(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2195(.a(s_235), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2196(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2197(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2198(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1611(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1612(.a(gate472inter0), .b(s_152), .O(gate472inter1));
  and2  gate1613(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1614(.a(s_152), .O(gate472inter3));
  inv1  gate1615(.a(s_153), .O(gate472inter4));
  nand2 gate1616(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1617(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1618(.a(G1114), .O(gate472inter7));
  inv1  gate1619(.a(G1210), .O(gate472inter8));
  nand2 gate1620(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1621(.a(s_153), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1622(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1623(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1624(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2577(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2578(.a(gate475inter0), .b(s_290), .O(gate475inter1));
  and2  gate2579(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2580(.a(s_290), .O(gate475inter3));
  inv1  gate2581(.a(s_291), .O(gate475inter4));
  nand2 gate2582(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2583(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2584(.a(G29), .O(gate475inter7));
  inv1  gate2585(.a(G1216), .O(gate475inter8));
  nand2 gate2586(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2587(.a(s_291), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2588(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2589(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2590(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1023(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1024(.a(gate476inter0), .b(s_68), .O(gate476inter1));
  and2  gate1025(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1026(.a(s_68), .O(gate476inter3));
  inv1  gate1027(.a(s_69), .O(gate476inter4));
  nand2 gate1028(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1029(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1030(.a(G1120), .O(gate476inter7));
  inv1  gate1031(.a(G1216), .O(gate476inter8));
  nand2 gate1032(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1033(.a(s_69), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1034(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1035(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1036(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1415(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1416(.a(gate477inter0), .b(s_124), .O(gate477inter1));
  and2  gate1417(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1418(.a(s_124), .O(gate477inter3));
  inv1  gate1419(.a(s_125), .O(gate477inter4));
  nand2 gate1420(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1421(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1422(.a(G30), .O(gate477inter7));
  inv1  gate1423(.a(G1219), .O(gate477inter8));
  nand2 gate1424(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1425(.a(s_125), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1426(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1427(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1428(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate799(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate800(.a(gate478inter0), .b(s_36), .O(gate478inter1));
  and2  gate801(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate802(.a(s_36), .O(gate478inter3));
  inv1  gate803(.a(s_37), .O(gate478inter4));
  nand2 gate804(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate805(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate806(.a(G1123), .O(gate478inter7));
  inv1  gate807(.a(G1219), .O(gate478inter8));
  nand2 gate808(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate809(.a(s_37), .b(gate478inter3), .O(gate478inter10));
  nor2  gate810(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate811(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate812(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1135(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1136(.a(gate480inter0), .b(s_84), .O(gate480inter1));
  and2  gate1137(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1138(.a(s_84), .O(gate480inter3));
  inv1  gate1139(.a(s_85), .O(gate480inter4));
  nand2 gate1140(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1141(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1142(.a(G1126), .O(gate480inter7));
  inv1  gate1143(.a(G1222), .O(gate480inter8));
  nand2 gate1144(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1145(.a(s_85), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1146(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1147(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1148(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1905(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1906(.a(gate483inter0), .b(s_194), .O(gate483inter1));
  and2  gate1907(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1908(.a(s_194), .O(gate483inter3));
  inv1  gate1909(.a(s_195), .O(gate483inter4));
  nand2 gate1910(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1911(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1912(.a(G1228), .O(gate483inter7));
  inv1  gate1913(.a(G1229), .O(gate483inter8));
  nand2 gate1914(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1915(.a(s_195), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1916(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1917(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1918(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1667(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1668(.a(gate486inter0), .b(s_160), .O(gate486inter1));
  and2  gate1669(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1670(.a(s_160), .O(gate486inter3));
  inv1  gate1671(.a(s_161), .O(gate486inter4));
  nand2 gate1672(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1673(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1674(.a(G1234), .O(gate486inter7));
  inv1  gate1675(.a(G1235), .O(gate486inter8));
  nand2 gate1676(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1677(.a(s_161), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1678(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1679(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1680(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1149(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1150(.a(gate489inter0), .b(s_86), .O(gate489inter1));
  and2  gate1151(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1152(.a(s_86), .O(gate489inter3));
  inv1  gate1153(.a(s_87), .O(gate489inter4));
  nand2 gate1154(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1155(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1156(.a(G1240), .O(gate489inter7));
  inv1  gate1157(.a(G1241), .O(gate489inter8));
  nand2 gate1158(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1159(.a(s_87), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1160(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1161(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1162(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1219(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1220(.a(gate493inter0), .b(s_96), .O(gate493inter1));
  and2  gate1221(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1222(.a(s_96), .O(gate493inter3));
  inv1  gate1223(.a(s_97), .O(gate493inter4));
  nand2 gate1224(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1225(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1226(.a(G1248), .O(gate493inter7));
  inv1  gate1227(.a(G1249), .O(gate493inter8));
  nand2 gate1228(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1229(.a(s_97), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1230(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1231(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1232(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate967(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate968(.a(gate496inter0), .b(s_60), .O(gate496inter1));
  and2  gate969(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate970(.a(s_60), .O(gate496inter3));
  inv1  gate971(.a(s_61), .O(gate496inter4));
  nand2 gate972(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate973(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate974(.a(G1254), .O(gate496inter7));
  inv1  gate975(.a(G1255), .O(gate496inter8));
  nand2 gate976(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate977(.a(s_61), .b(gate496inter3), .O(gate496inter10));
  nor2  gate978(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate979(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate980(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2255(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2256(.a(gate499inter0), .b(s_244), .O(gate499inter1));
  and2  gate2257(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2258(.a(s_244), .O(gate499inter3));
  inv1  gate2259(.a(s_245), .O(gate499inter4));
  nand2 gate2260(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2261(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2262(.a(G1260), .O(gate499inter7));
  inv1  gate2263(.a(G1261), .O(gate499inter8));
  nand2 gate2264(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2265(.a(s_245), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2266(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2267(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2268(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1303(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1304(.a(gate500inter0), .b(s_108), .O(gate500inter1));
  and2  gate1305(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1306(.a(s_108), .O(gate500inter3));
  inv1  gate1307(.a(s_109), .O(gate500inter4));
  nand2 gate1308(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1309(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1310(.a(G1262), .O(gate500inter7));
  inv1  gate1311(.a(G1263), .O(gate500inter8));
  nand2 gate1312(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1313(.a(s_109), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1314(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1315(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1316(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1177(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1178(.a(gate503inter0), .b(s_90), .O(gate503inter1));
  and2  gate1179(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1180(.a(s_90), .O(gate503inter3));
  inv1  gate1181(.a(s_91), .O(gate503inter4));
  nand2 gate1182(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1183(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1184(.a(G1268), .O(gate503inter7));
  inv1  gate1185(.a(G1269), .O(gate503inter8));
  nand2 gate1186(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1187(.a(s_91), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1188(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1189(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1190(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1513(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1514(.a(gate506inter0), .b(s_138), .O(gate506inter1));
  and2  gate1515(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1516(.a(s_138), .O(gate506inter3));
  inv1  gate1517(.a(s_139), .O(gate506inter4));
  nand2 gate1518(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1519(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1520(.a(G1274), .O(gate506inter7));
  inv1  gate1521(.a(G1275), .O(gate506inter8));
  nand2 gate1522(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1523(.a(s_139), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1524(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1525(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1526(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2227(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2228(.a(gate511inter0), .b(s_240), .O(gate511inter1));
  and2  gate2229(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2230(.a(s_240), .O(gate511inter3));
  inv1  gate2231(.a(s_241), .O(gate511inter4));
  nand2 gate2232(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2233(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2234(.a(G1284), .O(gate511inter7));
  inv1  gate2235(.a(G1285), .O(gate511inter8));
  nand2 gate2236(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2237(.a(s_241), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2238(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2239(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2240(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate575(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate576(.a(gate512inter0), .b(s_4), .O(gate512inter1));
  and2  gate577(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate578(.a(s_4), .O(gate512inter3));
  inv1  gate579(.a(s_5), .O(gate512inter4));
  nand2 gate580(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate581(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate582(.a(G1286), .O(gate512inter7));
  inv1  gate583(.a(G1287), .O(gate512inter8));
  nand2 gate584(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate585(.a(s_5), .b(gate512inter3), .O(gate512inter10));
  nor2  gate586(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate587(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate588(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule