module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate589(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate590(.a(gate18inter0), .b(s_6), .O(gate18inter1));
  and2  gate591(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate592(.a(s_6), .O(gate18inter3));
  inv1  gate593(.a(s_7), .O(gate18inter4));
  nand2 gate594(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate595(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate596(.a(G19), .O(gate18inter7));
  inv1  gate597(.a(G20), .O(gate18inter8));
  nand2 gate598(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate599(.a(s_7), .b(gate18inter3), .O(gate18inter10));
  nor2  gate600(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate601(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate602(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate687(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate688(.a(gate19inter0), .b(s_20), .O(gate19inter1));
  and2  gate689(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate690(.a(s_20), .O(gate19inter3));
  inv1  gate691(.a(s_21), .O(gate19inter4));
  nand2 gate692(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate693(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate694(.a(G21), .O(gate19inter7));
  inv1  gate695(.a(G22), .O(gate19inter8));
  nand2 gate696(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate697(.a(s_21), .b(gate19inter3), .O(gate19inter10));
  nor2  gate698(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate699(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate700(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1093(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1094(.a(gate37inter0), .b(s_78), .O(gate37inter1));
  and2  gate1095(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1096(.a(s_78), .O(gate37inter3));
  inv1  gate1097(.a(s_79), .O(gate37inter4));
  nand2 gate1098(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1099(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1100(.a(G19), .O(gate37inter7));
  inv1  gate1101(.a(G23), .O(gate37inter8));
  nand2 gate1102(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1103(.a(s_79), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1104(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1105(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1106(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate897(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate898(.a(gate55inter0), .b(s_50), .O(gate55inter1));
  and2  gate899(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate900(.a(s_50), .O(gate55inter3));
  inv1  gate901(.a(s_51), .O(gate55inter4));
  nand2 gate902(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate903(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate904(.a(G15), .O(gate55inter7));
  inv1  gate905(.a(G287), .O(gate55inter8));
  nand2 gate906(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate907(.a(s_51), .b(gate55inter3), .O(gate55inter10));
  nor2  gate908(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate909(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate910(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate785(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate786(.a(gate63inter0), .b(s_34), .O(gate63inter1));
  and2  gate787(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate788(.a(s_34), .O(gate63inter3));
  inv1  gate789(.a(s_35), .O(gate63inter4));
  nand2 gate790(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate791(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate792(.a(G23), .O(gate63inter7));
  inv1  gate793(.a(G299), .O(gate63inter8));
  nand2 gate794(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate795(.a(s_35), .b(gate63inter3), .O(gate63inter10));
  nor2  gate796(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate797(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate798(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1121(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1122(.a(gate67inter0), .b(s_82), .O(gate67inter1));
  and2  gate1123(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1124(.a(s_82), .O(gate67inter3));
  inv1  gate1125(.a(s_83), .O(gate67inter4));
  nand2 gate1126(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1127(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1128(.a(G27), .O(gate67inter7));
  inv1  gate1129(.a(G305), .O(gate67inter8));
  nand2 gate1130(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1131(.a(s_83), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1132(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1133(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1134(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate813(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate814(.a(gate81inter0), .b(s_38), .O(gate81inter1));
  and2  gate815(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate816(.a(s_38), .O(gate81inter3));
  inv1  gate817(.a(s_39), .O(gate81inter4));
  nand2 gate818(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate819(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate820(.a(G3), .O(gate81inter7));
  inv1  gate821(.a(G326), .O(gate81inter8));
  nand2 gate822(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate823(.a(s_39), .b(gate81inter3), .O(gate81inter10));
  nor2  gate824(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate825(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate826(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate939(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate940(.a(gate83inter0), .b(s_56), .O(gate83inter1));
  and2  gate941(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate942(.a(s_56), .O(gate83inter3));
  inv1  gate943(.a(s_57), .O(gate83inter4));
  nand2 gate944(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate945(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate946(.a(G11), .O(gate83inter7));
  inv1  gate947(.a(G329), .O(gate83inter8));
  nand2 gate948(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate949(.a(s_57), .b(gate83inter3), .O(gate83inter10));
  nor2  gate950(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate951(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate952(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate645(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate646(.a(gate87inter0), .b(s_14), .O(gate87inter1));
  and2  gate647(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate648(.a(s_14), .O(gate87inter3));
  inv1  gate649(.a(s_15), .O(gate87inter4));
  nand2 gate650(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate651(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate652(.a(G12), .O(gate87inter7));
  inv1  gate653(.a(G335), .O(gate87inter8));
  nand2 gate654(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate655(.a(s_15), .b(gate87inter3), .O(gate87inter10));
  nor2  gate656(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate657(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate658(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate729(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate730(.a(gate98inter0), .b(s_26), .O(gate98inter1));
  and2  gate731(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate732(.a(s_26), .O(gate98inter3));
  inv1  gate733(.a(s_27), .O(gate98inter4));
  nand2 gate734(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate735(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate736(.a(G23), .O(gate98inter7));
  inv1  gate737(.a(G350), .O(gate98inter8));
  nand2 gate738(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate739(.a(s_27), .b(gate98inter3), .O(gate98inter10));
  nor2  gate740(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate741(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate742(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate995(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate996(.a(gate100inter0), .b(s_64), .O(gate100inter1));
  and2  gate997(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate998(.a(s_64), .O(gate100inter3));
  inv1  gate999(.a(s_65), .O(gate100inter4));
  nand2 gate1000(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1001(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1002(.a(G31), .O(gate100inter7));
  inv1  gate1003(.a(G353), .O(gate100inter8));
  nand2 gate1004(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1005(.a(s_65), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1006(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1007(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1008(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1135(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1136(.a(gate109inter0), .b(s_84), .O(gate109inter1));
  and2  gate1137(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1138(.a(s_84), .O(gate109inter3));
  inv1  gate1139(.a(s_85), .O(gate109inter4));
  nand2 gate1140(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1141(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1142(.a(G370), .O(gate109inter7));
  inv1  gate1143(.a(G371), .O(gate109inter8));
  nand2 gate1144(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1145(.a(s_85), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1146(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1147(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1148(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate869(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate870(.a(gate111inter0), .b(s_46), .O(gate111inter1));
  and2  gate871(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate872(.a(s_46), .O(gate111inter3));
  inv1  gate873(.a(s_47), .O(gate111inter4));
  nand2 gate874(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate875(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate876(.a(G374), .O(gate111inter7));
  inv1  gate877(.a(G375), .O(gate111inter8));
  nand2 gate878(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate879(.a(s_47), .b(gate111inter3), .O(gate111inter10));
  nor2  gate880(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate881(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate882(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate953(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate954(.a(gate117inter0), .b(s_58), .O(gate117inter1));
  and2  gate955(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate956(.a(s_58), .O(gate117inter3));
  inv1  gate957(.a(s_59), .O(gate117inter4));
  nand2 gate958(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate959(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate960(.a(G386), .O(gate117inter7));
  inv1  gate961(.a(G387), .O(gate117inter8));
  nand2 gate962(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate963(.a(s_59), .b(gate117inter3), .O(gate117inter10));
  nor2  gate964(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate965(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate966(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1065(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1066(.a(gate120inter0), .b(s_74), .O(gate120inter1));
  and2  gate1067(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1068(.a(s_74), .O(gate120inter3));
  inv1  gate1069(.a(s_75), .O(gate120inter4));
  nand2 gate1070(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1071(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1072(.a(G392), .O(gate120inter7));
  inv1  gate1073(.a(G393), .O(gate120inter8));
  nand2 gate1074(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1075(.a(s_75), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1076(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1077(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1078(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate771(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate772(.a(gate134inter0), .b(s_32), .O(gate134inter1));
  and2  gate773(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate774(.a(s_32), .O(gate134inter3));
  inv1  gate775(.a(s_33), .O(gate134inter4));
  nand2 gate776(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate777(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate778(.a(G420), .O(gate134inter7));
  inv1  gate779(.a(G421), .O(gate134inter8));
  nand2 gate780(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate781(.a(s_33), .b(gate134inter3), .O(gate134inter10));
  nor2  gate782(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate783(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate784(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate967(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate968(.a(gate137inter0), .b(s_60), .O(gate137inter1));
  and2  gate969(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate970(.a(s_60), .O(gate137inter3));
  inv1  gate971(.a(s_61), .O(gate137inter4));
  nand2 gate972(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate973(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate974(.a(G426), .O(gate137inter7));
  inv1  gate975(.a(G429), .O(gate137inter8));
  nand2 gate976(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate977(.a(s_61), .b(gate137inter3), .O(gate137inter10));
  nor2  gate978(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate979(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate980(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1009(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1010(.a(gate139inter0), .b(s_66), .O(gate139inter1));
  and2  gate1011(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1012(.a(s_66), .O(gate139inter3));
  inv1  gate1013(.a(s_67), .O(gate139inter4));
  nand2 gate1014(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1015(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1016(.a(G438), .O(gate139inter7));
  inv1  gate1017(.a(G441), .O(gate139inter8));
  nand2 gate1018(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1019(.a(s_67), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1020(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1021(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1022(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate827(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate828(.a(gate157inter0), .b(s_40), .O(gate157inter1));
  and2  gate829(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate830(.a(s_40), .O(gate157inter3));
  inv1  gate831(.a(s_41), .O(gate157inter4));
  nand2 gate832(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate833(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate834(.a(G438), .O(gate157inter7));
  inv1  gate835(.a(G528), .O(gate157inter8));
  nand2 gate836(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate837(.a(s_41), .b(gate157inter3), .O(gate157inter10));
  nor2  gate838(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate839(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate840(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1023(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1024(.a(gate186inter0), .b(s_68), .O(gate186inter1));
  and2  gate1025(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1026(.a(s_68), .O(gate186inter3));
  inv1  gate1027(.a(s_69), .O(gate186inter4));
  nand2 gate1028(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1029(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1030(.a(G572), .O(gate186inter7));
  inv1  gate1031(.a(G573), .O(gate186inter8));
  nand2 gate1032(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1033(.a(s_69), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1034(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1035(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1036(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate561(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate562(.a(gate187inter0), .b(s_2), .O(gate187inter1));
  and2  gate563(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate564(.a(s_2), .O(gate187inter3));
  inv1  gate565(.a(s_3), .O(gate187inter4));
  nand2 gate566(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate567(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate568(.a(G574), .O(gate187inter7));
  inv1  gate569(.a(G575), .O(gate187inter8));
  nand2 gate570(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate571(.a(s_3), .b(gate187inter3), .O(gate187inter10));
  nor2  gate572(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate573(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate574(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1163(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1164(.a(gate193inter0), .b(s_88), .O(gate193inter1));
  and2  gate1165(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1166(.a(s_88), .O(gate193inter3));
  inv1  gate1167(.a(s_89), .O(gate193inter4));
  nand2 gate1168(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1169(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1170(.a(G586), .O(gate193inter7));
  inv1  gate1171(.a(G587), .O(gate193inter8));
  nand2 gate1172(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1173(.a(s_89), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1174(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1175(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1176(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate757(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate758(.a(gate196inter0), .b(s_30), .O(gate196inter1));
  and2  gate759(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate760(.a(s_30), .O(gate196inter3));
  inv1  gate761(.a(s_31), .O(gate196inter4));
  nand2 gate762(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate763(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate764(.a(G592), .O(gate196inter7));
  inv1  gate765(.a(G593), .O(gate196inter8));
  nand2 gate766(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate767(.a(s_31), .b(gate196inter3), .O(gate196inter10));
  nor2  gate768(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate769(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate770(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate631(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate632(.a(gate209inter0), .b(s_12), .O(gate209inter1));
  and2  gate633(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate634(.a(s_12), .O(gate209inter3));
  inv1  gate635(.a(s_13), .O(gate209inter4));
  nand2 gate636(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate637(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate638(.a(G602), .O(gate209inter7));
  inv1  gate639(.a(G666), .O(gate209inter8));
  nand2 gate640(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate641(.a(s_13), .b(gate209inter3), .O(gate209inter10));
  nor2  gate642(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate643(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate644(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate603(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate604(.a(gate223inter0), .b(s_8), .O(gate223inter1));
  and2  gate605(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate606(.a(s_8), .O(gate223inter3));
  inv1  gate607(.a(s_9), .O(gate223inter4));
  nand2 gate608(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate609(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate610(.a(G627), .O(gate223inter7));
  inv1  gate611(.a(G687), .O(gate223inter8));
  nand2 gate612(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate613(.a(s_9), .b(gate223inter3), .O(gate223inter10));
  nor2  gate614(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate615(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate616(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate925(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate926(.a(gate225inter0), .b(s_54), .O(gate225inter1));
  and2  gate927(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate928(.a(s_54), .O(gate225inter3));
  inv1  gate929(.a(s_55), .O(gate225inter4));
  nand2 gate930(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate931(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate932(.a(G690), .O(gate225inter7));
  inv1  gate933(.a(G691), .O(gate225inter8));
  nand2 gate934(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate935(.a(s_55), .b(gate225inter3), .O(gate225inter10));
  nor2  gate936(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate937(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate938(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate617(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate618(.a(gate228inter0), .b(s_10), .O(gate228inter1));
  and2  gate619(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate620(.a(s_10), .O(gate228inter3));
  inv1  gate621(.a(s_11), .O(gate228inter4));
  nand2 gate622(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate623(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate624(.a(G696), .O(gate228inter7));
  inv1  gate625(.a(G697), .O(gate228inter8));
  nand2 gate626(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate627(.a(s_11), .b(gate228inter3), .O(gate228inter10));
  nor2  gate628(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate629(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate630(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate799(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate800(.a(gate232inter0), .b(s_36), .O(gate232inter1));
  and2  gate801(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate802(.a(s_36), .O(gate232inter3));
  inv1  gate803(.a(s_37), .O(gate232inter4));
  nand2 gate804(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate805(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate806(.a(G704), .O(gate232inter7));
  inv1  gate807(.a(G705), .O(gate232inter8));
  nand2 gate808(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate809(.a(s_37), .b(gate232inter3), .O(gate232inter10));
  nor2  gate810(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate811(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate812(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1079(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1080(.a(gate253inter0), .b(s_76), .O(gate253inter1));
  and2  gate1081(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1082(.a(s_76), .O(gate253inter3));
  inv1  gate1083(.a(s_77), .O(gate253inter4));
  nand2 gate1084(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1085(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1086(.a(G260), .O(gate253inter7));
  inv1  gate1087(.a(G748), .O(gate253inter8));
  nand2 gate1088(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1089(.a(s_77), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1090(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1091(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1092(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate673(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate674(.a(gate256inter0), .b(s_18), .O(gate256inter1));
  and2  gate675(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate676(.a(s_18), .O(gate256inter3));
  inv1  gate677(.a(s_19), .O(gate256inter4));
  nand2 gate678(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate679(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate680(.a(G715), .O(gate256inter7));
  inv1  gate681(.a(G751), .O(gate256inter8));
  nand2 gate682(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate683(.a(s_19), .b(gate256inter3), .O(gate256inter10));
  nor2  gate684(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate685(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate686(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1051(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1052(.a(gate267inter0), .b(s_72), .O(gate267inter1));
  and2  gate1053(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1054(.a(s_72), .O(gate267inter3));
  inv1  gate1055(.a(s_73), .O(gate267inter4));
  nand2 gate1056(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1057(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1058(.a(G648), .O(gate267inter7));
  inv1  gate1059(.a(G776), .O(gate267inter8));
  nand2 gate1060(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1061(.a(s_73), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1062(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1063(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1064(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate743(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate744(.a(gate274inter0), .b(s_28), .O(gate274inter1));
  and2  gate745(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate746(.a(s_28), .O(gate274inter3));
  inv1  gate747(.a(s_29), .O(gate274inter4));
  nand2 gate748(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate749(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate750(.a(G770), .O(gate274inter7));
  inv1  gate751(.a(G794), .O(gate274inter8));
  nand2 gate752(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate753(.a(s_29), .b(gate274inter3), .O(gate274inter10));
  nor2  gate754(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate755(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate756(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate855(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate856(.a(gate290inter0), .b(s_44), .O(gate290inter1));
  and2  gate857(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate858(.a(s_44), .O(gate290inter3));
  inv1  gate859(.a(s_45), .O(gate290inter4));
  nand2 gate860(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate861(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate862(.a(G820), .O(gate290inter7));
  inv1  gate863(.a(G821), .O(gate290inter8));
  nand2 gate864(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate865(.a(s_45), .b(gate290inter3), .O(gate290inter10));
  nor2  gate866(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate867(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate868(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate701(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate702(.a(gate291inter0), .b(s_22), .O(gate291inter1));
  and2  gate703(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate704(.a(s_22), .O(gate291inter3));
  inv1  gate705(.a(s_23), .O(gate291inter4));
  nand2 gate706(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate707(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate708(.a(G822), .O(gate291inter7));
  inv1  gate709(.a(G823), .O(gate291inter8));
  nand2 gate710(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate711(.a(s_23), .b(gate291inter3), .O(gate291inter10));
  nor2  gate712(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate713(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate714(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate547(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate548(.a(gate403inter0), .b(s_0), .O(gate403inter1));
  and2  gate549(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate550(.a(s_0), .O(gate403inter3));
  inv1  gate551(.a(s_1), .O(gate403inter4));
  nand2 gate552(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate553(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate554(.a(G17), .O(gate403inter7));
  inv1  gate555(.a(G1084), .O(gate403inter8));
  nand2 gate556(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate557(.a(s_1), .b(gate403inter3), .O(gate403inter10));
  nor2  gate558(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate559(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate560(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate659(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate660(.a(gate408inter0), .b(s_16), .O(gate408inter1));
  and2  gate661(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate662(.a(s_16), .O(gate408inter3));
  inv1  gate663(.a(s_17), .O(gate408inter4));
  nand2 gate664(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate665(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate666(.a(G22), .O(gate408inter7));
  inv1  gate667(.a(G1099), .O(gate408inter8));
  nand2 gate668(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate669(.a(s_17), .b(gate408inter3), .O(gate408inter10));
  nor2  gate670(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate671(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate672(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1037(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1038(.a(gate410inter0), .b(s_70), .O(gate410inter1));
  and2  gate1039(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1040(.a(s_70), .O(gate410inter3));
  inv1  gate1041(.a(s_71), .O(gate410inter4));
  nand2 gate1042(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1043(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1044(.a(G24), .O(gate410inter7));
  inv1  gate1045(.a(G1105), .O(gate410inter8));
  nand2 gate1046(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1047(.a(s_71), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1048(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1049(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1050(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate981(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate982(.a(gate439inter0), .b(s_62), .O(gate439inter1));
  and2  gate983(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate984(.a(s_62), .O(gate439inter3));
  inv1  gate985(.a(s_63), .O(gate439inter4));
  nand2 gate986(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate987(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate988(.a(G11), .O(gate439inter7));
  inv1  gate989(.a(G1162), .O(gate439inter8));
  nand2 gate990(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate991(.a(s_63), .b(gate439inter3), .O(gate439inter10));
  nor2  gate992(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate993(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate994(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate883(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate884(.a(gate443inter0), .b(s_48), .O(gate443inter1));
  and2  gate885(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate886(.a(s_48), .O(gate443inter3));
  inv1  gate887(.a(s_49), .O(gate443inter4));
  nand2 gate888(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate889(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate890(.a(G13), .O(gate443inter7));
  inv1  gate891(.a(G1168), .O(gate443inter8));
  nand2 gate892(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate893(.a(s_49), .b(gate443inter3), .O(gate443inter10));
  nor2  gate894(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate895(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate896(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate715(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate716(.a(gate447inter0), .b(s_24), .O(gate447inter1));
  and2  gate717(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate718(.a(s_24), .O(gate447inter3));
  inv1  gate719(.a(s_25), .O(gate447inter4));
  nand2 gate720(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate721(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate722(.a(G15), .O(gate447inter7));
  inv1  gate723(.a(G1174), .O(gate447inter8));
  nand2 gate724(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate725(.a(s_25), .b(gate447inter3), .O(gate447inter10));
  nor2  gate726(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate727(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate728(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1107(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1108(.a(gate458inter0), .b(s_80), .O(gate458inter1));
  and2  gate1109(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1110(.a(s_80), .O(gate458inter3));
  inv1  gate1111(.a(s_81), .O(gate458inter4));
  nand2 gate1112(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1113(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1114(.a(G1093), .O(gate458inter7));
  inv1  gate1115(.a(G1189), .O(gate458inter8));
  nand2 gate1116(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1117(.a(s_81), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1118(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1119(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1120(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate575(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate576(.a(gate463inter0), .b(s_4), .O(gate463inter1));
  and2  gate577(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate578(.a(s_4), .O(gate463inter3));
  inv1  gate579(.a(s_5), .O(gate463inter4));
  nand2 gate580(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate581(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate582(.a(G23), .O(gate463inter7));
  inv1  gate583(.a(G1198), .O(gate463inter8));
  nand2 gate584(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate585(.a(s_5), .b(gate463inter3), .O(gate463inter10));
  nor2  gate586(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate587(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate588(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1149(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1150(.a(gate480inter0), .b(s_86), .O(gate480inter1));
  and2  gate1151(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1152(.a(s_86), .O(gate480inter3));
  inv1  gate1153(.a(s_87), .O(gate480inter4));
  nand2 gate1154(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1155(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1156(.a(G1126), .O(gate480inter7));
  inv1  gate1157(.a(G1222), .O(gate480inter8));
  nand2 gate1158(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1159(.a(s_87), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1160(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1161(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1162(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1177(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1178(.a(gate487inter0), .b(s_90), .O(gate487inter1));
  and2  gate1179(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1180(.a(s_90), .O(gate487inter3));
  inv1  gate1181(.a(s_91), .O(gate487inter4));
  nand2 gate1182(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1183(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1184(.a(G1236), .O(gate487inter7));
  inv1  gate1185(.a(G1237), .O(gate487inter8));
  nand2 gate1186(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1187(.a(s_91), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1188(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1189(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1190(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate911(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate912(.a(gate501inter0), .b(s_52), .O(gate501inter1));
  and2  gate913(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate914(.a(s_52), .O(gate501inter3));
  inv1  gate915(.a(s_53), .O(gate501inter4));
  nand2 gate916(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate917(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate918(.a(G1264), .O(gate501inter7));
  inv1  gate919(.a(G1265), .O(gate501inter8));
  nand2 gate920(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate921(.a(s_53), .b(gate501inter3), .O(gate501inter10));
  nor2  gate922(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate923(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate924(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate841(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate842(.a(gate503inter0), .b(s_42), .O(gate503inter1));
  and2  gate843(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate844(.a(s_42), .O(gate503inter3));
  inv1  gate845(.a(s_43), .O(gate503inter4));
  nand2 gate846(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate847(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate848(.a(G1268), .O(gate503inter7));
  inv1  gate849(.a(G1269), .O(gate503inter8));
  nand2 gate850(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate851(.a(s_43), .b(gate503inter3), .O(gate503inter10));
  nor2  gate852(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate853(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate854(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule