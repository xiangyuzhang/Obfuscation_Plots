module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate617(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate618(.a(gate16inter0), .b(s_10), .O(gate16inter1));
  and2  gate619(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate620(.a(s_10), .O(gate16inter3));
  inv1  gate621(.a(s_11), .O(gate16inter4));
  nand2 gate622(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate623(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate624(.a(G15), .O(gate16inter7));
  inv1  gate625(.a(G16), .O(gate16inter8));
  nand2 gate626(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate627(.a(s_11), .b(gate16inter3), .O(gate16inter10));
  nor2  gate628(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate629(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate630(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate659(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate660(.a(gate17inter0), .b(s_16), .O(gate17inter1));
  and2  gate661(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate662(.a(s_16), .O(gate17inter3));
  inv1  gate663(.a(s_17), .O(gate17inter4));
  nand2 gate664(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate665(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate666(.a(G17), .O(gate17inter7));
  inv1  gate667(.a(G18), .O(gate17inter8));
  nand2 gate668(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate669(.a(s_17), .b(gate17inter3), .O(gate17inter10));
  nor2  gate670(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate671(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate672(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate729(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate730(.a(gate19inter0), .b(s_26), .O(gate19inter1));
  and2  gate731(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate732(.a(s_26), .O(gate19inter3));
  inv1  gate733(.a(s_27), .O(gate19inter4));
  nand2 gate734(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate735(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate736(.a(G21), .O(gate19inter7));
  inv1  gate737(.a(G22), .O(gate19inter8));
  nand2 gate738(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate739(.a(s_27), .b(gate19inter3), .O(gate19inter10));
  nor2  gate740(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate741(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate742(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1513(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1514(.a(gate24inter0), .b(s_138), .O(gate24inter1));
  and2  gate1515(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1516(.a(s_138), .O(gate24inter3));
  inv1  gate1517(.a(s_139), .O(gate24inter4));
  nand2 gate1518(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1519(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1520(.a(G31), .O(gate24inter7));
  inv1  gate1521(.a(G32), .O(gate24inter8));
  nand2 gate1522(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1523(.a(s_139), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1524(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1525(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1526(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate561(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate562(.a(gate27inter0), .b(s_2), .O(gate27inter1));
  and2  gate563(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate564(.a(s_2), .O(gate27inter3));
  inv1  gate565(.a(s_3), .O(gate27inter4));
  nand2 gate566(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate567(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate568(.a(G2), .O(gate27inter7));
  inv1  gate569(.a(G6), .O(gate27inter8));
  nand2 gate570(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate571(.a(s_3), .b(gate27inter3), .O(gate27inter10));
  nor2  gate572(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate573(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate574(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate631(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate632(.a(gate33inter0), .b(s_12), .O(gate33inter1));
  and2  gate633(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate634(.a(s_12), .O(gate33inter3));
  inv1  gate635(.a(s_13), .O(gate33inter4));
  nand2 gate636(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate637(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate638(.a(G17), .O(gate33inter7));
  inv1  gate639(.a(G21), .O(gate33inter8));
  nand2 gate640(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate641(.a(s_13), .b(gate33inter3), .O(gate33inter10));
  nor2  gate642(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate643(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate644(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1527(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1528(.a(gate37inter0), .b(s_140), .O(gate37inter1));
  and2  gate1529(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1530(.a(s_140), .O(gate37inter3));
  inv1  gate1531(.a(s_141), .O(gate37inter4));
  nand2 gate1532(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1533(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1534(.a(G19), .O(gate37inter7));
  inv1  gate1535(.a(G23), .O(gate37inter8));
  nand2 gate1536(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1537(.a(s_141), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1538(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1539(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1540(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1345(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1346(.a(gate38inter0), .b(s_114), .O(gate38inter1));
  and2  gate1347(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1348(.a(s_114), .O(gate38inter3));
  inv1  gate1349(.a(s_115), .O(gate38inter4));
  nand2 gate1350(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1351(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1352(.a(G27), .O(gate38inter7));
  inv1  gate1353(.a(G31), .O(gate38inter8));
  nand2 gate1354(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1355(.a(s_115), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1356(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1357(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1358(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate757(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate758(.a(gate44inter0), .b(s_30), .O(gate44inter1));
  and2  gate759(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate760(.a(s_30), .O(gate44inter3));
  inv1  gate761(.a(s_31), .O(gate44inter4));
  nand2 gate762(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate763(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate764(.a(G4), .O(gate44inter7));
  inv1  gate765(.a(G269), .O(gate44inter8));
  nand2 gate766(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate767(.a(s_31), .b(gate44inter3), .O(gate44inter10));
  nor2  gate768(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate769(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate770(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate967(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate968(.a(gate54inter0), .b(s_60), .O(gate54inter1));
  and2  gate969(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate970(.a(s_60), .O(gate54inter3));
  inv1  gate971(.a(s_61), .O(gate54inter4));
  nand2 gate972(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate973(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate974(.a(G14), .O(gate54inter7));
  inv1  gate975(.a(G284), .O(gate54inter8));
  nand2 gate976(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate977(.a(s_61), .b(gate54inter3), .O(gate54inter10));
  nor2  gate978(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate979(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate980(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate603(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate604(.a(gate59inter0), .b(s_8), .O(gate59inter1));
  and2  gate605(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate606(.a(s_8), .O(gate59inter3));
  inv1  gate607(.a(s_9), .O(gate59inter4));
  nand2 gate608(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate609(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate610(.a(G19), .O(gate59inter7));
  inv1  gate611(.a(G293), .O(gate59inter8));
  nand2 gate612(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate613(.a(s_9), .b(gate59inter3), .O(gate59inter10));
  nor2  gate614(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate615(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate616(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate897(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate898(.a(gate66inter0), .b(s_50), .O(gate66inter1));
  and2  gate899(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate900(.a(s_50), .O(gate66inter3));
  inv1  gate901(.a(s_51), .O(gate66inter4));
  nand2 gate902(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate903(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate904(.a(G26), .O(gate66inter7));
  inv1  gate905(.a(G302), .O(gate66inter8));
  nand2 gate906(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate907(.a(s_51), .b(gate66inter3), .O(gate66inter10));
  nor2  gate908(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate909(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate910(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1373(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1374(.a(gate68inter0), .b(s_118), .O(gate68inter1));
  and2  gate1375(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1376(.a(s_118), .O(gate68inter3));
  inv1  gate1377(.a(s_119), .O(gate68inter4));
  nand2 gate1378(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1379(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1380(.a(G28), .O(gate68inter7));
  inv1  gate1381(.a(G305), .O(gate68inter8));
  nand2 gate1382(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1383(.a(s_119), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1384(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1385(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1386(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1191(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1192(.a(gate73inter0), .b(s_92), .O(gate73inter1));
  and2  gate1193(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1194(.a(s_92), .O(gate73inter3));
  inv1  gate1195(.a(s_93), .O(gate73inter4));
  nand2 gate1196(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1197(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1198(.a(G1), .O(gate73inter7));
  inv1  gate1199(.a(G314), .O(gate73inter8));
  nand2 gate1200(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1201(.a(s_93), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1202(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1203(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1204(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate687(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate688(.a(gate80inter0), .b(s_20), .O(gate80inter1));
  and2  gate689(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate690(.a(s_20), .O(gate80inter3));
  inv1  gate691(.a(s_21), .O(gate80inter4));
  nand2 gate692(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate693(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate694(.a(G14), .O(gate80inter7));
  inv1  gate695(.a(G323), .O(gate80inter8));
  nand2 gate696(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate697(.a(s_21), .b(gate80inter3), .O(gate80inter10));
  nor2  gate698(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate699(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate700(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate673(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate674(.a(gate88inter0), .b(s_18), .O(gate88inter1));
  and2  gate675(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate676(.a(s_18), .O(gate88inter3));
  inv1  gate677(.a(s_19), .O(gate88inter4));
  nand2 gate678(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate679(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate680(.a(G16), .O(gate88inter7));
  inv1  gate681(.a(G335), .O(gate88inter8));
  nand2 gate682(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate683(.a(s_19), .b(gate88inter3), .O(gate88inter10));
  nor2  gate684(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate685(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate686(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate575(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate576(.a(gate94inter0), .b(s_4), .O(gate94inter1));
  and2  gate577(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate578(.a(s_4), .O(gate94inter3));
  inv1  gate579(.a(s_5), .O(gate94inter4));
  nand2 gate580(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate581(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate582(.a(G22), .O(gate94inter7));
  inv1  gate583(.a(G344), .O(gate94inter8));
  nand2 gate584(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate585(.a(s_5), .b(gate94inter3), .O(gate94inter10));
  nor2  gate586(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate587(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate588(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1429(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1430(.a(gate96inter0), .b(s_126), .O(gate96inter1));
  and2  gate1431(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1432(.a(s_126), .O(gate96inter3));
  inv1  gate1433(.a(s_127), .O(gate96inter4));
  nand2 gate1434(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1435(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1436(.a(G30), .O(gate96inter7));
  inv1  gate1437(.a(G347), .O(gate96inter8));
  nand2 gate1438(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1439(.a(s_127), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1440(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1441(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1442(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1219(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1220(.a(gate105inter0), .b(s_96), .O(gate105inter1));
  and2  gate1221(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1222(.a(s_96), .O(gate105inter3));
  inv1  gate1223(.a(s_97), .O(gate105inter4));
  nand2 gate1224(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1225(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1226(.a(G362), .O(gate105inter7));
  inv1  gate1227(.a(G363), .O(gate105inter8));
  nand2 gate1228(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1229(.a(s_97), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1230(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1231(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1232(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1247(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1248(.a(gate111inter0), .b(s_100), .O(gate111inter1));
  and2  gate1249(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1250(.a(s_100), .O(gate111inter3));
  inv1  gate1251(.a(s_101), .O(gate111inter4));
  nand2 gate1252(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1253(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1254(.a(G374), .O(gate111inter7));
  inv1  gate1255(.a(G375), .O(gate111inter8));
  nand2 gate1256(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1257(.a(s_101), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1258(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1259(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1260(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1149(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1150(.a(gate115inter0), .b(s_86), .O(gate115inter1));
  and2  gate1151(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1152(.a(s_86), .O(gate115inter3));
  inv1  gate1153(.a(s_87), .O(gate115inter4));
  nand2 gate1154(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1155(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1156(.a(G382), .O(gate115inter7));
  inv1  gate1157(.a(G383), .O(gate115inter8));
  nand2 gate1158(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1159(.a(s_87), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1160(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1161(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1162(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate785(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate786(.a(gate125inter0), .b(s_34), .O(gate125inter1));
  and2  gate787(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate788(.a(s_34), .O(gate125inter3));
  inv1  gate789(.a(s_35), .O(gate125inter4));
  nand2 gate790(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate791(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate792(.a(G402), .O(gate125inter7));
  inv1  gate793(.a(G403), .O(gate125inter8));
  nand2 gate794(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate795(.a(s_35), .b(gate125inter3), .O(gate125inter10));
  nor2  gate796(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate797(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate798(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1289(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1290(.a(gate126inter0), .b(s_106), .O(gate126inter1));
  and2  gate1291(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1292(.a(s_106), .O(gate126inter3));
  inv1  gate1293(.a(s_107), .O(gate126inter4));
  nand2 gate1294(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1295(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1296(.a(G404), .O(gate126inter7));
  inv1  gate1297(.a(G405), .O(gate126inter8));
  nand2 gate1298(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1299(.a(s_107), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1300(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1301(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1302(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1499(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1500(.a(gate129inter0), .b(s_136), .O(gate129inter1));
  and2  gate1501(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1502(.a(s_136), .O(gate129inter3));
  inv1  gate1503(.a(s_137), .O(gate129inter4));
  nand2 gate1504(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1505(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1506(.a(G410), .O(gate129inter7));
  inv1  gate1507(.a(G411), .O(gate129inter8));
  nand2 gate1508(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1509(.a(s_137), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1510(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1511(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1512(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1485(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1486(.a(gate131inter0), .b(s_134), .O(gate131inter1));
  and2  gate1487(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1488(.a(s_134), .O(gate131inter3));
  inv1  gate1489(.a(s_135), .O(gate131inter4));
  nand2 gate1490(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1491(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1492(.a(G414), .O(gate131inter7));
  inv1  gate1493(.a(G415), .O(gate131inter8));
  nand2 gate1494(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1495(.a(s_135), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1496(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1497(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1498(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1331(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1332(.a(gate134inter0), .b(s_112), .O(gate134inter1));
  and2  gate1333(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1334(.a(s_112), .O(gate134inter3));
  inv1  gate1335(.a(s_113), .O(gate134inter4));
  nand2 gate1336(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1337(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1338(.a(G420), .O(gate134inter7));
  inv1  gate1339(.a(G421), .O(gate134inter8));
  nand2 gate1340(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1341(.a(s_113), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1342(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1343(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1344(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1359(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1360(.a(gate137inter0), .b(s_116), .O(gate137inter1));
  and2  gate1361(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1362(.a(s_116), .O(gate137inter3));
  inv1  gate1363(.a(s_117), .O(gate137inter4));
  nand2 gate1364(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1365(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1366(.a(G426), .O(gate137inter7));
  inv1  gate1367(.a(G429), .O(gate137inter8));
  nand2 gate1368(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1369(.a(s_117), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1370(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1371(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1372(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate715(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate716(.a(gate141inter0), .b(s_24), .O(gate141inter1));
  and2  gate717(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate718(.a(s_24), .O(gate141inter3));
  inv1  gate719(.a(s_25), .O(gate141inter4));
  nand2 gate720(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate721(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate722(.a(G450), .O(gate141inter7));
  inv1  gate723(.a(G453), .O(gate141inter8));
  nand2 gate724(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate725(.a(s_25), .b(gate141inter3), .O(gate141inter10));
  nor2  gate726(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate727(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate728(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1107(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1108(.a(gate155inter0), .b(s_80), .O(gate155inter1));
  and2  gate1109(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1110(.a(s_80), .O(gate155inter3));
  inv1  gate1111(.a(s_81), .O(gate155inter4));
  nand2 gate1112(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1113(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1114(.a(G432), .O(gate155inter7));
  inv1  gate1115(.a(G525), .O(gate155inter8));
  nand2 gate1116(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1117(.a(s_81), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1118(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1119(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1120(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate981(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate982(.a(gate156inter0), .b(s_62), .O(gate156inter1));
  and2  gate983(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate984(.a(s_62), .O(gate156inter3));
  inv1  gate985(.a(s_63), .O(gate156inter4));
  nand2 gate986(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate987(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate988(.a(G435), .O(gate156inter7));
  inv1  gate989(.a(G525), .O(gate156inter8));
  nand2 gate990(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate991(.a(s_63), .b(gate156inter3), .O(gate156inter10));
  nor2  gate992(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate993(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate994(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate911(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate912(.a(gate157inter0), .b(s_52), .O(gate157inter1));
  and2  gate913(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate914(.a(s_52), .O(gate157inter3));
  inv1  gate915(.a(s_53), .O(gate157inter4));
  nand2 gate916(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate917(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate918(.a(G438), .O(gate157inter7));
  inv1  gate919(.a(G528), .O(gate157inter8));
  nand2 gate920(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate921(.a(s_53), .b(gate157inter3), .O(gate157inter10));
  nor2  gate922(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate923(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate924(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate799(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate800(.a(gate158inter0), .b(s_36), .O(gate158inter1));
  and2  gate801(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate802(.a(s_36), .O(gate158inter3));
  inv1  gate803(.a(s_37), .O(gate158inter4));
  nand2 gate804(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate805(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate806(.a(G441), .O(gate158inter7));
  inv1  gate807(.a(G528), .O(gate158inter8));
  nand2 gate808(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate809(.a(s_37), .b(gate158inter3), .O(gate158inter10));
  nor2  gate810(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate811(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate812(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1177(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1178(.a(gate159inter0), .b(s_90), .O(gate159inter1));
  and2  gate1179(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1180(.a(s_90), .O(gate159inter3));
  inv1  gate1181(.a(s_91), .O(gate159inter4));
  nand2 gate1182(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1183(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1184(.a(G444), .O(gate159inter7));
  inv1  gate1185(.a(G531), .O(gate159inter8));
  nand2 gate1186(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1187(.a(s_91), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1188(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1189(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1190(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1009(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1010(.a(gate165inter0), .b(s_66), .O(gate165inter1));
  and2  gate1011(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1012(.a(s_66), .O(gate165inter3));
  inv1  gate1013(.a(s_67), .O(gate165inter4));
  nand2 gate1014(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1015(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1016(.a(G462), .O(gate165inter7));
  inv1  gate1017(.a(G540), .O(gate165inter8));
  nand2 gate1018(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1019(.a(s_67), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1020(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1021(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1022(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate589(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate590(.a(gate168inter0), .b(s_6), .O(gate168inter1));
  and2  gate591(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate592(.a(s_6), .O(gate168inter3));
  inv1  gate593(.a(s_7), .O(gate168inter4));
  nand2 gate594(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate595(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate596(.a(G471), .O(gate168inter7));
  inv1  gate597(.a(G543), .O(gate168inter8));
  nand2 gate598(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate599(.a(s_7), .b(gate168inter3), .O(gate168inter10));
  nor2  gate600(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate601(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate602(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1135(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1136(.a(gate170inter0), .b(s_84), .O(gate170inter1));
  and2  gate1137(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1138(.a(s_84), .O(gate170inter3));
  inv1  gate1139(.a(s_85), .O(gate170inter4));
  nand2 gate1140(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1141(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1142(.a(G477), .O(gate170inter7));
  inv1  gate1143(.a(G546), .O(gate170inter8));
  nand2 gate1144(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1145(.a(s_85), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1146(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1147(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1148(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1415(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1416(.a(gate181inter0), .b(s_124), .O(gate181inter1));
  and2  gate1417(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1418(.a(s_124), .O(gate181inter3));
  inv1  gate1419(.a(s_125), .O(gate181inter4));
  nand2 gate1420(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1421(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1422(.a(G510), .O(gate181inter7));
  inv1  gate1423(.a(G564), .O(gate181inter8));
  nand2 gate1424(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1425(.a(s_125), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1426(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1427(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1428(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1275(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1276(.a(gate184inter0), .b(s_104), .O(gate184inter1));
  and2  gate1277(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1278(.a(s_104), .O(gate184inter3));
  inv1  gate1279(.a(s_105), .O(gate184inter4));
  nand2 gate1280(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1281(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1282(.a(G519), .O(gate184inter7));
  inv1  gate1283(.a(G567), .O(gate184inter8));
  nand2 gate1284(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1285(.a(s_105), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1286(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1287(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1288(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate925(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate926(.a(gate190inter0), .b(s_54), .O(gate190inter1));
  and2  gate927(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate928(.a(s_54), .O(gate190inter3));
  inv1  gate929(.a(s_55), .O(gate190inter4));
  nand2 gate930(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate931(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate932(.a(G580), .O(gate190inter7));
  inv1  gate933(.a(G581), .O(gate190inter8));
  nand2 gate934(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate935(.a(s_55), .b(gate190inter3), .O(gate190inter10));
  nor2  gate936(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate937(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate938(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1387(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1388(.a(gate196inter0), .b(s_120), .O(gate196inter1));
  and2  gate1389(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1390(.a(s_120), .O(gate196inter3));
  inv1  gate1391(.a(s_121), .O(gate196inter4));
  nand2 gate1392(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1393(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1394(.a(G592), .O(gate196inter7));
  inv1  gate1395(.a(G593), .O(gate196inter8));
  nand2 gate1396(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1397(.a(s_121), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1398(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1399(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1400(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1093(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1094(.a(gate201inter0), .b(s_78), .O(gate201inter1));
  and2  gate1095(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1096(.a(s_78), .O(gate201inter3));
  inv1  gate1097(.a(s_79), .O(gate201inter4));
  nand2 gate1098(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1099(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1100(.a(G602), .O(gate201inter7));
  inv1  gate1101(.a(G607), .O(gate201inter8));
  nand2 gate1102(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1103(.a(s_79), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1104(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1105(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1106(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1233(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1234(.a(gate206inter0), .b(s_98), .O(gate206inter1));
  and2  gate1235(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1236(.a(s_98), .O(gate206inter3));
  inv1  gate1237(.a(s_99), .O(gate206inter4));
  nand2 gate1238(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1239(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1240(.a(G632), .O(gate206inter7));
  inv1  gate1241(.a(G637), .O(gate206inter8));
  nand2 gate1242(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1243(.a(s_99), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1244(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1245(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1246(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1471(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1472(.a(gate209inter0), .b(s_132), .O(gate209inter1));
  and2  gate1473(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1474(.a(s_132), .O(gate209inter3));
  inv1  gate1475(.a(s_133), .O(gate209inter4));
  nand2 gate1476(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1477(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1478(.a(G602), .O(gate209inter7));
  inv1  gate1479(.a(G666), .O(gate209inter8));
  nand2 gate1480(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1481(.a(s_133), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1482(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1483(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1484(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1037(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1038(.a(gate212inter0), .b(s_70), .O(gate212inter1));
  and2  gate1039(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1040(.a(s_70), .O(gate212inter3));
  inv1  gate1041(.a(s_71), .O(gate212inter4));
  nand2 gate1042(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1043(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1044(.a(G617), .O(gate212inter7));
  inv1  gate1045(.a(G669), .O(gate212inter8));
  nand2 gate1046(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1047(.a(s_71), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1048(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1049(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1050(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate645(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate646(.a(gate214inter0), .b(s_14), .O(gate214inter1));
  and2  gate647(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate648(.a(s_14), .O(gate214inter3));
  inv1  gate649(.a(s_15), .O(gate214inter4));
  nand2 gate650(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate651(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate652(.a(G612), .O(gate214inter7));
  inv1  gate653(.a(G672), .O(gate214inter8));
  nand2 gate654(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate655(.a(s_15), .b(gate214inter3), .O(gate214inter10));
  nor2  gate656(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate657(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate658(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate701(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate702(.a(gate231inter0), .b(s_22), .O(gate231inter1));
  and2  gate703(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate704(.a(s_22), .O(gate231inter3));
  inv1  gate705(.a(s_23), .O(gate231inter4));
  nand2 gate706(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate707(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate708(.a(G702), .O(gate231inter7));
  inv1  gate709(.a(G703), .O(gate231inter8));
  nand2 gate710(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate711(.a(s_23), .b(gate231inter3), .O(gate231inter10));
  nor2  gate712(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate713(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate714(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1023(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1024(.a(gate232inter0), .b(s_68), .O(gate232inter1));
  and2  gate1025(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1026(.a(s_68), .O(gate232inter3));
  inv1  gate1027(.a(s_69), .O(gate232inter4));
  nand2 gate1028(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1029(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1030(.a(G704), .O(gate232inter7));
  inv1  gate1031(.a(G705), .O(gate232inter8));
  nand2 gate1032(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1033(.a(s_69), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1034(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1035(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1036(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1205(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1206(.a(gate242inter0), .b(s_94), .O(gate242inter1));
  and2  gate1207(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1208(.a(s_94), .O(gate242inter3));
  inv1  gate1209(.a(s_95), .O(gate242inter4));
  nand2 gate1210(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1211(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1212(.a(G718), .O(gate242inter7));
  inv1  gate1213(.a(G730), .O(gate242inter8));
  nand2 gate1214(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1215(.a(s_95), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1216(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1217(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1218(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1065(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1066(.a(gate244inter0), .b(s_74), .O(gate244inter1));
  and2  gate1067(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1068(.a(s_74), .O(gate244inter3));
  inv1  gate1069(.a(s_75), .O(gate244inter4));
  nand2 gate1070(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1071(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1072(.a(G721), .O(gate244inter7));
  inv1  gate1073(.a(G733), .O(gate244inter8));
  nand2 gate1074(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1075(.a(s_75), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1076(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1077(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1078(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate827(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate828(.a(gate253inter0), .b(s_40), .O(gate253inter1));
  and2  gate829(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate830(.a(s_40), .O(gate253inter3));
  inv1  gate831(.a(s_41), .O(gate253inter4));
  nand2 gate832(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate833(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate834(.a(G260), .O(gate253inter7));
  inv1  gate835(.a(G748), .O(gate253inter8));
  nand2 gate836(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate837(.a(s_41), .b(gate253inter3), .O(gate253inter10));
  nor2  gate838(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate839(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate840(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1261(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1262(.a(gate255inter0), .b(s_102), .O(gate255inter1));
  and2  gate1263(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1264(.a(s_102), .O(gate255inter3));
  inv1  gate1265(.a(s_103), .O(gate255inter4));
  nand2 gate1266(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1267(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1268(.a(G263), .O(gate255inter7));
  inv1  gate1269(.a(G751), .O(gate255inter8));
  nand2 gate1270(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1271(.a(s_103), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1272(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1273(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1274(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate813(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate814(.a(gate258inter0), .b(s_38), .O(gate258inter1));
  and2  gate815(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate816(.a(s_38), .O(gate258inter3));
  inv1  gate817(.a(s_39), .O(gate258inter4));
  nand2 gate818(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate819(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate820(.a(G756), .O(gate258inter7));
  inv1  gate821(.a(G757), .O(gate258inter8));
  nand2 gate822(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate823(.a(s_39), .b(gate258inter3), .O(gate258inter10));
  nor2  gate824(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate825(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate826(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1443(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1444(.a(gate263inter0), .b(s_128), .O(gate263inter1));
  and2  gate1445(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1446(.a(s_128), .O(gate263inter3));
  inv1  gate1447(.a(s_129), .O(gate263inter4));
  nand2 gate1448(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1449(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1450(.a(G766), .O(gate263inter7));
  inv1  gate1451(.a(G767), .O(gate263inter8));
  nand2 gate1452(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1453(.a(s_129), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1454(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1455(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1456(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate743(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate744(.a(gate267inter0), .b(s_28), .O(gate267inter1));
  and2  gate745(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate746(.a(s_28), .O(gate267inter3));
  inv1  gate747(.a(s_29), .O(gate267inter4));
  nand2 gate748(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate749(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate750(.a(G648), .O(gate267inter7));
  inv1  gate751(.a(G776), .O(gate267inter8));
  nand2 gate752(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate753(.a(s_29), .b(gate267inter3), .O(gate267inter10));
  nor2  gate754(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate755(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate756(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1317(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1318(.a(gate274inter0), .b(s_110), .O(gate274inter1));
  and2  gate1319(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1320(.a(s_110), .O(gate274inter3));
  inv1  gate1321(.a(s_111), .O(gate274inter4));
  nand2 gate1322(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1323(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1324(.a(G770), .O(gate274inter7));
  inv1  gate1325(.a(G794), .O(gate274inter8));
  nand2 gate1326(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1327(.a(s_111), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1328(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1329(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1330(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1051(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1052(.a(gate279inter0), .b(s_72), .O(gate279inter1));
  and2  gate1053(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1054(.a(s_72), .O(gate279inter3));
  inv1  gate1055(.a(s_73), .O(gate279inter4));
  nand2 gate1056(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1057(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1058(.a(G651), .O(gate279inter7));
  inv1  gate1059(.a(G803), .O(gate279inter8));
  nand2 gate1060(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1061(.a(s_73), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1062(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1063(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1064(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1457(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1458(.a(gate281inter0), .b(s_130), .O(gate281inter1));
  and2  gate1459(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1460(.a(s_130), .O(gate281inter3));
  inv1  gate1461(.a(s_131), .O(gate281inter4));
  nand2 gate1462(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1463(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1464(.a(G654), .O(gate281inter7));
  inv1  gate1465(.a(G806), .O(gate281inter8));
  nand2 gate1466(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1467(.a(s_131), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1468(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1469(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1470(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1163(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1164(.a(gate292inter0), .b(s_88), .O(gate292inter1));
  and2  gate1165(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1166(.a(s_88), .O(gate292inter3));
  inv1  gate1167(.a(s_89), .O(gate292inter4));
  nand2 gate1168(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1169(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1170(.a(G824), .O(gate292inter7));
  inv1  gate1171(.a(G825), .O(gate292inter8));
  nand2 gate1172(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1173(.a(s_89), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1174(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1175(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1176(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate855(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate856(.a(gate387inter0), .b(s_44), .O(gate387inter1));
  and2  gate857(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate858(.a(s_44), .O(gate387inter3));
  inv1  gate859(.a(s_45), .O(gate387inter4));
  nand2 gate860(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate861(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate862(.a(G1), .O(gate387inter7));
  inv1  gate863(.a(G1036), .O(gate387inter8));
  nand2 gate864(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate865(.a(s_45), .b(gate387inter3), .O(gate387inter10));
  nor2  gate866(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate867(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate868(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1079(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1080(.a(gate390inter0), .b(s_76), .O(gate390inter1));
  and2  gate1081(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1082(.a(s_76), .O(gate390inter3));
  inv1  gate1083(.a(s_77), .O(gate390inter4));
  nand2 gate1084(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1085(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1086(.a(G4), .O(gate390inter7));
  inv1  gate1087(.a(G1045), .O(gate390inter8));
  nand2 gate1088(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1089(.a(s_77), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1090(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1091(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1092(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1401(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1402(.a(gate391inter0), .b(s_122), .O(gate391inter1));
  and2  gate1403(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1404(.a(s_122), .O(gate391inter3));
  inv1  gate1405(.a(s_123), .O(gate391inter4));
  nand2 gate1406(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1407(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1408(.a(G5), .O(gate391inter7));
  inv1  gate1409(.a(G1048), .O(gate391inter8));
  nand2 gate1410(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1411(.a(s_123), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1412(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1413(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1414(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1303(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1304(.a(gate394inter0), .b(s_108), .O(gate394inter1));
  and2  gate1305(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1306(.a(s_108), .O(gate394inter3));
  inv1  gate1307(.a(s_109), .O(gate394inter4));
  nand2 gate1308(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1309(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1310(.a(G8), .O(gate394inter7));
  inv1  gate1311(.a(G1057), .O(gate394inter8));
  nand2 gate1312(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1313(.a(s_109), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1314(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1315(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1316(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate939(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate940(.a(gate415inter0), .b(s_56), .O(gate415inter1));
  and2  gate941(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate942(.a(s_56), .O(gate415inter3));
  inv1  gate943(.a(s_57), .O(gate415inter4));
  nand2 gate944(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate945(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate946(.a(G29), .O(gate415inter7));
  inv1  gate947(.a(G1120), .O(gate415inter8));
  nand2 gate948(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate949(.a(s_57), .b(gate415inter3), .O(gate415inter10));
  nor2  gate950(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate951(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate952(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate771(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate772(.a(gate426inter0), .b(s_32), .O(gate426inter1));
  and2  gate773(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate774(.a(s_32), .O(gate426inter3));
  inv1  gate775(.a(s_33), .O(gate426inter4));
  nand2 gate776(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate777(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate778(.a(G1045), .O(gate426inter7));
  inv1  gate779(.a(G1141), .O(gate426inter8));
  nand2 gate780(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate781(.a(s_33), .b(gate426inter3), .O(gate426inter10));
  nor2  gate782(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate783(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate784(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate953(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate954(.a(gate441inter0), .b(s_58), .O(gate441inter1));
  and2  gate955(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate956(.a(s_58), .O(gate441inter3));
  inv1  gate957(.a(s_59), .O(gate441inter4));
  nand2 gate958(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate959(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate960(.a(G12), .O(gate441inter7));
  inv1  gate961(.a(G1165), .O(gate441inter8));
  nand2 gate962(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate963(.a(s_59), .b(gate441inter3), .O(gate441inter10));
  nor2  gate964(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate965(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate966(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate841(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate842(.a(gate478inter0), .b(s_42), .O(gate478inter1));
  and2  gate843(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate844(.a(s_42), .O(gate478inter3));
  inv1  gate845(.a(s_43), .O(gate478inter4));
  nand2 gate846(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate847(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate848(.a(G1123), .O(gate478inter7));
  inv1  gate849(.a(G1219), .O(gate478inter8));
  nand2 gate850(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate851(.a(s_43), .b(gate478inter3), .O(gate478inter10));
  nor2  gate852(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate853(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate854(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1121(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1122(.a(gate479inter0), .b(s_82), .O(gate479inter1));
  and2  gate1123(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1124(.a(s_82), .O(gate479inter3));
  inv1  gate1125(.a(s_83), .O(gate479inter4));
  nand2 gate1126(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1127(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1128(.a(G31), .O(gate479inter7));
  inv1  gate1129(.a(G1222), .O(gate479inter8));
  nand2 gate1130(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1131(.a(s_83), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1132(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1133(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1134(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate995(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate996(.a(gate483inter0), .b(s_64), .O(gate483inter1));
  and2  gate997(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate998(.a(s_64), .O(gate483inter3));
  inv1  gate999(.a(s_65), .O(gate483inter4));
  nand2 gate1000(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1001(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1002(.a(G1228), .O(gate483inter7));
  inv1  gate1003(.a(G1229), .O(gate483inter8));
  nand2 gate1004(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1005(.a(s_65), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1006(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1007(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1008(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate869(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate870(.a(gate491inter0), .b(s_46), .O(gate491inter1));
  and2  gate871(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate872(.a(s_46), .O(gate491inter3));
  inv1  gate873(.a(s_47), .O(gate491inter4));
  nand2 gate874(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate875(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate876(.a(G1244), .O(gate491inter7));
  inv1  gate877(.a(G1245), .O(gate491inter8));
  nand2 gate878(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate879(.a(s_47), .b(gate491inter3), .O(gate491inter10));
  nor2  gate880(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate881(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate882(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate883(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate884(.a(gate493inter0), .b(s_48), .O(gate493inter1));
  and2  gate885(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate886(.a(s_48), .O(gate493inter3));
  inv1  gate887(.a(s_49), .O(gate493inter4));
  nand2 gate888(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate889(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate890(.a(G1248), .O(gate493inter7));
  inv1  gate891(.a(G1249), .O(gate493inter8));
  nand2 gate892(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate893(.a(s_49), .b(gate493inter3), .O(gate493inter10));
  nor2  gate894(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate895(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate896(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate547(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate548(.a(gate512inter0), .b(s_0), .O(gate512inter1));
  and2  gate549(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate550(.a(s_0), .O(gate512inter3));
  inv1  gate551(.a(s_1), .O(gate512inter4));
  nand2 gate552(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate553(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate554(.a(G1286), .O(gate512inter7));
  inv1  gate555(.a(G1287), .O(gate512inter8));
  nand2 gate556(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate557(.a(s_1), .b(gate512inter3), .O(gate512inter10));
  nor2  gate558(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate559(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate560(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule