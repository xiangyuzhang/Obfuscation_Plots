module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12;

  xor2  gate203(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate204(.a(gate1inter0), .b(s_0), .O(gate1inter1));
  and2  gate205(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate206(.a(s_0), .O(gate1inter3));
  inv1  gate207(.a(s_1), .O(gate1inter4));
  nand2 gate208(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate209(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate210(.a(N1), .O(gate1inter7));
  inv1  gate211(.a(N5), .O(gate1inter8));
  nand2 gate212(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate213(.a(s_1), .b(gate1inter3), .O(gate1inter10));
  nor2  gate214(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate215(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate216(.a(gate1inter12), .b(gate1inter1), .O(N250));

  xor2  gate609(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate610(.a(gate2inter0), .b(s_58), .O(gate2inter1));
  and2  gate611(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate612(.a(s_58), .O(gate2inter3));
  inv1  gate613(.a(s_59), .O(gate2inter4));
  nand2 gate614(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate615(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate616(.a(N9), .O(gate2inter7));
  inv1  gate617(.a(N13), .O(gate2inter8));
  nand2 gate618(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate619(.a(s_59), .b(gate2inter3), .O(gate2inter10));
  nor2  gate620(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate621(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate622(.a(gate2inter12), .b(gate2inter1), .O(N251));
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate553(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate554(.a(gate4inter0), .b(s_50), .O(gate4inter1));
  and2  gate555(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate556(.a(s_50), .O(gate4inter3));
  inv1  gate557(.a(s_51), .O(gate4inter4));
  nand2 gate558(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate559(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate560(.a(N25), .O(gate4inter7));
  inv1  gate561(.a(N29), .O(gate4inter8));
  nand2 gate562(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate563(.a(s_51), .b(gate4inter3), .O(gate4inter10));
  nor2  gate564(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate565(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate566(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate525(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate526(.a(gate8inter0), .b(s_46), .O(gate8inter1));
  and2  gate527(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate528(.a(s_46), .O(gate8inter3));
  inv1  gate529(.a(s_47), .O(gate8inter4));
  nand2 gate530(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate531(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate532(.a(N57), .O(gate8inter7));
  inv1  gate533(.a(N61), .O(gate8inter8));
  nand2 gate534(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate535(.a(s_47), .b(gate8inter3), .O(gate8inter10));
  nor2  gate536(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate537(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate538(.a(gate8inter12), .b(gate8inter1), .O(N257));
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );

  xor2  gate469(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate470(.a(gate11inter0), .b(s_38), .O(gate11inter1));
  and2  gate471(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate472(.a(s_38), .O(gate11inter3));
  inv1  gate473(.a(s_39), .O(gate11inter4));
  nand2 gate474(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate475(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate476(.a(N81), .O(gate11inter7));
  inv1  gate477(.a(N85), .O(gate11inter8));
  nand2 gate478(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate479(.a(s_39), .b(gate11inter3), .O(gate11inter10));
  nor2  gate480(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate481(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate482(.a(gate11inter12), .b(gate11inter1), .O(N260));
xor2 gate12( .a(N89), .b(N93), .O(N261) );

  xor2  gate623(.a(N101), .b(N97), .O(gate13inter0));
  nand2 gate624(.a(gate13inter0), .b(s_60), .O(gate13inter1));
  and2  gate625(.a(N101), .b(N97), .O(gate13inter2));
  inv1  gate626(.a(s_60), .O(gate13inter3));
  inv1  gate627(.a(s_61), .O(gate13inter4));
  nand2 gate628(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate629(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate630(.a(N97), .O(gate13inter7));
  inv1  gate631(.a(N101), .O(gate13inter8));
  nand2 gate632(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate633(.a(s_61), .b(gate13inter3), .O(gate13inter10));
  nor2  gate634(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate635(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate636(.a(gate13inter12), .b(gate13inter1), .O(N262));
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate385(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate386(.a(gate30inter0), .b(s_26), .O(gate30inter1));
  and2  gate387(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate388(.a(s_26), .O(gate30inter3));
  inv1  gate389(.a(s_27), .O(gate30inter4));
  nand2 gate390(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate391(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate392(.a(N41), .O(gate30inter7));
  inv1  gate393(.a(N57), .O(gate30inter8));
  nand2 gate394(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate395(.a(s_27), .b(gate30inter3), .O(gate30inter10));
  nor2  gate396(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate397(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate398(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );

  xor2  gate455(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate456(.a(gate38inter0), .b(s_36), .O(gate38inter1));
  and2  gate457(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate458(.a(s_36), .O(gate38inter3));
  inv1  gate459(.a(s_37), .O(gate38inter4));
  nand2 gate460(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate461(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate462(.a(N105), .O(gate38inter7));
  inv1  gate463(.a(N121), .O(gate38inter8));
  nand2 gate464(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate465(.a(s_37), .b(gate38inter3), .O(gate38inter10));
  nor2  gate466(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate467(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate468(.a(gate38inter12), .b(gate38inter1), .O(N287));

  xor2  gate217(.a(N93), .b(N77), .O(gate39inter0));
  nand2 gate218(.a(gate39inter0), .b(s_2), .O(gate39inter1));
  and2  gate219(.a(N93), .b(N77), .O(gate39inter2));
  inv1  gate220(.a(s_2), .O(gate39inter3));
  inv1  gate221(.a(s_3), .O(gate39inter4));
  nand2 gate222(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate223(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate224(.a(N77), .O(gate39inter7));
  inv1  gate225(.a(N93), .O(gate39inter8));
  nand2 gate226(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate227(.a(s_3), .b(gate39inter3), .O(gate39inter10));
  nor2  gate228(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate229(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate230(.a(gate39inter12), .b(gate39inter1), .O(N288));

  xor2  gate511(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate512(.a(gate40inter0), .b(s_44), .O(gate40inter1));
  and2  gate513(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate514(.a(s_44), .O(gate40inter3));
  inv1  gate515(.a(s_45), .O(gate40inter4));
  nand2 gate516(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate517(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate518(.a(N109), .O(gate40inter7));
  inv1  gate519(.a(N125), .O(gate40inter8));
  nand2 gate520(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate521(.a(s_45), .b(gate40inter3), .O(gate40inter10));
  nor2  gate522(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate523(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate524(.a(gate40inter12), .b(gate40inter1), .O(N289));
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );

  xor2  gate595(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate596(.a(gate43inter0), .b(s_56), .O(gate43inter1));
  and2  gate597(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate598(.a(s_56), .O(gate43inter3));
  inv1  gate599(.a(s_57), .O(gate43inter4));
  nand2 gate600(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate601(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate602(.a(N254), .O(gate43inter7));
  inv1  gate603(.a(N255), .O(gate43inter8));
  nand2 gate604(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate605(.a(s_57), .b(gate43inter3), .O(gate43inter10));
  nor2  gate606(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate607(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate608(.a(gate43inter12), .b(gate43inter1), .O(N296));
xor2 gate44( .a(N256), .b(N257), .O(N299) );

  xor2  gate245(.a(N259), .b(N258), .O(gate45inter0));
  nand2 gate246(.a(gate45inter0), .b(s_6), .O(gate45inter1));
  and2  gate247(.a(N259), .b(N258), .O(gate45inter2));
  inv1  gate248(.a(s_6), .O(gate45inter3));
  inv1  gate249(.a(s_7), .O(gate45inter4));
  nand2 gate250(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate251(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate252(.a(N258), .O(gate45inter7));
  inv1  gate253(.a(N259), .O(gate45inter8));
  nand2 gate254(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate255(.a(s_7), .b(gate45inter3), .O(gate45inter10));
  nor2  gate256(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate257(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate258(.a(gate45inter12), .b(gate45inter1), .O(N302));
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate483(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate484(.a(gate47inter0), .b(s_40), .O(gate47inter1));
  and2  gate485(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate486(.a(s_40), .O(gate47inter3));
  inv1  gate487(.a(s_41), .O(gate47inter4));
  nand2 gate488(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate489(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate490(.a(N262), .O(gate47inter7));
  inv1  gate491(.a(N263), .O(gate47inter8));
  nand2 gate492(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate493(.a(s_41), .b(gate47inter3), .O(gate47inter10));
  nor2  gate494(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate495(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate496(.a(gate47inter12), .b(gate47inter1), .O(N308));
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );

  xor2  gate287(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate288(.a(gate51inter0), .b(s_12), .O(gate51inter1));
  and2  gate289(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate290(.a(s_12), .O(gate51inter3));
  inv1  gate291(.a(s_13), .O(gate51inter4));
  nand2 gate292(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate293(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate294(.a(N278), .O(gate51inter7));
  inv1  gate295(.a(N279), .O(gate51inter8));
  nand2 gate296(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate297(.a(s_13), .b(gate51inter3), .O(gate51inter10));
  nor2  gate298(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate299(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate300(.a(gate51inter12), .b(gate51inter1), .O(N316));
xor2 gate52( .a(N280), .b(N281), .O(N317) );

  xor2  gate539(.a(N283), .b(N282), .O(gate53inter0));
  nand2 gate540(.a(gate53inter0), .b(s_48), .O(gate53inter1));
  and2  gate541(.a(N283), .b(N282), .O(gate53inter2));
  inv1  gate542(.a(s_48), .O(gate53inter3));
  inv1  gate543(.a(s_49), .O(gate53inter4));
  nand2 gate544(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate545(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate546(.a(N282), .O(gate53inter7));
  inv1  gate547(.a(N283), .O(gate53inter8));
  nand2 gate548(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate549(.a(s_49), .b(gate53inter3), .O(gate53inter10));
  nor2  gate550(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate551(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate552(.a(gate53inter12), .b(gate53inter1), .O(N318));
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate301(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate302(.a(gate59inter0), .b(s_14), .O(gate59inter1));
  and2  gate303(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate304(.a(s_14), .O(gate59inter3));
  inv1  gate305(.a(s_15), .O(gate59inter4));
  nand2 gate306(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate307(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate308(.a(N290), .O(gate59inter7));
  inv1  gate309(.a(N296), .O(gate59inter8));
  nand2 gate310(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate311(.a(s_15), .b(gate59inter3), .O(gate59inter10));
  nor2  gate312(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate313(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate314(.a(gate59inter12), .b(gate59inter1), .O(N340));

  xor2  gate497(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate498(.a(gate60inter0), .b(s_42), .O(gate60inter1));
  and2  gate499(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate500(.a(s_42), .O(gate60inter3));
  inv1  gate501(.a(s_43), .O(gate60inter4));
  nand2 gate502(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate503(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate504(.a(N293), .O(gate60inter7));
  inv1  gate505(.a(N299), .O(gate60inter8));
  nand2 gate506(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate507(.a(s_43), .b(gate60inter3), .O(gate60inter10));
  nor2  gate508(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate509(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate510(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate273(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate274(.a(gate62inter0), .b(s_10), .O(gate62inter1));
  and2  gate275(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate276(.a(s_10), .O(gate62inter3));
  inv1  gate277(.a(s_11), .O(gate62inter4));
  nand2 gate278(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate279(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate280(.a(N308), .O(gate62inter7));
  inv1  gate281(.a(N311), .O(gate62inter8));
  nand2 gate282(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate283(.a(s_11), .b(gate62inter3), .O(gate62inter10));
  nor2  gate284(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate285(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate286(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );

  xor2  gate371(.a(N343), .b(N267), .O(gate66inter0));
  nand2 gate372(.a(gate66inter0), .b(s_24), .O(gate66inter1));
  and2  gate373(.a(N343), .b(N267), .O(gate66inter2));
  inv1  gate374(.a(s_24), .O(gate66inter3));
  inv1  gate375(.a(s_25), .O(gate66inter4));
  nand2 gate376(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate377(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate378(.a(N267), .O(gate66inter7));
  inv1  gate379(.a(N343), .O(gate66inter8));
  nand2 gate380(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate381(.a(s_25), .b(gate66inter3), .O(gate66inter10));
  nor2  gate382(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate383(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate384(.a(gate66inter12), .b(gate66inter1), .O(N347));

  xor2  gate357(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate358(.a(gate67inter0), .b(s_22), .O(gate67inter1));
  and2  gate359(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate360(.a(s_22), .O(gate67inter3));
  inv1  gate361(.a(s_23), .O(gate67inter4));
  nand2 gate362(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate363(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate364(.a(N268), .O(gate67inter7));
  inv1  gate365(.a(N344), .O(gate67inter8));
  nand2 gate366(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate367(.a(s_23), .b(gate67inter3), .O(gate67inter10));
  nor2  gate368(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate369(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate370(.a(gate67inter12), .b(gate67inter1), .O(N348));

  xor2  gate259(.a(N345), .b(N269), .O(gate68inter0));
  nand2 gate260(.a(gate68inter0), .b(s_8), .O(gate68inter1));
  and2  gate261(.a(N345), .b(N269), .O(gate68inter2));
  inv1  gate262(.a(s_8), .O(gate68inter3));
  inv1  gate263(.a(s_9), .O(gate68inter4));
  nand2 gate264(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate265(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate266(.a(N269), .O(gate68inter7));
  inv1  gate267(.a(N345), .O(gate68inter8));
  nand2 gate268(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate269(.a(s_9), .b(gate68inter3), .O(gate68inter10));
  nor2  gate270(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate271(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate272(.a(gate68inter12), .b(gate68inter1), .O(N349));
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate329(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate330(.a(gate75inter0), .b(s_18), .O(gate75inter1));
  and2  gate331(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate332(.a(s_18), .O(gate75inter3));
  inv1  gate333(.a(s_19), .O(gate75inter4));
  nand2 gate334(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate335(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate336(.a(N316), .O(gate75inter7));
  inv1  gate337(.a(N348), .O(gate75inter8));
  nand2 gate338(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate339(.a(s_19), .b(gate75inter3), .O(gate75inter10));
  nor2  gate340(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate341(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate342(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate315(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate316(.a(gate172inter0), .b(s_16), .O(gate172inter1));
  and2  gate317(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate318(.a(s_16), .O(gate172inter3));
  inv1  gate319(.a(s_17), .O(gate172inter4));
  nand2 gate320(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate321(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate322(.a(N5), .O(gate172inter7));
  inv1  gate323(.a(N693), .O(gate172inter8));
  nand2 gate324(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate325(.a(s_17), .b(gate172inter3), .O(gate172inter10));
  nor2  gate326(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate327(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate328(.a(gate172inter12), .b(gate172inter1), .O(N725));
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );

  xor2  gate427(.a(N697), .b(N21), .O(gate176inter0));
  nand2 gate428(.a(gate176inter0), .b(s_32), .O(gate176inter1));
  and2  gate429(.a(N697), .b(N21), .O(gate176inter2));
  inv1  gate430(.a(s_32), .O(gate176inter3));
  inv1  gate431(.a(s_33), .O(gate176inter4));
  nand2 gate432(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate433(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate434(.a(N21), .O(gate176inter7));
  inv1  gate435(.a(N697), .O(gate176inter8));
  nand2 gate436(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate437(.a(s_33), .b(gate176inter3), .O(gate176inter10));
  nor2  gate438(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate439(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate440(.a(gate176inter12), .b(gate176inter1), .O(N729));
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );
xor2 gate184( .a(N53), .b(N705), .O(N737) );

  xor2  gate567(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate568(.a(gate185inter0), .b(s_52), .O(gate185inter1));
  and2  gate569(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate570(.a(s_52), .O(gate185inter3));
  inv1  gate571(.a(s_53), .O(gate185inter4));
  nand2 gate572(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate573(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate574(.a(N57), .O(gate185inter7));
  inv1  gate575(.a(N706), .O(gate185inter8));
  nand2 gate576(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate577(.a(s_53), .b(gate185inter3), .O(gate185inter10));
  nor2  gate578(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate579(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate580(.a(gate185inter12), .b(gate185inter1), .O(N738));
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );

  xor2  gate581(.a(N709), .b(N69), .O(gate188inter0));
  nand2 gate582(.a(gate188inter0), .b(s_54), .O(gate188inter1));
  and2  gate583(.a(N709), .b(N69), .O(gate188inter2));
  inv1  gate584(.a(s_54), .O(gate188inter3));
  inv1  gate585(.a(s_55), .O(gate188inter4));
  nand2 gate586(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate587(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate588(.a(N69), .O(gate188inter7));
  inv1  gate589(.a(N709), .O(gate188inter8));
  nand2 gate590(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate591(.a(s_55), .b(gate188inter3), .O(gate188inter10));
  nor2  gate592(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate593(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate594(.a(gate188inter12), .b(gate188inter1), .O(N741));

  xor2  gate399(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate400(.a(gate189inter0), .b(s_28), .O(gate189inter1));
  and2  gate401(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate402(.a(s_28), .O(gate189inter3));
  inv1  gate403(.a(s_29), .O(gate189inter4));
  nand2 gate404(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate405(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate406(.a(N73), .O(gate189inter7));
  inv1  gate407(.a(N710), .O(gate189inter8));
  nand2 gate408(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate409(.a(s_29), .b(gate189inter3), .O(gate189inter10));
  nor2  gate410(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate411(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate412(.a(gate189inter12), .b(gate189inter1), .O(N742));
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );

  xor2  gate343(.a(N714), .b(N89), .O(gate193inter0));
  nand2 gate344(.a(gate193inter0), .b(s_20), .O(gate193inter1));
  and2  gate345(.a(N714), .b(N89), .O(gate193inter2));
  inv1  gate346(.a(s_20), .O(gate193inter3));
  inv1  gate347(.a(s_21), .O(gate193inter4));
  nand2 gate348(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate349(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate350(.a(N89), .O(gate193inter7));
  inv1  gate351(.a(N714), .O(gate193inter8));
  nand2 gate352(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate353(.a(s_21), .b(gate193inter3), .O(gate193inter10));
  nor2  gate354(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate355(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate356(.a(gate193inter12), .b(gate193inter1), .O(N746));

  xor2  gate413(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate414(.a(gate194inter0), .b(s_30), .O(gate194inter1));
  and2  gate415(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate416(.a(s_30), .O(gate194inter3));
  inv1  gate417(.a(s_31), .O(gate194inter4));
  nand2 gate418(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate419(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate420(.a(N93), .O(gate194inter7));
  inv1  gate421(.a(N715), .O(gate194inter8));
  nand2 gate422(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate423(.a(s_31), .b(gate194inter3), .O(gate194inter10));
  nor2  gate424(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate425(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate426(.a(gate194inter12), .b(gate194inter1), .O(N747));

  xor2  gate441(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate442(.a(gate195inter0), .b(s_34), .O(gate195inter1));
  and2  gate443(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate444(.a(s_34), .O(gate195inter3));
  inv1  gate445(.a(s_35), .O(gate195inter4));
  nand2 gate446(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate447(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate448(.a(N97), .O(gate195inter7));
  inv1  gate449(.a(N716), .O(gate195inter8));
  nand2 gate450(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate451(.a(s_35), .b(gate195inter3), .O(gate195inter10));
  nor2  gate452(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate453(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate454(.a(gate195inter12), .b(gate195inter1), .O(N748));

  xor2  gate231(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate232(.a(gate196inter0), .b(s_4), .O(gate196inter1));
  and2  gate233(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate234(.a(s_4), .O(gate196inter3));
  inv1  gate235(.a(s_5), .O(gate196inter4));
  nand2 gate236(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate237(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate238(.a(N101), .O(gate196inter7));
  inv1  gate239(.a(N717), .O(gate196inter8));
  nand2 gate240(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate241(.a(s_5), .b(gate196inter3), .O(gate196inter10));
  nor2  gate242(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate243(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate244(.a(gate196inter12), .b(gate196inter1), .O(N749));
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule