module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate729(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate730(.a(gate19inter0), .b(s_26), .O(gate19inter1));
  and2  gate731(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate732(.a(s_26), .O(gate19inter3));
  inv1  gate733(.a(s_27), .O(gate19inter4));
  nand2 gate734(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate735(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate736(.a(G21), .O(gate19inter7));
  inv1  gate737(.a(G22), .O(gate19inter8));
  nand2 gate738(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate739(.a(s_27), .b(gate19inter3), .O(gate19inter10));
  nor2  gate740(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate741(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate742(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1331(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1332(.a(gate24inter0), .b(s_112), .O(gate24inter1));
  and2  gate1333(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1334(.a(s_112), .O(gate24inter3));
  inv1  gate1335(.a(s_113), .O(gate24inter4));
  nand2 gate1336(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1337(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1338(.a(G31), .O(gate24inter7));
  inv1  gate1339(.a(G32), .O(gate24inter8));
  nand2 gate1340(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1341(.a(s_113), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1342(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1343(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1344(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate673(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate674(.a(gate27inter0), .b(s_18), .O(gate27inter1));
  and2  gate675(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate676(.a(s_18), .O(gate27inter3));
  inv1  gate677(.a(s_19), .O(gate27inter4));
  nand2 gate678(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate679(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate680(.a(G2), .O(gate27inter7));
  inv1  gate681(.a(G6), .O(gate27inter8));
  nand2 gate682(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate683(.a(s_19), .b(gate27inter3), .O(gate27inter10));
  nor2  gate684(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate685(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate686(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1163(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1164(.a(gate31inter0), .b(s_88), .O(gate31inter1));
  and2  gate1165(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1166(.a(s_88), .O(gate31inter3));
  inv1  gate1167(.a(s_89), .O(gate31inter4));
  nand2 gate1168(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1169(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1170(.a(G4), .O(gate31inter7));
  inv1  gate1171(.a(G8), .O(gate31inter8));
  nand2 gate1172(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1173(.a(s_89), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1174(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1175(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1176(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate659(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate660(.a(gate37inter0), .b(s_16), .O(gate37inter1));
  and2  gate661(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate662(.a(s_16), .O(gate37inter3));
  inv1  gate663(.a(s_17), .O(gate37inter4));
  nand2 gate664(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate665(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate666(.a(G19), .O(gate37inter7));
  inv1  gate667(.a(G23), .O(gate37inter8));
  nand2 gate668(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate669(.a(s_17), .b(gate37inter3), .O(gate37inter10));
  nor2  gate670(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate671(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate672(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1387(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1388(.a(gate38inter0), .b(s_120), .O(gate38inter1));
  and2  gate1389(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1390(.a(s_120), .O(gate38inter3));
  inv1  gate1391(.a(s_121), .O(gate38inter4));
  nand2 gate1392(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1393(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1394(.a(G27), .O(gate38inter7));
  inv1  gate1395(.a(G31), .O(gate38inter8));
  nand2 gate1396(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1397(.a(s_121), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1398(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1399(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1400(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate589(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate590(.a(gate51inter0), .b(s_6), .O(gate51inter1));
  and2  gate591(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate592(.a(s_6), .O(gate51inter3));
  inv1  gate593(.a(s_7), .O(gate51inter4));
  nand2 gate594(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate595(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate596(.a(G11), .O(gate51inter7));
  inv1  gate597(.a(G281), .O(gate51inter8));
  nand2 gate598(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate599(.a(s_7), .b(gate51inter3), .O(gate51inter10));
  nor2  gate600(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate601(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate602(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1191(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1192(.a(gate52inter0), .b(s_92), .O(gate52inter1));
  and2  gate1193(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1194(.a(s_92), .O(gate52inter3));
  inv1  gate1195(.a(s_93), .O(gate52inter4));
  nand2 gate1196(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1197(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1198(.a(G12), .O(gate52inter7));
  inv1  gate1199(.a(G281), .O(gate52inter8));
  nand2 gate1200(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1201(.a(s_93), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1202(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1203(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1204(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate715(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate716(.a(gate54inter0), .b(s_24), .O(gate54inter1));
  and2  gate717(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate718(.a(s_24), .O(gate54inter3));
  inv1  gate719(.a(s_25), .O(gate54inter4));
  nand2 gate720(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate721(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate722(.a(G14), .O(gate54inter7));
  inv1  gate723(.a(G284), .O(gate54inter8));
  nand2 gate724(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate725(.a(s_25), .b(gate54inter3), .O(gate54inter10));
  nor2  gate726(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate727(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate728(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate687(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate688(.a(gate55inter0), .b(s_20), .O(gate55inter1));
  and2  gate689(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate690(.a(s_20), .O(gate55inter3));
  inv1  gate691(.a(s_21), .O(gate55inter4));
  nand2 gate692(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate693(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate694(.a(G15), .O(gate55inter7));
  inv1  gate695(.a(G287), .O(gate55inter8));
  nand2 gate696(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate697(.a(s_21), .b(gate55inter3), .O(gate55inter10));
  nor2  gate698(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate699(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate700(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1107(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1108(.a(gate59inter0), .b(s_80), .O(gate59inter1));
  and2  gate1109(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1110(.a(s_80), .O(gate59inter3));
  inv1  gate1111(.a(s_81), .O(gate59inter4));
  nand2 gate1112(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1113(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1114(.a(G19), .O(gate59inter7));
  inv1  gate1115(.a(G293), .O(gate59inter8));
  nand2 gate1116(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1117(.a(s_81), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1118(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1119(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1120(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1541(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1542(.a(gate64inter0), .b(s_142), .O(gate64inter1));
  and2  gate1543(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1544(.a(s_142), .O(gate64inter3));
  inv1  gate1545(.a(s_143), .O(gate64inter4));
  nand2 gate1546(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1547(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1548(.a(G24), .O(gate64inter7));
  inv1  gate1549(.a(G299), .O(gate64inter8));
  nand2 gate1550(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1551(.a(s_143), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1552(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1553(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1554(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1555(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1556(.a(gate67inter0), .b(s_144), .O(gate67inter1));
  and2  gate1557(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1558(.a(s_144), .O(gate67inter3));
  inv1  gate1559(.a(s_145), .O(gate67inter4));
  nand2 gate1560(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1561(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1562(.a(G27), .O(gate67inter7));
  inv1  gate1563(.a(G305), .O(gate67inter8));
  nand2 gate1564(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1565(.a(s_145), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1566(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1567(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1568(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate785(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate786(.a(gate68inter0), .b(s_34), .O(gate68inter1));
  and2  gate787(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate788(.a(s_34), .O(gate68inter3));
  inv1  gate789(.a(s_35), .O(gate68inter4));
  nand2 gate790(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate791(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate792(.a(G28), .O(gate68inter7));
  inv1  gate793(.a(G305), .O(gate68inter8));
  nand2 gate794(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate795(.a(s_35), .b(gate68inter3), .O(gate68inter10));
  nor2  gate796(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate797(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate798(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate813(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate814(.a(gate83inter0), .b(s_38), .O(gate83inter1));
  and2  gate815(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate816(.a(s_38), .O(gate83inter3));
  inv1  gate817(.a(s_39), .O(gate83inter4));
  nand2 gate818(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate819(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate820(.a(G11), .O(gate83inter7));
  inv1  gate821(.a(G329), .O(gate83inter8));
  nand2 gate822(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate823(.a(s_39), .b(gate83inter3), .O(gate83inter10));
  nor2  gate824(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate825(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate826(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate561(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate562(.a(gate85inter0), .b(s_2), .O(gate85inter1));
  and2  gate563(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate564(.a(s_2), .O(gate85inter3));
  inv1  gate565(.a(s_3), .O(gate85inter4));
  nand2 gate566(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate567(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate568(.a(G4), .O(gate85inter7));
  inv1  gate569(.a(G332), .O(gate85inter8));
  nand2 gate570(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate571(.a(s_3), .b(gate85inter3), .O(gate85inter10));
  nor2  gate572(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate573(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate574(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1499(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1500(.a(gate87inter0), .b(s_136), .O(gate87inter1));
  and2  gate1501(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1502(.a(s_136), .O(gate87inter3));
  inv1  gate1503(.a(s_137), .O(gate87inter4));
  nand2 gate1504(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1505(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1506(.a(G12), .O(gate87inter7));
  inv1  gate1507(.a(G335), .O(gate87inter8));
  nand2 gate1508(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1509(.a(s_137), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1510(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1511(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1512(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1051(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1052(.a(gate99inter0), .b(s_72), .O(gate99inter1));
  and2  gate1053(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1054(.a(s_72), .O(gate99inter3));
  inv1  gate1055(.a(s_73), .O(gate99inter4));
  nand2 gate1056(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1057(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1058(.a(G27), .O(gate99inter7));
  inv1  gate1059(.a(G353), .O(gate99inter8));
  nand2 gate1060(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1061(.a(s_73), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1062(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1063(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1064(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate841(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate842(.a(gate103inter0), .b(s_42), .O(gate103inter1));
  and2  gate843(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate844(.a(s_42), .O(gate103inter3));
  inv1  gate845(.a(s_43), .O(gate103inter4));
  nand2 gate846(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate847(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate848(.a(G28), .O(gate103inter7));
  inv1  gate849(.a(G359), .O(gate103inter8));
  nand2 gate850(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate851(.a(s_43), .b(gate103inter3), .O(gate103inter10));
  nor2  gate852(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate853(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate854(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate967(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate968(.a(gate104inter0), .b(s_60), .O(gate104inter1));
  and2  gate969(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate970(.a(s_60), .O(gate104inter3));
  inv1  gate971(.a(s_61), .O(gate104inter4));
  nand2 gate972(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate973(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate974(.a(G32), .O(gate104inter7));
  inv1  gate975(.a(G359), .O(gate104inter8));
  nand2 gate976(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate977(.a(s_61), .b(gate104inter3), .O(gate104inter10));
  nor2  gate978(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate979(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate980(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1023(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1024(.a(gate105inter0), .b(s_68), .O(gate105inter1));
  and2  gate1025(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1026(.a(s_68), .O(gate105inter3));
  inv1  gate1027(.a(s_69), .O(gate105inter4));
  nand2 gate1028(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1029(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1030(.a(G362), .O(gate105inter7));
  inv1  gate1031(.a(G363), .O(gate105inter8));
  nand2 gate1032(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1033(.a(s_69), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1034(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1035(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1036(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1219(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1220(.a(gate108inter0), .b(s_96), .O(gate108inter1));
  and2  gate1221(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1222(.a(s_96), .O(gate108inter3));
  inv1  gate1223(.a(s_97), .O(gate108inter4));
  nand2 gate1224(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1225(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1226(.a(G368), .O(gate108inter7));
  inv1  gate1227(.a(G369), .O(gate108inter8));
  nand2 gate1228(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1229(.a(s_97), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1230(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1231(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1232(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1289(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1290(.a(gate113inter0), .b(s_106), .O(gate113inter1));
  and2  gate1291(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1292(.a(s_106), .O(gate113inter3));
  inv1  gate1293(.a(s_107), .O(gate113inter4));
  nand2 gate1294(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1295(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1296(.a(G378), .O(gate113inter7));
  inv1  gate1297(.a(G379), .O(gate113inter8));
  nand2 gate1298(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1299(.a(s_107), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1300(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1301(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1302(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate925(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate926(.a(gate115inter0), .b(s_54), .O(gate115inter1));
  and2  gate927(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate928(.a(s_54), .O(gate115inter3));
  inv1  gate929(.a(s_55), .O(gate115inter4));
  nand2 gate930(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate931(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate932(.a(G382), .O(gate115inter7));
  inv1  gate933(.a(G383), .O(gate115inter8));
  nand2 gate934(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate935(.a(s_55), .b(gate115inter3), .O(gate115inter10));
  nor2  gate936(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate937(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate938(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1303(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1304(.a(gate119inter0), .b(s_108), .O(gate119inter1));
  and2  gate1305(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1306(.a(s_108), .O(gate119inter3));
  inv1  gate1307(.a(s_109), .O(gate119inter4));
  nand2 gate1308(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1309(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1310(.a(G390), .O(gate119inter7));
  inv1  gate1311(.a(G391), .O(gate119inter8));
  nand2 gate1312(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1313(.a(s_109), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1314(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1315(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1316(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1597(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1598(.a(gate121inter0), .b(s_150), .O(gate121inter1));
  and2  gate1599(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1600(.a(s_150), .O(gate121inter3));
  inv1  gate1601(.a(s_151), .O(gate121inter4));
  nand2 gate1602(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1603(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1604(.a(G394), .O(gate121inter7));
  inv1  gate1605(.a(G395), .O(gate121inter8));
  nand2 gate1606(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1607(.a(s_151), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1608(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1609(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1610(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1373(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1374(.a(gate131inter0), .b(s_118), .O(gate131inter1));
  and2  gate1375(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1376(.a(s_118), .O(gate131inter3));
  inv1  gate1377(.a(s_119), .O(gate131inter4));
  nand2 gate1378(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1379(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1380(.a(G414), .O(gate131inter7));
  inv1  gate1381(.a(G415), .O(gate131inter8));
  nand2 gate1382(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1383(.a(s_119), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1384(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1385(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1386(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1247(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1248(.a(gate137inter0), .b(s_100), .O(gate137inter1));
  and2  gate1249(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1250(.a(s_100), .O(gate137inter3));
  inv1  gate1251(.a(s_101), .O(gate137inter4));
  nand2 gate1252(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1253(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1254(.a(G426), .O(gate137inter7));
  inv1  gate1255(.a(G429), .O(gate137inter8));
  nand2 gate1256(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1257(.a(s_101), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1258(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1259(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1260(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1583(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1584(.a(gate140inter0), .b(s_148), .O(gate140inter1));
  and2  gate1585(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1586(.a(s_148), .O(gate140inter3));
  inv1  gate1587(.a(s_149), .O(gate140inter4));
  nand2 gate1588(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1589(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1590(.a(G444), .O(gate140inter7));
  inv1  gate1591(.a(G447), .O(gate140inter8));
  nand2 gate1592(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1593(.a(s_149), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1594(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1595(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1596(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate799(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate800(.a(gate145inter0), .b(s_36), .O(gate145inter1));
  and2  gate801(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate802(.a(s_36), .O(gate145inter3));
  inv1  gate803(.a(s_37), .O(gate145inter4));
  nand2 gate804(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate805(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate806(.a(G474), .O(gate145inter7));
  inv1  gate807(.a(G477), .O(gate145inter8));
  nand2 gate808(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate809(.a(s_37), .b(gate145inter3), .O(gate145inter10));
  nor2  gate810(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate811(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate812(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1177(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1178(.a(gate157inter0), .b(s_90), .O(gate157inter1));
  and2  gate1179(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1180(.a(s_90), .O(gate157inter3));
  inv1  gate1181(.a(s_91), .O(gate157inter4));
  nand2 gate1182(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1183(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1184(.a(G438), .O(gate157inter7));
  inv1  gate1185(.a(G528), .O(gate157inter8));
  nand2 gate1186(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1187(.a(s_91), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1188(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1189(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1190(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate995(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate996(.a(gate158inter0), .b(s_64), .O(gate158inter1));
  and2  gate997(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate998(.a(s_64), .O(gate158inter3));
  inv1  gate999(.a(s_65), .O(gate158inter4));
  nand2 gate1000(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1001(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1002(.a(G441), .O(gate158inter7));
  inv1  gate1003(.a(G528), .O(gate158inter8));
  nand2 gate1004(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1005(.a(s_65), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1006(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1007(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1008(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1471(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1472(.a(gate165inter0), .b(s_132), .O(gate165inter1));
  and2  gate1473(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1474(.a(s_132), .O(gate165inter3));
  inv1  gate1475(.a(s_133), .O(gate165inter4));
  nand2 gate1476(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1477(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1478(.a(G462), .O(gate165inter7));
  inv1  gate1479(.a(G540), .O(gate165inter8));
  nand2 gate1480(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1481(.a(s_133), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1482(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1483(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1484(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1037(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1038(.a(gate175inter0), .b(s_70), .O(gate175inter1));
  and2  gate1039(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1040(.a(s_70), .O(gate175inter3));
  inv1  gate1041(.a(s_71), .O(gate175inter4));
  nand2 gate1042(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1043(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1044(.a(G492), .O(gate175inter7));
  inv1  gate1045(.a(G555), .O(gate175inter8));
  nand2 gate1046(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1047(.a(s_71), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1048(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1049(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1050(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate827(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate828(.a(gate176inter0), .b(s_40), .O(gate176inter1));
  and2  gate829(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate830(.a(s_40), .O(gate176inter3));
  inv1  gate831(.a(s_41), .O(gate176inter4));
  nand2 gate832(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate833(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate834(.a(G495), .O(gate176inter7));
  inv1  gate835(.a(G555), .O(gate176inter8));
  nand2 gate836(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate837(.a(s_41), .b(gate176inter3), .O(gate176inter10));
  nor2  gate838(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate839(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate840(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate603(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate604(.a(gate180inter0), .b(s_8), .O(gate180inter1));
  and2  gate605(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate606(.a(s_8), .O(gate180inter3));
  inv1  gate607(.a(s_9), .O(gate180inter4));
  nand2 gate608(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate609(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate610(.a(G507), .O(gate180inter7));
  inv1  gate611(.a(G561), .O(gate180inter8));
  nand2 gate612(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate613(.a(s_9), .b(gate180inter3), .O(gate180inter10));
  nor2  gate614(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate615(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate616(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1149(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1150(.a(gate191inter0), .b(s_86), .O(gate191inter1));
  and2  gate1151(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1152(.a(s_86), .O(gate191inter3));
  inv1  gate1153(.a(s_87), .O(gate191inter4));
  nand2 gate1154(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1155(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1156(.a(G582), .O(gate191inter7));
  inv1  gate1157(.a(G583), .O(gate191inter8));
  nand2 gate1158(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1159(.a(s_87), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1160(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1161(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1162(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate575(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate576(.a(gate197inter0), .b(s_4), .O(gate197inter1));
  and2  gate577(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate578(.a(s_4), .O(gate197inter3));
  inv1  gate579(.a(s_5), .O(gate197inter4));
  nand2 gate580(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate581(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate582(.a(G594), .O(gate197inter7));
  inv1  gate583(.a(G595), .O(gate197inter8));
  nand2 gate584(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate585(.a(s_5), .b(gate197inter3), .O(gate197inter10));
  nor2  gate586(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate587(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate588(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate757(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate758(.a(gate199inter0), .b(s_30), .O(gate199inter1));
  and2  gate759(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate760(.a(s_30), .O(gate199inter3));
  inv1  gate761(.a(s_31), .O(gate199inter4));
  nand2 gate762(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate763(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate764(.a(G598), .O(gate199inter7));
  inv1  gate765(.a(G599), .O(gate199inter8));
  nand2 gate766(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate767(.a(s_31), .b(gate199inter3), .O(gate199inter10));
  nor2  gate768(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate769(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate770(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate645(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate646(.a(gate200inter0), .b(s_14), .O(gate200inter1));
  and2  gate647(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate648(.a(s_14), .O(gate200inter3));
  inv1  gate649(.a(s_15), .O(gate200inter4));
  nand2 gate650(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate651(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate652(.a(G600), .O(gate200inter7));
  inv1  gate653(.a(G601), .O(gate200inter8));
  nand2 gate654(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate655(.a(s_15), .b(gate200inter3), .O(gate200inter10));
  nor2  gate656(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate657(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate658(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate883(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate884(.a(gate201inter0), .b(s_48), .O(gate201inter1));
  and2  gate885(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate886(.a(s_48), .O(gate201inter3));
  inv1  gate887(.a(s_49), .O(gate201inter4));
  nand2 gate888(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate889(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate890(.a(G602), .O(gate201inter7));
  inv1  gate891(.a(G607), .O(gate201inter8));
  nand2 gate892(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate893(.a(s_49), .b(gate201inter3), .O(gate201inter10));
  nor2  gate894(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate895(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate896(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate981(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate982(.a(gate224inter0), .b(s_62), .O(gate224inter1));
  and2  gate983(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate984(.a(s_62), .O(gate224inter3));
  inv1  gate985(.a(s_63), .O(gate224inter4));
  nand2 gate986(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate987(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate988(.a(G637), .O(gate224inter7));
  inv1  gate989(.a(G687), .O(gate224inter8));
  nand2 gate990(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate991(.a(s_63), .b(gate224inter3), .O(gate224inter10));
  nor2  gate992(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate993(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate994(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate771(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate772(.a(gate226inter0), .b(s_32), .O(gate226inter1));
  and2  gate773(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate774(.a(s_32), .O(gate226inter3));
  inv1  gate775(.a(s_33), .O(gate226inter4));
  nand2 gate776(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate777(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate778(.a(G692), .O(gate226inter7));
  inv1  gate779(.a(G693), .O(gate226inter8));
  nand2 gate780(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate781(.a(s_33), .b(gate226inter3), .O(gate226inter10));
  nor2  gate782(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate783(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate784(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1415(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1416(.a(gate237inter0), .b(s_124), .O(gate237inter1));
  and2  gate1417(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1418(.a(s_124), .O(gate237inter3));
  inv1  gate1419(.a(s_125), .O(gate237inter4));
  nand2 gate1420(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1421(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1422(.a(G254), .O(gate237inter7));
  inv1  gate1423(.a(G706), .O(gate237inter8));
  nand2 gate1424(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1425(.a(s_125), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1426(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1427(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1428(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate631(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate632(.a(gate238inter0), .b(s_12), .O(gate238inter1));
  and2  gate633(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate634(.a(s_12), .O(gate238inter3));
  inv1  gate635(.a(s_13), .O(gate238inter4));
  nand2 gate636(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate637(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate638(.a(G257), .O(gate238inter7));
  inv1  gate639(.a(G709), .O(gate238inter8));
  nand2 gate640(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate641(.a(s_13), .b(gate238inter3), .O(gate238inter10));
  nor2  gate642(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate643(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate644(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1205(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1206(.a(gate239inter0), .b(s_94), .O(gate239inter1));
  and2  gate1207(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1208(.a(s_94), .O(gate239inter3));
  inv1  gate1209(.a(s_95), .O(gate239inter4));
  nand2 gate1210(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1211(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1212(.a(G260), .O(gate239inter7));
  inv1  gate1213(.a(G712), .O(gate239inter8));
  nand2 gate1214(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1215(.a(s_95), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1216(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1217(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1218(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1233(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1234(.a(gate248inter0), .b(s_98), .O(gate248inter1));
  and2  gate1235(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1236(.a(s_98), .O(gate248inter3));
  inv1  gate1237(.a(s_99), .O(gate248inter4));
  nand2 gate1238(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1239(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1240(.a(G727), .O(gate248inter7));
  inv1  gate1241(.a(G739), .O(gate248inter8));
  nand2 gate1242(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1243(.a(s_99), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1244(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1245(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1246(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate743(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate744(.a(gate249inter0), .b(s_28), .O(gate249inter1));
  and2  gate745(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate746(.a(s_28), .O(gate249inter3));
  inv1  gate747(.a(s_29), .O(gate249inter4));
  nand2 gate748(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate749(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate750(.a(G254), .O(gate249inter7));
  inv1  gate751(.a(G742), .O(gate249inter8));
  nand2 gate752(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate753(.a(s_29), .b(gate249inter3), .O(gate249inter10));
  nor2  gate754(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate755(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate756(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate897(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate898(.a(gate252inter0), .b(s_50), .O(gate252inter1));
  and2  gate899(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate900(.a(s_50), .O(gate252inter3));
  inv1  gate901(.a(s_51), .O(gate252inter4));
  nand2 gate902(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate903(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate904(.a(G709), .O(gate252inter7));
  inv1  gate905(.a(G745), .O(gate252inter8));
  nand2 gate906(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate907(.a(s_51), .b(gate252inter3), .O(gate252inter10));
  nor2  gate908(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate909(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate910(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1065(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1066(.a(gate290inter0), .b(s_74), .O(gate290inter1));
  and2  gate1067(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1068(.a(s_74), .O(gate290inter3));
  inv1  gate1069(.a(s_75), .O(gate290inter4));
  nand2 gate1070(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1071(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1072(.a(G820), .O(gate290inter7));
  inv1  gate1073(.a(G821), .O(gate290inter8));
  nand2 gate1074(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1075(.a(s_75), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1076(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1077(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1078(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate617(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate618(.a(gate296inter0), .b(s_10), .O(gate296inter1));
  and2  gate619(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate620(.a(s_10), .O(gate296inter3));
  inv1  gate621(.a(s_11), .O(gate296inter4));
  nand2 gate622(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate623(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate624(.a(G826), .O(gate296inter7));
  inv1  gate625(.a(G827), .O(gate296inter8));
  nand2 gate626(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate627(.a(s_11), .b(gate296inter3), .O(gate296inter10));
  nor2  gate628(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate629(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate630(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate939(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate940(.a(gate388inter0), .b(s_56), .O(gate388inter1));
  and2  gate941(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate942(.a(s_56), .O(gate388inter3));
  inv1  gate943(.a(s_57), .O(gate388inter4));
  nand2 gate944(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate945(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate946(.a(G2), .O(gate388inter7));
  inv1  gate947(.a(G1039), .O(gate388inter8));
  nand2 gate948(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate949(.a(s_57), .b(gate388inter3), .O(gate388inter10));
  nor2  gate950(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate951(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate952(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1443(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1444(.a(gate407inter0), .b(s_128), .O(gate407inter1));
  and2  gate1445(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1446(.a(s_128), .O(gate407inter3));
  inv1  gate1447(.a(s_129), .O(gate407inter4));
  nand2 gate1448(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1449(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1450(.a(G21), .O(gate407inter7));
  inv1  gate1451(.a(G1096), .O(gate407inter8));
  nand2 gate1452(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1453(.a(s_129), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1454(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1455(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1456(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1093(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1094(.a(gate410inter0), .b(s_78), .O(gate410inter1));
  and2  gate1095(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1096(.a(s_78), .O(gate410inter3));
  inv1  gate1097(.a(s_79), .O(gate410inter4));
  nand2 gate1098(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1099(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1100(.a(G24), .O(gate410inter7));
  inv1  gate1101(.a(G1105), .O(gate410inter8));
  nand2 gate1102(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1103(.a(s_79), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1104(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1105(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1106(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1275(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1276(.a(gate415inter0), .b(s_104), .O(gate415inter1));
  and2  gate1277(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1278(.a(s_104), .O(gate415inter3));
  inv1  gate1279(.a(s_105), .O(gate415inter4));
  nand2 gate1280(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1281(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1282(.a(G29), .O(gate415inter7));
  inv1  gate1283(.a(G1120), .O(gate415inter8));
  nand2 gate1284(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1285(.a(s_105), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1286(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1287(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1288(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1345(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1346(.a(gate422inter0), .b(s_114), .O(gate422inter1));
  and2  gate1347(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1348(.a(s_114), .O(gate422inter3));
  inv1  gate1349(.a(s_115), .O(gate422inter4));
  nand2 gate1350(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1351(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1352(.a(G1039), .O(gate422inter7));
  inv1  gate1353(.a(G1135), .O(gate422inter8));
  nand2 gate1354(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1355(.a(s_115), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1356(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1357(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1358(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate701(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate702(.a(gate427inter0), .b(s_22), .O(gate427inter1));
  and2  gate703(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate704(.a(s_22), .O(gate427inter3));
  inv1  gate705(.a(s_23), .O(gate427inter4));
  nand2 gate706(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate707(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate708(.a(G5), .O(gate427inter7));
  inv1  gate709(.a(G1144), .O(gate427inter8));
  nand2 gate710(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate711(.a(s_23), .b(gate427inter3), .O(gate427inter10));
  nor2  gate712(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate713(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate714(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1009(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1010(.a(gate428inter0), .b(s_66), .O(gate428inter1));
  and2  gate1011(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1012(.a(s_66), .O(gate428inter3));
  inv1  gate1013(.a(s_67), .O(gate428inter4));
  nand2 gate1014(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1015(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1016(.a(G1048), .O(gate428inter7));
  inv1  gate1017(.a(G1144), .O(gate428inter8));
  nand2 gate1018(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1019(.a(s_67), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1020(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1021(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1022(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1485(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1486(.a(gate439inter0), .b(s_134), .O(gate439inter1));
  and2  gate1487(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1488(.a(s_134), .O(gate439inter3));
  inv1  gate1489(.a(s_135), .O(gate439inter4));
  nand2 gate1490(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1491(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1492(.a(G11), .O(gate439inter7));
  inv1  gate1493(.a(G1162), .O(gate439inter8));
  nand2 gate1494(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1495(.a(s_135), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1496(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1497(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1498(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1527(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1528(.a(gate443inter0), .b(s_140), .O(gate443inter1));
  and2  gate1529(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1530(.a(s_140), .O(gate443inter3));
  inv1  gate1531(.a(s_141), .O(gate443inter4));
  nand2 gate1532(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1533(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1534(.a(G13), .O(gate443inter7));
  inv1  gate1535(.a(G1168), .O(gate443inter8));
  nand2 gate1536(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1537(.a(s_141), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1538(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1539(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1540(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1429(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1430(.a(gate451inter0), .b(s_126), .O(gate451inter1));
  and2  gate1431(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1432(.a(s_126), .O(gate451inter3));
  inv1  gate1433(.a(s_127), .O(gate451inter4));
  nand2 gate1434(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1435(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1436(.a(G17), .O(gate451inter7));
  inv1  gate1437(.a(G1180), .O(gate451inter8));
  nand2 gate1438(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1439(.a(s_127), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1440(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1441(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1442(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate869(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate870(.a(gate453inter0), .b(s_46), .O(gate453inter1));
  and2  gate871(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate872(.a(s_46), .O(gate453inter3));
  inv1  gate873(.a(s_47), .O(gate453inter4));
  nand2 gate874(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate875(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate876(.a(G18), .O(gate453inter7));
  inv1  gate877(.a(G1183), .O(gate453inter8));
  nand2 gate878(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate879(.a(s_47), .b(gate453inter3), .O(gate453inter10));
  nor2  gate880(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate881(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate882(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1513(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1514(.a(gate456inter0), .b(s_138), .O(gate456inter1));
  and2  gate1515(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1516(.a(s_138), .O(gate456inter3));
  inv1  gate1517(.a(s_139), .O(gate456inter4));
  nand2 gate1518(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1519(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1520(.a(G1090), .O(gate456inter7));
  inv1  gate1521(.a(G1186), .O(gate456inter8));
  nand2 gate1522(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1523(.a(s_139), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1524(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1525(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1526(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1121(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1122(.a(gate458inter0), .b(s_82), .O(gate458inter1));
  and2  gate1123(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1124(.a(s_82), .O(gate458inter3));
  inv1  gate1125(.a(s_83), .O(gate458inter4));
  nand2 gate1126(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1127(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1128(.a(G1093), .O(gate458inter7));
  inv1  gate1129(.a(G1189), .O(gate458inter8));
  nand2 gate1130(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1131(.a(s_83), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1132(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1133(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1134(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1401(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1402(.a(gate462inter0), .b(s_122), .O(gate462inter1));
  and2  gate1403(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1404(.a(s_122), .O(gate462inter3));
  inv1  gate1405(.a(s_123), .O(gate462inter4));
  nand2 gate1406(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1407(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1408(.a(G1099), .O(gate462inter7));
  inv1  gate1409(.a(G1195), .O(gate462inter8));
  nand2 gate1410(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1411(.a(s_123), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1412(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1413(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1414(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1569(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1570(.a(gate468inter0), .b(s_146), .O(gate468inter1));
  and2  gate1571(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1572(.a(s_146), .O(gate468inter3));
  inv1  gate1573(.a(s_147), .O(gate468inter4));
  nand2 gate1574(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1575(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1576(.a(G1108), .O(gate468inter7));
  inv1  gate1577(.a(G1204), .O(gate468inter8));
  nand2 gate1578(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1579(.a(s_147), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1580(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1581(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1582(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate911(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate912(.a(gate471inter0), .b(s_52), .O(gate471inter1));
  and2  gate913(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate914(.a(s_52), .O(gate471inter3));
  inv1  gate915(.a(s_53), .O(gate471inter4));
  nand2 gate916(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate917(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate918(.a(G27), .O(gate471inter7));
  inv1  gate919(.a(G1210), .O(gate471inter8));
  nand2 gate920(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate921(.a(s_53), .b(gate471inter3), .O(gate471inter10));
  nor2  gate922(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate923(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate924(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1079(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1080(.a(gate476inter0), .b(s_76), .O(gate476inter1));
  and2  gate1081(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1082(.a(s_76), .O(gate476inter3));
  inv1  gate1083(.a(s_77), .O(gate476inter4));
  nand2 gate1084(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1085(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1086(.a(G1120), .O(gate476inter7));
  inv1  gate1087(.a(G1216), .O(gate476inter8));
  nand2 gate1088(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1089(.a(s_77), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1090(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1091(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1092(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate547(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate548(.a(gate479inter0), .b(s_0), .O(gate479inter1));
  and2  gate549(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate550(.a(s_0), .O(gate479inter3));
  inv1  gate551(.a(s_1), .O(gate479inter4));
  nand2 gate552(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate553(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate554(.a(G31), .O(gate479inter7));
  inv1  gate555(.a(G1222), .O(gate479inter8));
  nand2 gate556(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate557(.a(s_1), .b(gate479inter3), .O(gate479inter10));
  nor2  gate558(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate559(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate560(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1317(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1318(.a(gate486inter0), .b(s_110), .O(gate486inter1));
  and2  gate1319(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1320(.a(s_110), .O(gate486inter3));
  inv1  gate1321(.a(s_111), .O(gate486inter4));
  nand2 gate1322(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1323(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1324(.a(G1234), .O(gate486inter7));
  inv1  gate1325(.a(G1235), .O(gate486inter8));
  nand2 gate1326(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1327(.a(s_111), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1328(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1329(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1330(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate855(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate856(.a(gate500inter0), .b(s_44), .O(gate500inter1));
  and2  gate857(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate858(.a(s_44), .O(gate500inter3));
  inv1  gate859(.a(s_45), .O(gate500inter4));
  nand2 gate860(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate861(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate862(.a(G1262), .O(gate500inter7));
  inv1  gate863(.a(G1263), .O(gate500inter8));
  nand2 gate864(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate865(.a(s_45), .b(gate500inter3), .O(gate500inter10));
  nor2  gate866(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate867(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate868(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1261(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1262(.a(gate501inter0), .b(s_102), .O(gate501inter1));
  and2  gate1263(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1264(.a(s_102), .O(gate501inter3));
  inv1  gate1265(.a(s_103), .O(gate501inter4));
  nand2 gate1266(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1267(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1268(.a(G1264), .O(gate501inter7));
  inv1  gate1269(.a(G1265), .O(gate501inter8));
  nand2 gate1270(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1271(.a(s_103), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1272(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1273(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1274(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate953(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate954(.a(gate502inter0), .b(s_58), .O(gate502inter1));
  and2  gate955(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate956(.a(s_58), .O(gate502inter3));
  inv1  gate957(.a(s_59), .O(gate502inter4));
  nand2 gate958(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate959(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate960(.a(G1266), .O(gate502inter7));
  inv1  gate961(.a(G1267), .O(gate502inter8));
  nand2 gate962(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate963(.a(s_59), .b(gate502inter3), .O(gate502inter10));
  nor2  gate964(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate965(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate966(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1359(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1360(.a(gate506inter0), .b(s_116), .O(gate506inter1));
  and2  gate1361(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1362(.a(s_116), .O(gate506inter3));
  inv1  gate1363(.a(s_117), .O(gate506inter4));
  nand2 gate1364(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1365(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1366(.a(G1274), .O(gate506inter7));
  inv1  gate1367(.a(G1275), .O(gate506inter8));
  nand2 gate1368(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1369(.a(s_117), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1370(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1371(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1372(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1457(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1458(.a(gate511inter0), .b(s_130), .O(gate511inter1));
  and2  gate1459(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1460(.a(s_130), .O(gate511inter3));
  inv1  gate1461(.a(s_131), .O(gate511inter4));
  nand2 gate1462(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1463(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1464(.a(G1284), .O(gate511inter7));
  inv1  gate1465(.a(G1285), .O(gate511inter8));
  nand2 gate1466(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1467(.a(s_131), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1468(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1469(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1470(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1135(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1136(.a(gate513inter0), .b(s_84), .O(gate513inter1));
  and2  gate1137(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1138(.a(s_84), .O(gate513inter3));
  inv1  gate1139(.a(s_85), .O(gate513inter4));
  nand2 gate1140(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1141(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1142(.a(G1288), .O(gate513inter7));
  inv1  gate1143(.a(G1289), .O(gate513inter8));
  nand2 gate1144(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1145(.a(s_85), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1146(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1147(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1148(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule