module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate701(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate702(.a(gate15inter0), .b(s_22), .O(gate15inter1));
  and2  gate703(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate704(.a(s_22), .O(gate15inter3));
  inv1  gate705(.a(s_23), .O(gate15inter4));
  nand2 gate706(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate707(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate708(.a(G13), .O(gate15inter7));
  inv1  gate709(.a(G14), .O(gate15inter8));
  nand2 gate710(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate711(.a(s_23), .b(gate15inter3), .O(gate15inter10));
  nor2  gate712(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate713(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate714(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1079(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1080(.a(gate28inter0), .b(s_76), .O(gate28inter1));
  and2  gate1081(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1082(.a(s_76), .O(gate28inter3));
  inv1  gate1083(.a(s_77), .O(gate28inter4));
  nand2 gate1084(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1085(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1086(.a(G10), .O(gate28inter7));
  inv1  gate1087(.a(G14), .O(gate28inter8));
  nand2 gate1088(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1089(.a(s_77), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1090(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1091(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1092(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1023(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1024(.a(gate31inter0), .b(s_68), .O(gate31inter1));
  and2  gate1025(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1026(.a(s_68), .O(gate31inter3));
  inv1  gate1027(.a(s_69), .O(gate31inter4));
  nand2 gate1028(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1029(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1030(.a(G4), .O(gate31inter7));
  inv1  gate1031(.a(G8), .O(gate31inter8));
  nand2 gate1032(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1033(.a(s_69), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1034(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1035(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1036(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate981(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate982(.a(gate38inter0), .b(s_62), .O(gate38inter1));
  and2  gate983(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate984(.a(s_62), .O(gate38inter3));
  inv1  gate985(.a(s_63), .O(gate38inter4));
  nand2 gate986(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate987(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate988(.a(G27), .O(gate38inter7));
  inv1  gate989(.a(G31), .O(gate38inter8));
  nand2 gate990(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate991(.a(s_63), .b(gate38inter3), .O(gate38inter10));
  nor2  gate992(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate993(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate994(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1205(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1206(.a(gate42inter0), .b(s_94), .O(gate42inter1));
  and2  gate1207(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1208(.a(s_94), .O(gate42inter3));
  inv1  gate1209(.a(s_95), .O(gate42inter4));
  nand2 gate1210(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1211(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1212(.a(G2), .O(gate42inter7));
  inv1  gate1213(.a(G266), .O(gate42inter8));
  nand2 gate1214(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1215(.a(s_95), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1216(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1217(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1218(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate575(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate576(.a(gate49inter0), .b(s_4), .O(gate49inter1));
  and2  gate577(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate578(.a(s_4), .O(gate49inter3));
  inv1  gate579(.a(s_5), .O(gate49inter4));
  nand2 gate580(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate581(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate582(.a(G9), .O(gate49inter7));
  inv1  gate583(.a(G278), .O(gate49inter8));
  nand2 gate584(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate585(.a(s_5), .b(gate49inter3), .O(gate49inter10));
  nor2  gate586(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate587(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate588(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate547(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate548(.a(gate51inter0), .b(s_0), .O(gate51inter1));
  and2  gate549(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate550(.a(s_0), .O(gate51inter3));
  inv1  gate551(.a(s_1), .O(gate51inter4));
  nand2 gate552(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate553(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate554(.a(G11), .O(gate51inter7));
  inv1  gate555(.a(G281), .O(gate51inter8));
  nand2 gate556(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate557(.a(s_1), .b(gate51inter3), .O(gate51inter10));
  nor2  gate558(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate559(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate560(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1009(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1010(.a(gate61inter0), .b(s_66), .O(gate61inter1));
  and2  gate1011(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1012(.a(s_66), .O(gate61inter3));
  inv1  gate1013(.a(s_67), .O(gate61inter4));
  nand2 gate1014(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1015(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1016(.a(G21), .O(gate61inter7));
  inv1  gate1017(.a(G296), .O(gate61inter8));
  nand2 gate1018(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1019(.a(s_67), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1020(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1021(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1022(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate939(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate940(.a(gate62inter0), .b(s_56), .O(gate62inter1));
  and2  gate941(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate942(.a(s_56), .O(gate62inter3));
  inv1  gate943(.a(s_57), .O(gate62inter4));
  nand2 gate944(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate945(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate946(.a(G22), .O(gate62inter7));
  inv1  gate947(.a(G296), .O(gate62inter8));
  nand2 gate948(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate949(.a(s_57), .b(gate62inter3), .O(gate62inter10));
  nor2  gate950(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate951(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate952(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1135(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1136(.a(gate64inter0), .b(s_84), .O(gate64inter1));
  and2  gate1137(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1138(.a(s_84), .O(gate64inter3));
  inv1  gate1139(.a(s_85), .O(gate64inter4));
  nand2 gate1140(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1141(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1142(.a(G24), .O(gate64inter7));
  inv1  gate1143(.a(G299), .O(gate64inter8));
  nand2 gate1144(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1145(.a(s_85), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1146(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1147(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1148(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate911(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate912(.a(gate66inter0), .b(s_52), .O(gate66inter1));
  and2  gate913(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate914(.a(s_52), .O(gate66inter3));
  inv1  gate915(.a(s_53), .O(gate66inter4));
  nand2 gate916(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate917(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate918(.a(G26), .O(gate66inter7));
  inv1  gate919(.a(G302), .O(gate66inter8));
  nand2 gate920(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate921(.a(s_53), .b(gate66inter3), .O(gate66inter10));
  nor2  gate922(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate923(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate924(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate883(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate884(.a(gate74inter0), .b(s_48), .O(gate74inter1));
  and2  gate885(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate886(.a(s_48), .O(gate74inter3));
  inv1  gate887(.a(s_49), .O(gate74inter4));
  nand2 gate888(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate889(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate890(.a(G5), .O(gate74inter7));
  inv1  gate891(.a(G314), .O(gate74inter8));
  nand2 gate892(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate893(.a(s_49), .b(gate74inter3), .O(gate74inter10));
  nor2  gate894(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate895(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate896(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate715(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate716(.a(gate80inter0), .b(s_24), .O(gate80inter1));
  and2  gate717(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate718(.a(s_24), .O(gate80inter3));
  inv1  gate719(.a(s_25), .O(gate80inter4));
  nand2 gate720(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate721(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate722(.a(G14), .O(gate80inter7));
  inv1  gate723(.a(G323), .O(gate80inter8));
  nand2 gate724(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate725(.a(s_25), .b(gate80inter3), .O(gate80inter10));
  nor2  gate726(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate727(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate728(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate603(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate604(.a(gate87inter0), .b(s_8), .O(gate87inter1));
  and2  gate605(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate606(.a(s_8), .O(gate87inter3));
  inv1  gate607(.a(s_9), .O(gate87inter4));
  nand2 gate608(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate609(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate610(.a(G12), .O(gate87inter7));
  inv1  gate611(.a(G335), .O(gate87inter8));
  nand2 gate612(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate613(.a(s_9), .b(gate87inter3), .O(gate87inter10));
  nor2  gate614(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate615(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate616(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate897(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate898(.a(gate104inter0), .b(s_50), .O(gate104inter1));
  and2  gate899(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate900(.a(s_50), .O(gate104inter3));
  inv1  gate901(.a(s_51), .O(gate104inter4));
  nand2 gate902(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate903(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate904(.a(G32), .O(gate104inter7));
  inv1  gate905(.a(G359), .O(gate104inter8));
  nand2 gate906(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate907(.a(s_51), .b(gate104inter3), .O(gate104inter10));
  nor2  gate908(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate909(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate910(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate743(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate744(.a(gate110inter0), .b(s_28), .O(gate110inter1));
  and2  gate745(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate746(.a(s_28), .O(gate110inter3));
  inv1  gate747(.a(s_29), .O(gate110inter4));
  nand2 gate748(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate749(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate750(.a(G372), .O(gate110inter7));
  inv1  gate751(.a(G373), .O(gate110inter8));
  nand2 gate752(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate753(.a(s_29), .b(gate110inter3), .O(gate110inter10));
  nor2  gate754(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate755(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate756(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate995(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate996(.a(gate113inter0), .b(s_64), .O(gate113inter1));
  and2  gate997(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate998(.a(s_64), .O(gate113inter3));
  inv1  gate999(.a(s_65), .O(gate113inter4));
  nand2 gate1000(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1001(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1002(.a(G378), .O(gate113inter7));
  inv1  gate1003(.a(G379), .O(gate113inter8));
  nand2 gate1004(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1005(.a(s_65), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1006(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1007(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1008(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate757(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate758(.a(gate118inter0), .b(s_30), .O(gate118inter1));
  and2  gate759(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate760(.a(s_30), .O(gate118inter3));
  inv1  gate761(.a(s_31), .O(gate118inter4));
  nand2 gate762(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate763(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate764(.a(G388), .O(gate118inter7));
  inv1  gate765(.a(G389), .O(gate118inter8));
  nand2 gate766(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate767(.a(s_31), .b(gate118inter3), .O(gate118inter10));
  nor2  gate768(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate769(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate770(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1037(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1038(.a(gate123inter0), .b(s_70), .O(gate123inter1));
  and2  gate1039(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1040(.a(s_70), .O(gate123inter3));
  inv1  gate1041(.a(s_71), .O(gate123inter4));
  nand2 gate1042(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1043(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1044(.a(G398), .O(gate123inter7));
  inv1  gate1045(.a(G399), .O(gate123inter8));
  nand2 gate1046(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1047(.a(s_71), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1048(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1049(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1050(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1163(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1164(.a(gate137inter0), .b(s_88), .O(gate137inter1));
  and2  gate1165(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1166(.a(s_88), .O(gate137inter3));
  inv1  gate1167(.a(s_89), .O(gate137inter4));
  nand2 gate1168(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1169(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1170(.a(G426), .O(gate137inter7));
  inv1  gate1171(.a(G429), .O(gate137inter8));
  nand2 gate1172(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1173(.a(s_89), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1174(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1175(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1176(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate631(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate632(.a(gate143inter0), .b(s_12), .O(gate143inter1));
  and2  gate633(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate634(.a(s_12), .O(gate143inter3));
  inv1  gate635(.a(s_13), .O(gate143inter4));
  nand2 gate636(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate637(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate638(.a(G462), .O(gate143inter7));
  inv1  gate639(.a(G465), .O(gate143inter8));
  nand2 gate640(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate641(.a(s_13), .b(gate143inter3), .O(gate143inter10));
  nor2  gate642(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate643(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate644(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate813(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate814(.a(gate152inter0), .b(s_38), .O(gate152inter1));
  and2  gate815(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate816(.a(s_38), .O(gate152inter3));
  inv1  gate817(.a(s_39), .O(gate152inter4));
  nand2 gate818(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate819(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate820(.a(G516), .O(gate152inter7));
  inv1  gate821(.a(G519), .O(gate152inter8));
  nand2 gate822(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate823(.a(s_39), .b(gate152inter3), .O(gate152inter10));
  nor2  gate824(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate825(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate826(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1093(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1094(.a(gate155inter0), .b(s_78), .O(gate155inter1));
  and2  gate1095(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1096(.a(s_78), .O(gate155inter3));
  inv1  gate1097(.a(s_79), .O(gate155inter4));
  nand2 gate1098(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1099(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1100(.a(G432), .O(gate155inter7));
  inv1  gate1101(.a(G525), .O(gate155inter8));
  nand2 gate1102(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1103(.a(s_79), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1104(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1105(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1106(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1247(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1248(.a(gate158inter0), .b(s_100), .O(gate158inter1));
  and2  gate1249(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1250(.a(s_100), .O(gate158inter3));
  inv1  gate1251(.a(s_101), .O(gate158inter4));
  nand2 gate1252(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1253(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1254(.a(G441), .O(gate158inter7));
  inv1  gate1255(.a(G528), .O(gate158inter8));
  nand2 gate1256(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1257(.a(s_101), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1258(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1259(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1260(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate785(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate786(.a(gate160inter0), .b(s_34), .O(gate160inter1));
  and2  gate787(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate788(.a(s_34), .O(gate160inter3));
  inv1  gate789(.a(s_35), .O(gate160inter4));
  nand2 gate790(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate791(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate792(.a(G447), .O(gate160inter7));
  inv1  gate793(.a(G531), .O(gate160inter8));
  nand2 gate794(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate795(.a(s_35), .b(gate160inter3), .O(gate160inter10));
  nor2  gate796(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate797(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate798(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate589(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate590(.a(gate188inter0), .b(s_6), .O(gate188inter1));
  and2  gate591(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate592(.a(s_6), .O(gate188inter3));
  inv1  gate593(.a(s_7), .O(gate188inter4));
  nand2 gate594(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate595(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate596(.a(G576), .O(gate188inter7));
  inv1  gate597(.a(G577), .O(gate188inter8));
  nand2 gate598(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate599(.a(s_7), .b(gate188inter3), .O(gate188inter10));
  nor2  gate600(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate601(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate602(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1065(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1066(.a(gate192inter0), .b(s_74), .O(gate192inter1));
  and2  gate1067(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1068(.a(s_74), .O(gate192inter3));
  inv1  gate1069(.a(s_75), .O(gate192inter4));
  nand2 gate1070(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1071(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1072(.a(G584), .O(gate192inter7));
  inv1  gate1073(.a(G585), .O(gate192inter8));
  nand2 gate1074(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1075(.a(s_75), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1076(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1077(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1078(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate799(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate800(.a(gate202inter0), .b(s_36), .O(gate202inter1));
  and2  gate801(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate802(.a(s_36), .O(gate202inter3));
  inv1  gate803(.a(s_37), .O(gate202inter4));
  nand2 gate804(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate805(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate806(.a(G612), .O(gate202inter7));
  inv1  gate807(.a(G617), .O(gate202inter8));
  nand2 gate808(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate809(.a(s_37), .b(gate202inter3), .O(gate202inter10));
  nor2  gate810(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate811(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate812(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1121(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1122(.a(gate203inter0), .b(s_82), .O(gate203inter1));
  and2  gate1123(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1124(.a(s_82), .O(gate203inter3));
  inv1  gate1125(.a(s_83), .O(gate203inter4));
  nand2 gate1126(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1127(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1128(.a(G602), .O(gate203inter7));
  inv1  gate1129(.a(G612), .O(gate203inter8));
  nand2 gate1130(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1131(.a(s_83), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1132(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1133(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1134(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1107(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1108(.a(gate219inter0), .b(s_80), .O(gate219inter1));
  and2  gate1109(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1110(.a(s_80), .O(gate219inter3));
  inv1  gate1111(.a(s_81), .O(gate219inter4));
  nand2 gate1112(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1113(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1114(.a(G632), .O(gate219inter7));
  inv1  gate1115(.a(G681), .O(gate219inter8));
  nand2 gate1116(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1117(.a(s_81), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1118(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1119(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1120(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate561(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate562(.a(gate228inter0), .b(s_2), .O(gate228inter1));
  and2  gate563(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate564(.a(s_2), .O(gate228inter3));
  inv1  gate565(.a(s_3), .O(gate228inter4));
  nand2 gate566(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate567(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate568(.a(G696), .O(gate228inter7));
  inv1  gate569(.a(G697), .O(gate228inter8));
  nand2 gate570(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate571(.a(s_3), .b(gate228inter3), .O(gate228inter10));
  nor2  gate572(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate573(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate574(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate869(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate870(.a(gate237inter0), .b(s_46), .O(gate237inter1));
  and2  gate871(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate872(.a(s_46), .O(gate237inter3));
  inv1  gate873(.a(s_47), .O(gate237inter4));
  nand2 gate874(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate875(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate876(.a(G254), .O(gate237inter7));
  inv1  gate877(.a(G706), .O(gate237inter8));
  nand2 gate878(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate879(.a(s_47), .b(gate237inter3), .O(gate237inter10));
  nor2  gate880(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate881(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate882(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1149(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1150(.a(gate240inter0), .b(s_86), .O(gate240inter1));
  and2  gate1151(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1152(.a(s_86), .O(gate240inter3));
  inv1  gate1153(.a(s_87), .O(gate240inter4));
  nand2 gate1154(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1155(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1156(.a(G263), .O(gate240inter7));
  inv1  gate1157(.a(G715), .O(gate240inter8));
  nand2 gate1158(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1159(.a(s_87), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1160(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1161(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1162(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate967(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate968(.a(gate266inter0), .b(s_60), .O(gate266inter1));
  and2  gate969(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate970(.a(s_60), .O(gate266inter3));
  inv1  gate971(.a(s_61), .O(gate266inter4));
  nand2 gate972(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate973(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate974(.a(G645), .O(gate266inter7));
  inv1  gate975(.a(G773), .O(gate266inter8));
  nand2 gate976(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate977(.a(s_61), .b(gate266inter3), .O(gate266inter10));
  nor2  gate978(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate979(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate980(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1233(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1234(.a(gate280inter0), .b(s_98), .O(gate280inter1));
  and2  gate1235(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1236(.a(s_98), .O(gate280inter3));
  inv1  gate1237(.a(s_99), .O(gate280inter4));
  nand2 gate1238(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1239(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1240(.a(G779), .O(gate280inter7));
  inv1  gate1241(.a(G803), .O(gate280inter8));
  nand2 gate1242(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1243(.a(s_99), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1244(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1245(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1246(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1051(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1052(.a(gate281inter0), .b(s_72), .O(gate281inter1));
  and2  gate1053(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1054(.a(s_72), .O(gate281inter3));
  inv1  gate1055(.a(s_73), .O(gate281inter4));
  nand2 gate1056(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1057(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1058(.a(G654), .O(gate281inter7));
  inv1  gate1059(.a(G806), .O(gate281inter8));
  nand2 gate1060(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1061(.a(s_73), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1062(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1063(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1064(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate855(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate856(.a(gate282inter0), .b(s_44), .O(gate282inter1));
  and2  gate857(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate858(.a(s_44), .O(gate282inter3));
  inv1  gate859(.a(s_45), .O(gate282inter4));
  nand2 gate860(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate861(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate862(.a(G782), .O(gate282inter7));
  inv1  gate863(.a(G806), .O(gate282inter8));
  nand2 gate864(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate865(.a(s_45), .b(gate282inter3), .O(gate282inter10));
  nor2  gate866(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate867(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate868(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate673(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate674(.a(gate287inter0), .b(s_18), .O(gate287inter1));
  and2  gate675(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate676(.a(s_18), .O(gate287inter3));
  inv1  gate677(.a(s_19), .O(gate287inter4));
  nand2 gate678(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate679(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate680(.a(G663), .O(gate287inter7));
  inv1  gate681(.a(G815), .O(gate287inter8));
  nand2 gate682(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate683(.a(s_19), .b(gate287inter3), .O(gate287inter10));
  nor2  gate684(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate685(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate686(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate617(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate618(.a(gate390inter0), .b(s_10), .O(gate390inter1));
  and2  gate619(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate620(.a(s_10), .O(gate390inter3));
  inv1  gate621(.a(s_11), .O(gate390inter4));
  nand2 gate622(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate623(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate624(.a(G4), .O(gate390inter7));
  inv1  gate625(.a(G1045), .O(gate390inter8));
  nand2 gate626(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate627(.a(s_11), .b(gate390inter3), .O(gate390inter10));
  nor2  gate628(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate629(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate630(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate771(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate772(.a(gate401inter0), .b(s_32), .O(gate401inter1));
  and2  gate773(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate774(.a(s_32), .O(gate401inter3));
  inv1  gate775(.a(s_33), .O(gate401inter4));
  nand2 gate776(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate777(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate778(.a(G15), .O(gate401inter7));
  inv1  gate779(.a(G1078), .O(gate401inter8));
  nand2 gate780(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate781(.a(s_33), .b(gate401inter3), .O(gate401inter10));
  nor2  gate782(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate783(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate784(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate659(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate660(.a(gate405inter0), .b(s_16), .O(gate405inter1));
  and2  gate661(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate662(.a(s_16), .O(gate405inter3));
  inv1  gate663(.a(s_17), .O(gate405inter4));
  nand2 gate664(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate665(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate666(.a(G19), .O(gate405inter7));
  inv1  gate667(.a(G1090), .O(gate405inter8));
  nand2 gate668(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate669(.a(s_17), .b(gate405inter3), .O(gate405inter10));
  nor2  gate670(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate671(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate672(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate827(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate828(.a(gate418inter0), .b(s_40), .O(gate418inter1));
  and2  gate829(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate830(.a(s_40), .O(gate418inter3));
  inv1  gate831(.a(s_41), .O(gate418inter4));
  nand2 gate832(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate833(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate834(.a(G32), .O(gate418inter7));
  inv1  gate835(.a(G1129), .O(gate418inter8));
  nand2 gate836(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate837(.a(s_41), .b(gate418inter3), .O(gate418inter10));
  nor2  gate838(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate839(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate840(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate841(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate842(.a(gate421inter0), .b(s_42), .O(gate421inter1));
  and2  gate843(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate844(.a(s_42), .O(gate421inter3));
  inv1  gate845(.a(s_43), .O(gate421inter4));
  nand2 gate846(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate847(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate848(.a(G2), .O(gate421inter7));
  inv1  gate849(.a(G1135), .O(gate421inter8));
  nand2 gate850(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate851(.a(s_43), .b(gate421inter3), .O(gate421inter10));
  nor2  gate852(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate853(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate854(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1191(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1192(.a(gate425inter0), .b(s_92), .O(gate425inter1));
  and2  gate1193(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1194(.a(s_92), .O(gate425inter3));
  inv1  gate1195(.a(s_93), .O(gate425inter4));
  nand2 gate1196(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1197(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1198(.a(G4), .O(gate425inter7));
  inv1  gate1199(.a(G1141), .O(gate425inter8));
  nand2 gate1200(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1201(.a(s_93), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1202(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1203(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1204(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate645(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate646(.a(gate429inter0), .b(s_14), .O(gate429inter1));
  and2  gate647(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate648(.a(s_14), .O(gate429inter3));
  inv1  gate649(.a(s_15), .O(gate429inter4));
  nand2 gate650(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate651(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate652(.a(G6), .O(gate429inter7));
  inv1  gate653(.a(G1147), .O(gate429inter8));
  nand2 gate654(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate655(.a(s_15), .b(gate429inter3), .O(gate429inter10));
  nor2  gate656(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate657(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate658(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate729(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate730(.a(gate445inter0), .b(s_26), .O(gate445inter1));
  and2  gate731(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate732(.a(s_26), .O(gate445inter3));
  inv1  gate733(.a(s_27), .O(gate445inter4));
  nand2 gate734(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate735(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate736(.a(G14), .O(gate445inter7));
  inv1  gate737(.a(G1171), .O(gate445inter8));
  nand2 gate738(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate739(.a(s_27), .b(gate445inter3), .O(gate445inter10));
  nor2  gate740(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate741(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate742(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate925(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate926(.a(gate453inter0), .b(s_54), .O(gate453inter1));
  and2  gate927(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate928(.a(s_54), .O(gate453inter3));
  inv1  gate929(.a(s_55), .O(gate453inter4));
  nand2 gate930(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate931(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate932(.a(G18), .O(gate453inter7));
  inv1  gate933(.a(G1183), .O(gate453inter8));
  nand2 gate934(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate935(.a(s_55), .b(gate453inter3), .O(gate453inter10));
  nor2  gate936(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate937(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate938(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate687(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate688(.a(gate466inter0), .b(s_20), .O(gate466inter1));
  and2  gate689(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate690(.a(s_20), .O(gate466inter3));
  inv1  gate691(.a(s_21), .O(gate466inter4));
  nand2 gate692(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate693(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate694(.a(G1105), .O(gate466inter7));
  inv1  gate695(.a(G1201), .O(gate466inter8));
  nand2 gate696(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate697(.a(s_21), .b(gate466inter3), .O(gate466inter10));
  nor2  gate698(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate699(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate700(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate953(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate954(.a(gate478inter0), .b(s_58), .O(gate478inter1));
  and2  gate955(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate956(.a(s_58), .O(gate478inter3));
  inv1  gate957(.a(s_59), .O(gate478inter4));
  nand2 gate958(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate959(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate960(.a(G1123), .O(gate478inter7));
  inv1  gate961(.a(G1219), .O(gate478inter8));
  nand2 gate962(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate963(.a(s_59), .b(gate478inter3), .O(gate478inter10));
  nor2  gate964(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate965(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate966(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1177(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1178(.a(gate493inter0), .b(s_90), .O(gate493inter1));
  and2  gate1179(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1180(.a(s_90), .O(gate493inter3));
  inv1  gate1181(.a(s_91), .O(gate493inter4));
  nand2 gate1182(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1183(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1184(.a(G1248), .O(gate493inter7));
  inv1  gate1185(.a(G1249), .O(gate493inter8));
  nand2 gate1186(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1187(.a(s_91), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1188(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1189(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1190(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1219(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1220(.a(gate495inter0), .b(s_96), .O(gate495inter1));
  and2  gate1221(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1222(.a(s_96), .O(gate495inter3));
  inv1  gate1223(.a(s_97), .O(gate495inter4));
  nand2 gate1224(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1225(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1226(.a(G1252), .O(gate495inter7));
  inv1  gate1227(.a(G1253), .O(gate495inter8));
  nand2 gate1228(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1229(.a(s_97), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1230(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1231(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1232(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule