module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2045(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2046(.a(gate9inter0), .b(s_214), .O(gate9inter1));
  and2  gate2047(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2048(.a(s_214), .O(gate9inter3));
  inv1  gate2049(.a(s_215), .O(gate9inter4));
  nand2 gate2050(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2051(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2052(.a(G1), .O(gate9inter7));
  inv1  gate2053(.a(G2), .O(gate9inter8));
  nand2 gate2054(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2055(.a(s_215), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2056(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2057(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2058(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1191(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1192(.a(gate12inter0), .b(s_92), .O(gate12inter1));
  and2  gate1193(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1194(.a(s_92), .O(gate12inter3));
  inv1  gate1195(.a(s_93), .O(gate12inter4));
  nand2 gate1196(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1197(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1198(.a(G7), .O(gate12inter7));
  inv1  gate1199(.a(G8), .O(gate12inter8));
  nand2 gate1200(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1201(.a(s_93), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1202(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1203(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1204(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate701(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate702(.a(gate13inter0), .b(s_22), .O(gate13inter1));
  and2  gate703(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate704(.a(s_22), .O(gate13inter3));
  inv1  gate705(.a(s_23), .O(gate13inter4));
  nand2 gate706(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate707(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate708(.a(G9), .O(gate13inter7));
  inv1  gate709(.a(G10), .O(gate13inter8));
  nand2 gate710(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate711(.a(s_23), .b(gate13inter3), .O(gate13inter10));
  nor2  gate712(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate713(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate714(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate855(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate856(.a(gate16inter0), .b(s_44), .O(gate16inter1));
  and2  gate857(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate858(.a(s_44), .O(gate16inter3));
  inv1  gate859(.a(s_45), .O(gate16inter4));
  nand2 gate860(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate861(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate862(.a(G15), .O(gate16inter7));
  inv1  gate863(.a(G16), .O(gate16inter8));
  nand2 gate864(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate865(.a(s_45), .b(gate16inter3), .O(gate16inter10));
  nor2  gate866(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate867(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate868(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate631(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate632(.a(gate19inter0), .b(s_12), .O(gate19inter1));
  and2  gate633(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate634(.a(s_12), .O(gate19inter3));
  inv1  gate635(.a(s_13), .O(gate19inter4));
  nand2 gate636(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate637(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate638(.a(G21), .O(gate19inter7));
  inv1  gate639(.a(G22), .O(gate19inter8));
  nand2 gate640(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate641(.a(s_13), .b(gate19inter3), .O(gate19inter10));
  nor2  gate642(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate643(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate644(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1933(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1934(.a(gate23inter0), .b(s_198), .O(gate23inter1));
  and2  gate1935(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1936(.a(s_198), .O(gate23inter3));
  inv1  gate1937(.a(s_199), .O(gate23inter4));
  nand2 gate1938(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1939(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1940(.a(G29), .O(gate23inter7));
  inv1  gate1941(.a(G30), .O(gate23inter8));
  nand2 gate1942(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1943(.a(s_199), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1944(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1945(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1946(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1275(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1276(.a(gate25inter0), .b(s_104), .O(gate25inter1));
  and2  gate1277(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1278(.a(s_104), .O(gate25inter3));
  inv1  gate1279(.a(s_105), .O(gate25inter4));
  nand2 gate1280(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1281(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1282(.a(G1), .O(gate25inter7));
  inv1  gate1283(.a(G5), .O(gate25inter8));
  nand2 gate1284(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1285(.a(s_105), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1286(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1287(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1288(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1163(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1164(.a(gate28inter0), .b(s_88), .O(gate28inter1));
  and2  gate1165(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1166(.a(s_88), .O(gate28inter3));
  inv1  gate1167(.a(s_89), .O(gate28inter4));
  nand2 gate1168(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1169(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1170(.a(G10), .O(gate28inter7));
  inv1  gate1171(.a(G14), .O(gate28inter8));
  nand2 gate1172(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1173(.a(s_89), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1174(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1175(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1176(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1905(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1906(.a(gate29inter0), .b(s_194), .O(gate29inter1));
  and2  gate1907(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1908(.a(s_194), .O(gate29inter3));
  inv1  gate1909(.a(s_195), .O(gate29inter4));
  nand2 gate1910(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1911(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1912(.a(G3), .O(gate29inter7));
  inv1  gate1913(.a(G7), .O(gate29inter8));
  nand2 gate1914(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1915(.a(s_195), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1916(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1917(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1918(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1989(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1990(.a(gate30inter0), .b(s_206), .O(gate30inter1));
  and2  gate1991(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1992(.a(s_206), .O(gate30inter3));
  inv1  gate1993(.a(s_207), .O(gate30inter4));
  nand2 gate1994(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1995(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1996(.a(G11), .O(gate30inter7));
  inv1  gate1997(.a(G15), .O(gate30inter8));
  nand2 gate1998(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1999(.a(s_207), .b(gate30inter3), .O(gate30inter10));
  nor2  gate2000(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate2001(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate2002(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1877(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1878(.a(gate31inter0), .b(s_190), .O(gate31inter1));
  and2  gate1879(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1880(.a(s_190), .O(gate31inter3));
  inv1  gate1881(.a(s_191), .O(gate31inter4));
  nand2 gate1882(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1883(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1884(.a(G4), .O(gate31inter7));
  inv1  gate1885(.a(G8), .O(gate31inter8));
  nand2 gate1886(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1887(.a(s_191), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1888(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1889(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1890(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1415(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1416(.a(gate33inter0), .b(s_124), .O(gate33inter1));
  and2  gate1417(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1418(.a(s_124), .O(gate33inter3));
  inv1  gate1419(.a(s_125), .O(gate33inter4));
  nand2 gate1420(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1421(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1422(.a(G17), .O(gate33inter7));
  inv1  gate1423(.a(G21), .O(gate33inter8));
  nand2 gate1424(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1425(.a(s_125), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1426(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1427(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1428(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1709(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1710(.a(gate37inter0), .b(s_166), .O(gate37inter1));
  and2  gate1711(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1712(.a(s_166), .O(gate37inter3));
  inv1  gate1713(.a(s_167), .O(gate37inter4));
  nand2 gate1714(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1715(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1716(.a(G19), .O(gate37inter7));
  inv1  gate1717(.a(G23), .O(gate37inter8));
  nand2 gate1718(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1719(.a(s_167), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1720(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1721(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1722(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1149(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1150(.a(gate45inter0), .b(s_86), .O(gate45inter1));
  and2  gate1151(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1152(.a(s_86), .O(gate45inter3));
  inv1  gate1153(.a(s_87), .O(gate45inter4));
  nand2 gate1154(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1155(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1156(.a(G5), .O(gate45inter7));
  inv1  gate1157(.a(G272), .O(gate45inter8));
  nand2 gate1158(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1159(.a(s_87), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1160(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1161(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1162(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1919(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1920(.a(gate53inter0), .b(s_196), .O(gate53inter1));
  and2  gate1921(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1922(.a(s_196), .O(gate53inter3));
  inv1  gate1923(.a(s_197), .O(gate53inter4));
  nand2 gate1924(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1925(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1926(.a(G13), .O(gate53inter7));
  inv1  gate1927(.a(G284), .O(gate53inter8));
  nand2 gate1928(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1929(.a(s_197), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1930(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1931(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1932(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate2129(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate2130(.a(gate55inter0), .b(s_226), .O(gate55inter1));
  and2  gate2131(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate2132(.a(s_226), .O(gate55inter3));
  inv1  gate2133(.a(s_227), .O(gate55inter4));
  nand2 gate2134(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate2135(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate2136(.a(G15), .O(gate55inter7));
  inv1  gate2137(.a(G287), .O(gate55inter8));
  nand2 gate2138(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate2139(.a(s_227), .b(gate55inter3), .O(gate55inter10));
  nor2  gate2140(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate2141(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate2142(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2073(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2074(.a(gate62inter0), .b(s_218), .O(gate62inter1));
  and2  gate2075(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2076(.a(s_218), .O(gate62inter3));
  inv1  gate2077(.a(s_219), .O(gate62inter4));
  nand2 gate2078(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2079(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2080(.a(G22), .O(gate62inter7));
  inv1  gate2081(.a(G296), .O(gate62inter8));
  nand2 gate2082(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2083(.a(s_219), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2084(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2085(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2086(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2003(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2004(.a(gate63inter0), .b(s_208), .O(gate63inter1));
  and2  gate2005(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2006(.a(s_208), .O(gate63inter3));
  inv1  gate2007(.a(s_209), .O(gate63inter4));
  nand2 gate2008(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2009(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2010(.a(G23), .O(gate63inter7));
  inv1  gate2011(.a(G299), .O(gate63inter8));
  nand2 gate2012(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2013(.a(s_209), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2014(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2015(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2016(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate2115(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2116(.a(gate65inter0), .b(s_224), .O(gate65inter1));
  and2  gate2117(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2118(.a(s_224), .O(gate65inter3));
  inv1  gate2119(.a(s_225), .O(gate65inter4));
  nand2 gate2120(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2121(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2122(.a(G25), .O(gate65inter7));
  inv1  gate2123(.a(G302), .O(gate65inter8));
  nand2 gate2124(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2125(.a(s_225), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2126(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2127(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2128(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1723(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1724(.a(gate67inter0), .b(s_168), .O(gate67inter1));
  and2  gate1725(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1726(.a(s_168), .O(gate67inter3));
  inv1  gate1727(.a(s_169), .O(gate67inter4));
  nand2 gate1728(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1729(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1730(.a(G27), .O(gate67inter7));
  inv1  gate1731(.a(G305), .O(gate67inter8));
  nand2 gate1732(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1733(.a(s_169), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1734(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1735(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1736(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2157(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2158(.a(gate71inter0), .b(s_230), .O(gate71inter1));
  and2  gate2159(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2160(.a(s_230), .O(gate71inter3));
  inv1  gate2161(.a(s_231), .O(gate71inter4));
  nand2 gate2162(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2163(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2164(.a(G31), .O(gate71inter7));
  inv1  gate2165(.a(G311), .O(gate71inter8));
  nand2 gate2166(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2167(.a(s_231), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2168(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2169(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2170(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1429(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1430(.a(gate72inter0), .b(s_126), .O(gate72inter1));
  and2  gate1431(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1432(.a(s_126), .O(gate72inter3));
  inv1  gate1433(.a(s_127), .O(gate72inter4));
  nand2 gate1434(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1435(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1436(.a(G32), .O(gate72inter7));
  inv1  gate1437(.a(G311), .O(gate72inter8));
  nand2 gate1438(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1439(.a(s_127), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1440(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1441(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1442(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate547(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate548(.a(gate73inter0), .b(s_0), .O(gate73inter1));
  and2  gate549(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate550(.a(s_0), .O(gate73inter3));
  inv1  gate551(.a(s_1), .O(gate73inter4));
  nand2 gate552(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate553(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate554(.a(G1), .O(gate73inter7));
  inv1  gate555(.a(G314), .O(gate73inter8));
  nand2 gate556(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate557(.a(s_1), .b(gate73inter3), .O(gate73inter10));
  nor2  gate558(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate559(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate560(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1891(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1892(.a(gate75inter0), .b(s_192), .O(gate75inter1));
  and2  gate1893(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1894(.a(s_192), .O(gate75inter3));
  inv1  gate1895(.a(s_193), .O(gate75inter4));
  nand2 gate1896(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1897(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1898(.a(G9), .O(gate75inter7));
  inv1  gate1899(.a(G317), .O(gate75inter8));
  nand2 gate1900(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1901(.a(s_193), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1902(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1903(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1904(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2031(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2032(.a(gate79inter0), .b(s_212), .O(gate79inter1));
  and2  gate2033(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2034(.a(s_212), .O(gate79inter3));
  inv1  gate2035(.a(s_213), .O(gate79inter4));
  nand2 gate2036(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2037(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2038(.a(G10), .O(gate79inter7));
  inv1  gate2039(.a(G323), .O(gate79inter8));
  nand2 gate2040(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2041(.a(s_213), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2042(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2043(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2044(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate687(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate688(.a(gate82inter0), .b(s_20), .O(gate82inter1));
  and2  gate689(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate690(.a(s_20), .O(gate82inter3));
  inv1  gate691(.a(s_21), .O(gate82inter4));
  nand2 gate692(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate693(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate694(.a(G7), .O(gate82inter7));
  inv1  gate695(.a(G326), .O(gate82inter8));
  nand2 gate696(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate697(.a(s_21), .b(gate82inter3), .O(gate82inter10));
  nor2  gate698(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate699(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate700(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1541(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1542(.a(gate85inter0), .b(s_142), .O(gate85inter1));
  and2  gate1543(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1544(.a(s_142), .O(gate85inter3));
  inv1  gate1545(.a(s_143), .O(gate85inter4));
  nand2 gate1546(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1547(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1548(.a(G4), .O(gate85inter7));
  inv1  gate1549(.a(G332), .O(gate85inter8));
  nand2 gate1550(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1551(.a(s_143), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1552(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1553(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1554(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1975(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1976(.a(gate90inter0), .b(s_204), .O(gate90inter1));
  and2  gate1977(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1978(.a(s_204), .O(gate90inter3));
  inv1  gate1979(.a(s_205), .O(gate90inter4));
  nand2 gate1980(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1981(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1982(.a(G21), .O(gate90inter7));
  inv1  gate1983(.a(G338), .O(gate90inter8));
  nand2 gate1984(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1985(.a(s_205), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1986(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1987(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1988(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate589(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate590(.a(gate96inter0), .b(s_6), .O(gate96inter1));
  and2  gate591(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate592(.a(s_6), .O(gate96inter3));
  inv1  gate593(.a(s_7), .O(gate96inter4));
  nand2 gate594(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate595(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate596(.a(G30), .O(gate96inter7));
  inv1  gate597(.a(G347), .O(gate96inter8));
  nand2 gate598(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate599(.a(s_7), .b(gate96inter3), .O(gate96inter10));
  nor2  gate600(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate601(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate602(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2101(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2102(.a(gate97inter0), .b(s_222), .O(gate97inter1));
  and2  gate2103(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2104(.a(s_222), .O(gate97inter3));
  inv1  gate2105(.a(s_223), .O(gate97inter4));
  nand2 gate2106(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2107(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2108(.a(G19), .O(gate97inter7));
  inv1  gate2109(.a(G350), .O(gate97inter8));
  nand2 gate2110(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2111(.a(s_223), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2112(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2113(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2114(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1051(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1052(.a(gate99inter0), .b(s_72), .O(gate99inter1));
  and2  gate1053(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1054(.a(s_72), .O(gate99inter3));
  inv1  gate1055(.a(s_73), .O(gate99inter4));
  nand2 gate1056(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1057(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1058(.a(G27), .O(gate99inter7));
  inv1  gate1059(.a(G353), .O(gate99inter8));
  nand2 gate1060(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1061(.a(s_73), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1062(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1063(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1064(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1821(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1822(.a(gate101inter0), .b(s_182), .O(gate101inter1));
  and2  gate1823(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1824(.a(s_182), .O(gate101inter3));
  inv1  gate1825(.a(s_183), .O(gate101inter4));
  nand2 gate1826(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1827(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1828(.a(G20), .O(gate101inter7));
  inv1  gate1829(.a(G356), .O(gate101inter8));
  nand2 gate1830(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1831(.a(s_183), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1832(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1833(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1834(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate897(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate898(.a(gate105inter0), .b(s_50), .O(gate105inter1));
  and2  gate899(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate900(.a(s_50), .O(gate105inter3));
  inv1  gate901(.a(s_51), .O(gate105inter4));
  nand2 gate902(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate903(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate904(.a(G362), .O(gate105inter7));
  inv1  gate905(.a(G363), .O(gate105inter8));
  nand2 gate906(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate907(.a(s_51), .b(gate105inter3), .O(gate105inter10));
  nor2  gate908(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate909(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate910(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1597(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1598(.a(gate107inter0), .b(s_150), .O(gate107inter1));
  and2  gate1599(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1600(.a(s_150), .O(gate107inter3));
  inv1  gate1601(.a(s_151), .O(gate107inter4));
  nand2 gate1602(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1603(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1604(.a(G366), .O(gate107inter7));
  inv1  gate1605(.a(G367), .O(gate107inter8));
  nand2 gate1606(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1607(.a(s_151), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1608(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1609(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1610(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate967(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate968(.a(gate115inter0), .b(s_60), .O(gate115inter1));
  and2  gate969(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate970(.a(s_60), .O(gate115inter3));
  inv1  gate971(.a(s_61), .O(gate115inter4));
  nand2 gate972(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate973(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate974(.a(G382), .O(gate115inter7));
  inv1  gate975(.a(G383), .O(gate115inter8));
  nand2 gate976(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate977(.a(s_61), .b(gate115inter3), .O(gate115inter10));
  nor2  gate978(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate979(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate980(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1331(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1332(.a(gate121inter0), .b(s_112), .O(gate121inter1));
  and2  gate1333(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1334(.a(s_112), .O(gate121inter3));
  inv1  gate1335(.a(s_113), .O(gate121inter4));
  nand2 gate1336(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1337(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1338(.a(G394), .O(gate121inter7));
  inv1  gate1339(.a(G395), .O(gate121inter8));
  nand2 gate1340(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1341(.a(s_113), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1342(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1343(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1344(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate561(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate562(.a(gate129inter0), .b(s_2), .O(gate129inter1));
  and2  gate563(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate564(.a(s_2), .O(gate129inter3));
  inv1  gate565(.a(s_3), .O(gate129inter4));
  nand2 gate566(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate567(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate568(.a(G410), .O(gate129inter7));
  inv1  gate569(.a(G411), .O(gate129inter8));
  nand2 gate570(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate571(.a(s_3), .b(gate129inter3), .O(gate129inter10));
  nor2  gate572(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate573(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate574(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate841(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate842(.a(gate139inter0), .b(s_42), .O(gate139inter1));
  and2  gate843(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate844(.a(s_42), .O(gate139inter3));
  inv1  gate845(.a(s_43), .O(gate139inter4));
  nand2 gate846(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate847(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate848(.a(G438), .O(gate139inter7));
  inv1  gate849(.a(G441), .O(gate139inter8));
  nand2 gate850(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate851(.a(s_43), .b(gate139inter3), .O(gate139inter10));
  nor2  gate852(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate853(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate854(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2087(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2088(.a(gate146inter0), .b(s_220), .O(gate146inter1));
  and2  gate2089(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2090(.a(s_220), .O(gate146inter3));
  inv1  gate2091(.a(s_221), .O(gate146inter4));
  nand2 gate2092(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2093(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2094(.a(G480), .O(gate146inter7));
  inv1  gate2095(.a(G483), .O(gate146inter8));
  nand2 gate2096(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2097(.a(s_221), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2098(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2099(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2100(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate785(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate786(.a(gate149inter0), .b(s_34), .O(gate149inter1));
  and2  gate787(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate788(.a(s_34), .O(gate149inter3));
  inv1  gate789(.a(s_35), .O(gate149inter4));
  nand2 gate790(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate791(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate792(.a(G498), .O(gate149inter7));
  inv1  gate793(.a(G501), .O(gate149inter8));
  nand2 gate794(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate795(.a(s_35), .b(gate149inter3), .O(gate149inter10));
  nor2  gate796(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate797(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate798(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1359(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1360(.a(gate155inter0), .b(s_116), .O(gate155inter1));
  and2  gate1361(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1362(.a(s_116), .O(gate155inter3));
  inv1  gate1363(.a(s_117), .O(gate155inter4));
  nand2 gate1364(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1365(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1366(.a(G432), .O(gate155inter7));
  inv1  gate1367(.a(G525), .O(gate155inter8));
  nand2 gate1368(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1369(.a(s_117), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1370(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1371(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1372(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1751(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1752(.a(gate158inter0), .b(s_172), .O(gate158inter1));
  and2  gate1753(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1754(.a(s_172), .O(gate158inter3));
  inv1  gate1755(.a(s_173), .O(gate158inter4));
  nand2 gate1756(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1757(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1758(.a(G441), .O(gate158inter7));
  inv1  gate1759(.a(G528), .O(gate158inter8));
  nand2 gate1760(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1761(.a(s_173), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1762(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1763(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1764(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate715(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate716(.a(gate160inter0), .b(s_24), .O(gate160inter1));
  and2  gate717(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate718(.a(s_24), .O(gate160inter3));
  inv1  gate719(.a(s_25), .O(gate160inter4));
  nand2 gate720(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate721(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate722(.a(G447), .O(gate160inter7));
  inv1  gate723(.a(G531), .O(gate160inter8));
  nand2 gate724(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate725(.a(s_25), .b(gate160inter3), .O(gate160inter10));
  nor2  gate726(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate727(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate728(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1569(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1570(.a(gate163inter0), .b(s_146), .O(gate163inter1));
  and2  gate1571(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1572(.a(s_146), .O(gate163inter3));
  inv1  gate1573(.a(s_147), .O(gate163inter4));
  nand2 gate1574(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1575(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1576(.a(G456), .O(gate163inter7));
  inv1  gate1577(.a(G537), .O(gate163inter8));
  nand2 gate1578(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1579(.a(s_147), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1580(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1581(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1582(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1513(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1514(.a(gate165inter0), .b(s_138), .O(gate165inter1));
  and2  gate1515(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1516(.a(s_138), .O(gate165inter3));
  inv1  gate1517(.a(s_139), .O(gate165inter4));
  nand2 gate1518(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1519(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1520(.a(G462), .O(gate165inter7));
  inv1  gate1521(.a(G540), .O(gate165inter8));
  nand2 gate1522(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1523(.a(s_139), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1524(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1525(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1526(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1121(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1122(.a(gate167inter0), .b(s_82), .O(gate167inter1));
  and2  gate1123(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1124(.a(s_82), .O(gate167inter3));
  inv1  gate1125(.a(s_83), .O(gate167inter4));
  nand2 gate1126(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1127(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1128(.a(G468), .O(gate167inter7));
  inv1  gate1129(.a(G543), .O(gate167inter8));
  nand2 gate1130(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1131(.a(s_83), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1132(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1133(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1134(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1289(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1290(.a(gate168inter0), .b(s_106), .O(gate168inter1));
  and2  gate1291(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1292(.a(s_106), .O(gate168inter3));
  inv1  gate1293(.a(s_107), .O(gate168inter4));
  nand2 gate1294(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1295(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1296(.a(G471), .O(gate168inter7));
  inv1  gate1297(.a(G543), .O(gate168inter8));
  nand2 gate1298(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1299(.a(s_107), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1300(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1301(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1302(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1093(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1094(.a(gate176inter0), .b(s_78), .O(gate176inter1));
  and2  gate1095(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1096(.a(s_78), .O(gate176inter3));
  inv1  gate1097(.a(s_79), .O(gate176inter4));
  nand2 gate1098(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1099(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1100(.a(G495), .O(gate176inter7));
  inv1  gate1101(.a(G555), .O(gate176inter8));
  nand2 gate1102(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1103(.a(s_79), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1104(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1105(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1106(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1863(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1864(.a(gate182inter0), .b(s_188), .O(gate182inter1));
  and2  gate1865(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1866(.a(s_188), .O(gate182inter3));
  inv1  gate1867(.a(s_189), .O(gate182inter4));
  nand2 gate1868(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1869(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1870(.a(G513), .O(gate182inter7));
  inv1  gate1871(.a(G564), .O(gate182inter8));
  nand2 gate1872(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1873(.a(s_189), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1874(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1875(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1876(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1205(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1206(.a(gate183inter0), .b(s_94), .O(gate183inter1));
  and2  gate1207(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1208(.a(s_94), .O(gate183inter3));
  inv1  gate1209(.a(s_95), .O(gate183inter4));
  nand2 gate1210(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1211(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1212(.a(G516), .O(gate183inter7));
  inv1  gate1213(.a(G567), .O(gate183inter8));
  nand2 gate1214(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1215(.a(s_95), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1216(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1217(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1218(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1485(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1486(.a(gate186inter0), .b(s_134), .O(gate186inter1));
  and2  gate1487(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1488(.a(s_134), .O(gate186inter3));
  inv1  gate1489(.a(s_135), .O(gate186inter4));
  nand2 gate1490(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1491(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1492(.a(G572), .O(gate186inter7));
  inv1  gate1493(.a(G573), .O(gate186inter8));
  nand2 gate1494(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1495(.a(s_135), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1496(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1497(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1498(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1779(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1780(.a(gate193inter0), .b(s_176), .O(gate193inter1));
  and2  gate1781(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1782(.a(s_176), .O(gate193inter3));
  inv1  gate1783(.a(s_177), .O(gate193inter4));
  nand2 gate1784(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1785(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1786(.a(G586), .O(gate193inter7));
  inv1  gate1787(.a(G587), .O(gate193inter8));
  nand2 gate1788(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1789(.a(s_177), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1790(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1791(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1792(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1317(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1318(.a(gate195inter0), .b(s_110), .O(gate195inter1));
  and2  gate1319(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1320(.a(s_110), .O(gate195inter3));
  inv1  gate1321(.a(s_111), .O(gate195inter4));
  nand2 gate1322(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1323(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1324(.a(G590), .O(gate195inter7));
  inv1  gate1325(.a(G591), .O(gate195inter8));
  nand2 gate1326(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1327(.a(s_111), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1328(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1329(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1330(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1639(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1640(.a(gate199inter0), .b(s_156), .O(gate199inter1));
  and2  gate1641(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1642(.a(s_156), .O(gate199inter3));
  inv1  gate1643(.a(s_157), .O(gate199inter4));
  nand2 gate1644(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1645(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1646(.a(G598), .O(gate199inter7));
  inv1  gate1647(.a(G599), .O(gate199inter8));
  nand2 gate1648(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1649(.a(s_157), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1650(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1651(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1652(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate827(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate828(.a(gate200inter0), .b(s_40), .O(gate200inter1));
  and2  gate829(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate830(.a(s_40), .O(gate200inter3));
  inv1  gate831(.a(s_41), .O(gate200inter4));
  nand2 gate832(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate833(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate834(.a(G600), .O(gate200inter7));
  inv1  gate835(.a(G601), .O(gate200inter8));
  nand2 gate836(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate837(.a(s_41), .b(gate200inter3), .O(gate200inter10));
  nor2  gate838(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate839(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate840(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1583(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1584(.a(gate203inter0), .b(s_148), .O(gate203inter1));
  and2  gate1585(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1586(.a(s_148), .O(gate203inter3));
  inv1  gate1587(.a(s_149), .O(gate203inter4));
  nand2 gate1588(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1589(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1590(.a(G602), .O(gate203inter7));
  inv1  gate1591(.a(G612), .O(gate203inter8));
  nand2 gate1592(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1593(.a(s_149), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1594(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1595(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1596(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate799(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate800(.a(gate206inter0), .b(s_36), .O(gate206inter1));
  and2  gate801(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate802(.a(s_36), .O(gate206inter3));
  inv1  gate803(.a(s_37), .O(gate206inter4));
  nand2 gate804(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate805(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate806(.a(G632), .O(gate206inter7));
  inv1  gate807(.a(G637), .O(gate206inter8));
  nand2 gate808(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate809(.a(s_37), .b(gate206inter3), .O(gate206inter10));
  nor2  gate810(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate811(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate812(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate981(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate982(.a(gate209inter0), .b(s_62), .O(gate209inter1));
  and2  gate983(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate984(.a(s_62), .O(gate209inter3));
  inv1  gate985(.a(s_63), .O(gate209inter4));
  nand2 gate986(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate987(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate988(.a(G602), .O(gate209inter7));
  inv1  gate989(.a(G666), .O(gate209inter8));
  nand2 gate990(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate991(.a(s_63), .b(gate209inter3), .O(gate209inter10));
  nor2  gate992(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate993(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate994(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1961(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1962(.a(gate213inter0), .b(s_202), .O(gate213inter1));
  and2  gate1963(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1964(.a(s_202), .O(gate213inter3));
  inv1  gate1965(.a(s_203), .O(gate213inter4));
  nand2 gate1966(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1967(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1968(.a(G602), .O(gate213inter7));
  inv1  gate1969(.a(G672), .O(gate213inter8));
  nand2 gate1970(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1971(.a(s_203), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1972(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1973(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1974(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1233(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1234(.a(gate221inter0), .b(s_98), .O(gate221inter1));
  and2  gate1235(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1236(.a(s_98), .O(gate221inter3));
  inv1  gate1237(.a(s_99), .O(gate221inter4));
  nand2 gate1238(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1239(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1240(.a(G622), .O(gate221inter7));
  inv1  gate1241(.a(G684), .O(gate221inter8));
  nand2 gate1242(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1243(.a(s_99), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1244(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1245(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1246(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1247(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1248(.a(gate233inter0), .b(s_100), .O(gate233inter1));
  and2  gate1249(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1250(.a(s_100), .O(gate233inter3));
  inv1  gate1251(.a(s_101), .O(gate233inter4));
  nand2 gate1252(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1253(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1254(.a(G242), .O(gate233inter7));
  inv1  gate1255(.a(G718), .O(gate233inter8));
  nand2 gate1256(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1257(.a(s_101), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1258(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1259(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1260(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1835(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1836(.a(gate241inter0), .b(s_184), .O(gate241inter1));
  and2  gate1837(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1838(.a(s_184), .O(gate241inter3));
  inv1  gate1839(.a(s_185), .O(gate241inter4));
  nand2 gate1840(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1841(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1842(.a(G242), .O(gate241inter7));
  inv1  gate1843(.a(G730), .O(gate241inter8));
  nand2 gate1844(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1845(.a(s_185), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1846(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1847(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1848(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate953(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate954(.a(gate247inter0), .b(s_58), .O(gate247inter1));
  and2  gate955(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate956(.a(s_58), .O(gate247inter3));
  inv1  gate957(.a(s_59), .O(gate247inter4));
  nand2 gate958(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate959(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate960(.a(G251), .O(gate247inter7));
  inv1  gate961(.a(G739), .O(gate247inter8));
  nand2 gate962(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate963(.a(s_59), .b(gate247inter3), .O(gate247inter10));
  nor2  gate964(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate965(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate966(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1443(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1444(.a(gate248inter0), .b(s_128), .O(gate248inter1));
  and2  gate1445(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1446(.a(s_128), .O(gate248inter3));
  inv1  gate1447(.a(s_129), .O(gate248inter4));
  nand2 gate1448(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1449(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1450(.a(G727), .O(gate248inter7));
  inv1  gate1451(.a(G739), .O(gate248inter8));
  nand2 gate1452(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1453(.a(s_129), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1454(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1455(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1456(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1345(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1346(.a(gate251inter0), .b(s_114), .O(gate251inter1));
  and2  gate1347(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1348(.a(s_114), .O(gate251inter3));
  inv1  gate1349(.a(s_115), .O(gate251inter4));
  nand2 gate1350(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1351(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1352(.a(G257), .O(gate251inter7));
  inv1  gate1353(.a(G745), .O(gate251inter8));
  nand2 gate1354(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1355(.a(s_115), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1356(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1357(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1358(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1611(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1612(.a(gate258inter0), .b(s_152), .O(gate258inter1));
  and2  gate1613(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1614(.a(s_152), .O(gate258inter3));
  inv1  gate1615(.a(s_153), .O(gate258inter4));
  nand2 gate1616(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1617(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1618(.a(G756), .O(gate258inter7));
  inv1  gate1619(.a(G757), .O(gate258inter8));
  nand2 gate1620(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1621(.a(s_153), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1622(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1623(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1624(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1107(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1108(.a(gate262inter0), .b(s_80), .O(gate262inter1));
  and2  gate1109(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1110(.a(s_80), .O(gate262inter3));
  inv1  gate1111(.a(s_81), .O(gate262inter4));
  nand2 gate1112(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1113(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1114(.a(G764), .O(gate262inter7));
  inv1  gate1115(.a(G765), .O(gate262inter8));
  nand2 gate1116(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1117(.a(s_81), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1118(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1119(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1120(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate813(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate814(.a(gate265inter0), .b(s_38), .O(gate265inter1));
  and2  gate815(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate816(.a(s_38), .O(gate265inter3));
  inv1  gate817(.a(s_39), .O(gate265inter4));
  nand2 gate818(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate819(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate820(.a(G642), .O(gate265inter7));
  inv1  gate821(.a(G770), .O(gate265inter8));
  nand2 gate822(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate823(.a(s_39), .b(gate265inter3), .O(gate265inter10));
  nor2  gate824(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate825(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate826(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate771(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate772(.a(gate266inter0), .b(s_32), .O(gate266inter1));
  and2  gate773(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate774(.a(s_32), .O(gate266inter3));
  inv1  gate775(.a(s_33), .O(gate266inter4));
  nand2 gate776(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate777(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate778(.a(G645), .O(gate266inter7));
  inv1  gate779(.a(G773), .O(gate266inter8));
  nand2 gate780(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate781(.a(s_33), .b(gate266inter3), .O(gate266inter10));
  nor2  gate782(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate783(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate784(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate925(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate926(.a(gate267inter0), .b(s_54), .O(gate267inter1));
  and2  gate927(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate928(.a(s_54), .O(gate267inter3));
  inv1  gate929(.a(s_55), .O(gate267inter4));
  nand2 gate930(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate931(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate932(.a(G648), .O(gate267inter7));
  inv1  gate933(.a(G776), .O(gate267inter8));
  nand2 gate934(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate935(.a(s_55), .b(gate267inter3), .O(gate267inter10));
  nor2  gate936(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate937(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate938(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate729(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate730(.a(gate270inter0), .b(s_26), .O(gate270inter1));
  and2  gate731(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate732(.a(s_26), .O(gate270inter3));
  inv1  gate733(.a(s_27), .O(gate270inter4));
  nand2 gate734(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate735(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate736(.a(G657), .O(gate270inter7));
  inv1  gate737(.a(G785), .O(gate270inter8));
  nand2 gate738(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate739(.a(s_27), .b(gate270inter3), .O(gate270inter10));
  nor2  gate740(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate741(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate742(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate995(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate996(.a(gate271inter0), .b(s_64), .O(gate271inter1));
  and2  gate997(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate998(.a(s_64), .O(gate271inter3));
  inv1  gate999(.a(s_65), .O(gate271inter4));
  nand2 gate1000(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1001(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1002(.a(G660), .O(gate271inter7));
  inv1  gate1003(.a(G788), .O(gate271inter8));
  nand2 gate1004(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1005(.a(s_65), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1006(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1007(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1008(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1009(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1010(.a(gate272inter0), .b(s_66), .O(gate272inter1));
  and2  gate1011(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1012(.a(s_66), .O(gate272inter3));
  inv1  gate1013(.a(s_67), .O(gate272inter4));
  nand2 gate1014(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1015(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1016(.a(G663), .O(gate272inter7));
  inv1  gate1017(.a(G791), .O(gate272inter8));
  nand2 gate1018(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1019(.a(s_67), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1020(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1021(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1022(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1667(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1668(.a(gate275inter0), .b(s_160), .O(gate275inter1));
  and2  gate1669(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1670(.a(s_160), .O(gate275inter3));
  inv1  gate1671(.a(s_161), .O(gate275inter4));
  nand2 gate1672(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1673(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1674(.a(G645), .O(gate275inter7));
  inv1  gate1675(.a(G797), .O(gate275inter8));
  nand2 gate1676(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1677(.a(s_161), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1678(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1679(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1680(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate659(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate660(.a(gate276inter0), .b(s_16), .O(gate276inter1));
  and2  gate661(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate662(.a(s_16), .O(gate276inter3));
  inv1  gate663(.a(s_17), .O(gate276inter4));
  nand2 gate664(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate665(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate666(.a(G773), .O(gate276inter7));
  inv1  gate667(.a(G797), .O(gate276inter8));
  nand2 gate668(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate669(.a(s_17), .b(gate276inter3), .O(gate276inter10));
  nor2  gate670(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate671(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate672(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate869(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate870(.a(gate279inter0), .b(s_46), .O(gate279inter1));
  and2  gate871(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate872(.a(s_46), .O(gate279inter3));
  inv1  gate873(.a(s_47), .O(gate279inter4));
  nand2 gate874(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate875(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate876(.a(G651), .O(gate279inter7));
  inv1  gate877(.a(G803), .O(gate279inter8));
  nand2 gate878(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate879(.a(s_47), .b(gate279inter3), .O(gate279inter10));
  nor2  gate880(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate881(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate882(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1499(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1500(.a(gate281inter0), .b(s_136), .O(gate281inter1));
  and2  gate1501(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1502(.a(s_136), .O(gate281inter3));
  inv1  gate1503(.a(s_137), .O(gate281inter4));
  nand2 gate1504(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1505(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1506(.a(G654), .O(gate281inter7));
  inv1  gate1507(.a(G806), .O(gate281inter8));
  nand2 gate1508(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1509(.a(s_137), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1510(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1511(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1512(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1527(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1528(.a(gate284inter0), .b(s_140), .O(gate284inter1));
  and2  gate1529(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1530(.a(s_140), .O(gate284inter3));
  inv1  gate1531(.a(s_141), .O(gate284inter4));
  nand2 gate1532(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1533(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1534(.a(G785), .O(gate284inter7));
  inv1  gate1535(.a(G809), .O(gate284inter8));
  nand2 gate1536(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1537(.a(s_141), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1538(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1539(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1540(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate673(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate674(.a(gate289inter0), .b(s_18), .O(gate289inter1));
  and2  gate675(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate676(.a(s_18), .O(gate289inter3));
  inv1  gate677(.a(s_19), .O(gate289inter4));
  nand2 gate678(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate679(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate680(.a(G818), .O(gate289inter7));
  inv1  gate681(.a(G819), .O(gate289inter8));
  nand2 gate682(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate683(.a(s_19), .b(gate289inter3), .O(gate289inter10));
  nor2  gate684(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate685(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate686(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1387(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1388(.a(gate292inter0), .b(s_120), .O(gate292inter1));
  and2  gate1389(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1390(.a(s_120), .O(gate292inter3));
  inv1  gate1391(.a(s_121), .O(gate292inter4));
  nand2 gate1392(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1393(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1394(.a(G824), .O(gate292inter7));
  inv1  gate1395(.a(G825), .O(gate292inter8));
  nand2 gate1396(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1397(.a(s_121), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1398(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1399(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1400(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1947(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1948(.a(gate387inter0), .b(s_200), .O(gate387inter1));
  and2  gate1949(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1950(.a(s_200), .O(gate387inter3));
  inv1  gate1951(.a(s_201), .O(gate387inter4));
  nand2 gate1952(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1953(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1954(.a(G1), .O(gate387inter7));
  inv1  gate1955(.a(G1036), .O(gate387inter8));
  nand2 gate1956(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1957(.a(s_201), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1958(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1959(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1960(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate939(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate940(.a(gate391inter0), .b(s_56), .O(gate391inter1));
  and2  gate941(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate942(.a(s_56), .O(gate391inter3));
  inv1  gate943(.a(s_57), .O(gate391inter4));
  nand2 gate944(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate945(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate946(.a(G5), .O(gate391inter7));
  inv1  gate947(.a(G1048), .O(gate391inter8));
  nand2 gate948(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate949(.a(s_57), .b(gate391inter3), .O(gate391inter10));
  nor2  gate950(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate951(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate952(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate617(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate618(.a(gate392inter0), .b(s_10), .O(gate392inter1));
  and2  gate619(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate620(.a(s_10), .O(gate392inter3));
  inv1  gate621(.a(s_11), .O(gate392inter4));
  nand2 gate622(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate623(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate624(.a(G6), .O(gate392inter7));
  inv1  gate625(.a(G1051), .O(gate392inter8));
  nand2 gate626(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate627(.a(s_11), .b(gate392inter3), .O(gate392inter10));
  nor2  gate628(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate629(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate630(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1625(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1626(.a(gate393inter0), .b(s_154), .O(gate393inter1));
  and2  gate1627(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1628(.a(s_154), .O(gate393inter3));
  inv1  gate1629(.a(s_155), .O(gate393inter4));
  nand2 gate1630(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1631(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1632(.a(G7), .O(gate393inter7));
  inv1  gate1633(.a(G1054), .O(gate393inter8));
  nand2 gate1634(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1635(.a(s_155), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1636(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1637(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1638(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2059(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2060(.a(gate395inter0), .b(s_216), .O(gate395inter1));
  and2  gate2061(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2062(.a(s_216), .O(gate395inter3));
  inv1  gate2063(.a(s_217), .O(gate395inter4));
  nand2 gate2064(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2065(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2066(.a(G9), .O(gate395inter7));
  inv1  gate2067(.a(G1060), .O(gate395inter8));
  nand2 gate2068(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2069(.a(s_217), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2070(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2071(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2072(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1807(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1808(.a(gate396inter0), .b(s_180), .O(gate396inter1));
  and2  gate1809(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1810(.a(s_180), .O(gate396inter3));
  inv1  gate1811(.a(s_181), .O(gate396inter4));
  nand2 gate1812(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1813(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1814(.a(G10), .O(gate396inter7));
  inv1  gate1815(.a(G1063), .O(gate396inter8));
  nand2 gate1816(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1817(.a(s_181), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1818(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1819(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1820(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1023(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1024(.a(gate400inter0), .b(s_68), .O(gate400inter1));
  and2  gate1025(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1026(.a(s_68), .O(gate400inter3));
  inv1  gate1027(.a(s_69), .O(gate400inter4));
  nand2 gate1028(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1029(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1030(.a(G14), .O(gate400inter7));
  inv1  gate1031(.a(G1075), .O(gate400inter8));
  nand2 gate1032(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1033(.a(s_69), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1034(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1035(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1036(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1219(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1220(.a(gate407inter0), .b(s_96), .O(gate407inter1));
  and2  gate1221(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1222(.a(s_96), .O(gate407inter3));
  inv1  gate1223(.a(s_97), .O(gate407inter4));
  nand2 gate1224(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1225(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1226(.a(G21), .O(gate407inter7));
  inv1  gate1227(.a(G1096), .O(gate407inter8));
  nand2 gate1228(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1229(.a(s_97), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1230(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1231(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1232(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1555(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1556(.a(gate409inter0), .b(s_144), .O(gate409inter1));
  and2  gate1557(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1558(.a(s_144), .O(gate409inter3));
  inv1  gate1559(.a(s_145), .O(gate409inter4));
  nand2 gate1560(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1561(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1562(.a(G23), .O(gate409inter7));
  inv1  gate1563(.a(G1102), .O(gate409inter8));
  nand2 gate1564(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1565(.a(s_145), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1566(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1567(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1568(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1177(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1178(.a(gate411inter0), .b(s_90), .O(gate411inter1));
  and2  gate1179(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1180(.a(s_90), .O(gate411inter3));
  inv1  gate1181(.a(s_91), .O(gate411inter4));
  nand2 gate1182(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1183(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1184(.a(G25), .O(gate411inter7));
  inv1  gate1185(.a(G1108), .O(gate411inter8));
  nand2 gate1186(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1187(.a(s_91), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1188(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1189(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1190(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1457(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1458(.a(gate413inter0), .b(s_130), .O(gate413inter1));
  and2  gate1459(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1460(.a(s_130), .O(gate413inter3));
  inv1  gate1461(.a(s_131), .O(gate413inter4));
  nand2 gate1462(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1463(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1464(.a(G27), .O(gate413inter7));
  inv1  gate1465(.a(G1114), .O(gate413inter8));
  nand2 gate1466(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1467(.a(s_131), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1468(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1469(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1470(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate743(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate744(.a(gate420inter0), .b(s_28), .O(gate420inter1));
  and2  gate745(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate746(.a(s_28), .O(gate420inter3));
  inv1  gate747(.a(s_29), .O(gate420inter4));
  nand2 gate748(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate749(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate750(.a(G1036), .O(gate420inter7));
  inv1  gate751(.a(G1132), .O(gate420inter8));
  nand2 gate752(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate753(.a(s_29), .b(gate420inter3), .O(gate420inter10));
  nor2  gate754(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate755(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate756(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1079(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1080(.a(gate424inter0), .b(s_76), .O(gate424inter1));
  and2  gate1081(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1082(.a(s_76), .O(gate424inter3));
  inv1  gate1083(.a(s_77), .O(gate424inter4));
  nand2 gate1084(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1085(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1086(.a(G1042), .O(gate424inter7));
  inv1  gate1087(.a(G1138), .O(gate424inter8));
  nand2 gate1088(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1089(.a(s_77), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1090(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1091(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1092(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1037(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1038(.a(gate440inter0), .b(s_70), .O(gate440inter1));
  and2  gate1039(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1040(.a(s_70), .O(gate440inter3));
  inv1  gate1041(.a(s_71), .O(gate440inter4));
  nand2 gate1042(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1043(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1044(.a(G1066), .O(gate440inter7));
  inv1  gate1045(.a(G1162), .O(gate440inter8));
  nand2 gate1046(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1047(.a(s_71), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1048(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1049(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1050(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate2143(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2144(.a(gate441inter0), .b(s_228), .O(gate441inter1));
  and2  gate2145(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2146(.a(s_228), .O(gate441inter3));
  inv1  gate2147(.a(s_229), .O(gate441inter4));
  nand2 gate2148(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2149(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2150(.a(G12), .O(gate441inter7));
  inv1  gate2151(.a(G1165), .O(gate441inter8));
  nand2 gate2152(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2153(.a(s_229), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2154(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2155(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2156(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1849(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1850(.a(gate443inter0), .b(s_186), .O(gate443inter1));
  and2  gate1851(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1852(.a(s_186), .O(gate443inter3));
  inv1  gate1853(.a(s_187), .O(gate443inter4));
  nand2 gate1854(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1855(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1856(.a(G13), .O(gate443inter7));
  inv1  gate1857(.a(G1168), .O(gate443inter8));
  nand2 gate1858(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1859(.a(s_187), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1860(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1861(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1862(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1653(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1654(.a(gate444inter0), .b(s_158), .O(gate444inter1));
  and2  gate1655(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1656(.a(s_158), .O(gate444inter3));
  inv1  gate1657(.a(s_159), .O(gate444inter4));
  nand2 gate1658(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1659(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1660(.a(G1072), .O(gate444inter7));
  inv1  gate1661(.a(G1168), .O(gate444inter8));
  nand2 gate1662(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1663(.a(s_159), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1664(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1665(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1666(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate883(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate884(.a(gate452inter0), .b(s_48), .O(gate452inter1));
  and2  gate885(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate886(.a(s_48), .O(gate452inter3));
  inv1  gate887(.a(s_49), .O(gate452inter4));
  nand2 gate888(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate889(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate890(.a(G1084), .O(gate452inter7));
  inv1  gate891(.a(G1180), .O(gate452inter8));
  nand2 gate892(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate893(.a(s_49), .b(gate452inter3), .O(gate452inter10));
  nor2  gate894(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate895(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate896(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate1695(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1696(.a(gate453inter0), .b(s_164), .O(gate453inter1));
  and2  gate1697(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1698(.a(s_164), .O(gate453inter3));
  inv1  gate1699(.a(s_165), .O(gate453inter4));
  nand2 gate1700(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1701(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1702(.a(G18), .O(gate453inter7));
  inv1  gate1703(.a(G1183), .O(gate453inter8));
  nand2 gate1704(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1705(.a(s_165), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1706(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1707(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1708(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1401(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1402(.a(gate454inter0), .b(s_122), .O(gate454inter1));
  and2  gate1403(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1404(.a(s_122), .O(gate454inter3));
  inv1  gate1405(.a(s_123), .O(gate454inter4));
  nand2 gate1406(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1407(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1408(.a(G1087), .O(gate454inter7));
  inv1  gate1409(.a(G1183), .O(gate454inter8));
  nand2 gate1410(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1411(.a(s_123), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1412(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1413(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1414(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate757(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate758(.a(gate456inter0), .b(s_30), .O(gate456inter1));
  and2  gate759(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate760(.a(s_30), .O(gate456inter3));
  inv1  gate761(.a(s_31), .O(gate456inter4));
  nand2 gate762(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate763(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate764(.a(G1090), .O(gate456inter7));
  inv1  gate765(.a(G1186), .O(gate456inter8));
  nand2 gate766(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate767(.a(s_31), .b(gate456inter3), .O(gate456inter10));
  nor2  gate768(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate769(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate770(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1135(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1136(.a(gate463inter0), .b(s_84), .O(gate463inter1));
  and2  gate1137(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1138(.a(s_84), .O(gate463inter3));
  inv1  gate1139(.a(s_85), .O(gate463inter4));
  nand2 gate1140(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1141(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1142(.a(G23), .O(gate463inter7));
  inv1  gate1143(.a(G1198), .O(gate463inter8));
  nand2 gate1144(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1145(.a(s_85), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1146(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1147(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1148(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1793(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1794(.a(gate464inter0), .b(s_178), .O(gate464inter1));
  and2  gate1795(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1796(.a(s_178), .O(gate464inter3));
  inv1  gate1797(.a(s_179), .O(gate464inter4));
  nand2 gate1798(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1799(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1800(.a(G1102), .O(gate464inter7));
  inv1  gate1801(.a(G1198), .O(gate464inter8));
  nand2 gate1802(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1803(.a(s_179), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1804(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1805(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1806(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1681(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1682(.a(gate466inter0), .b(s_162), .O(gate466inter1));
  and2  gate1683(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1684(.a(s_162), .O(gate466inter3));
  inv1  gate1685(.a(s_163), .O(gate466inter4));
  nand2 gate1686(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1687(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1688(.a(G1105), .O(gate466inter7));
  inv1  gate1689(.a(G1201), .O(gate466inter8));
  nand2 gate1690(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1691(.a(s_163), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1692(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1693(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1694(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1373(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1374(.a(gate467inter0), .b(s_118), .O(gate467inter1));
  and2  gate1375(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1376(.a(s_118), .O(gate467inter3));
  inv1  gate1377(.a(s_119), .O(gate467inter4));
  nand2 gate1378(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1379(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1380(.a(G25), .O(gate467inter7));
  inv1  gate1381(.a(G1204), .O(gate467inter8));
  nand2 gate1382(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1383(.a(s_119), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1384(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1385(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1386(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate2017(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2018(.a(gate469inter0), .b(s_210), .O(gate469inter1));
  and2  gate2019(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2020(.a(s_210), .O(gate469inter3));
  inv1  gate2021(.a(s_211), .O(gate469inter4));
  nand2 gate2022(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2023(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2024(.a(G26), .O(gate469inter7));
  inv1  gate2025(.a(G1207), .O(gate469inter8));
  nand2 gate2026(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2027(.a(s_211), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2028(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2029(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2030(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1737(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1738(.a(gate471inter0), .b(s_170), .O(gate471inter1));
  and2  gate1739(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1740(.a(s_170), .O(gate471inter3));
  inv1  gate1741(.a(s_171), .O(gate471inter4));
  nand2 gate1742(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1743(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1744(.a(G27), .O(gate471inter7));
  inv1  gate1745(.a(G1210), .O(gate471inter8));
  nand2 gate1746(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1747(.a(s_171), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1748(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1749(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1750(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate911(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate912(.a(gate473inter0), .b(s_52), .O(gate473inter1));
  and2  gate913(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate914(.a(s_52), .O(gate473inter3));
  inv1  gate915(.a(s_53), .O(gate473inter4));
  nand2 gate916(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate917(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate918(.a(G28), .O(gate473inter7));
  inv1  gate919(.a(G1213), .O(gate473inter8));
  nand2 gate920(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate921(.a(s_53), .b(gate473inter3), .O(gate473inter10));
  nor2  gate922(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate923(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate924(.a(gate473inter12), .b(gate473inter1), .O(G1282));

  xor2  gate1261(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1262(.a(gate474inter0), .b(s_102), .O(gate474inter1));
  and2  gate1263(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1264(.a(s_102), .O(gate474inter3));
  inv1  gate1265(.a(s_103), .O(gate474inter4));
  nand2 gate1266(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1267(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1268(.a(G1117), .O(gate474inter7));
  inv1  gate1269(.a(G1213), .O(gate474inter8));
  nand2 gate1270(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1271(.a(s_103), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1272(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1273(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1274(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate645(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate646(.a(gate482inter0), .b(s_14), .O(gate482inter1));
  and2  gate647(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate648(.a(s_14), .O(gate482inter3));
  inv1  gate649(.a(s_15), .O(gate482inter4));
  nand2 gate650(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate651(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate652(.a(G1129), .O(gate482inter7));
  inv1  gate653(.a(G1225), .O(gate482inter8));
  nand2 gate654(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate655(.a(s_15), .b(gate482inter3), .O(gate482inter10));
  nor2  gate656(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate657(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate658(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1765(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1766(.a(gate485inter0), .b(s_174), .O(gate485inter1));
  and2  gate1767(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1768(.a(s_174), .O(gate485inter3));
  inv1  gate1769(.a(s_175), .O(gate485inter4));
  nand2 gate1770(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1771(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1772(.a(G1232), .O(gate485inter7));
  inv1  gate1773(.a(G1233), .O(gate485inter8));
  nand2 gate1774(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1775(.a(s_175), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1776(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1777(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1778(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate575(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate576(.a(gate488inter0), .b(s_4), .O(gate488inter1));
  and2  gate577(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate578(.a(s_4), .O(gate488inter3));
  inv1  gate579(.a(s_5), .O(gate488inter4));
  nand2 gate580(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate581(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate582(.a(G1238), .O(gate488inter7));
  inv1  gate583(.a(G1239), .O(gate488inter8));
  nand2 gate584(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate585(.a(s_5), .b(gate488inter3), .O(gate488inter10));
  nor2  gate586(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate587(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate588(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate603(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate604(.a(gate489inter0), .b(s_8), .O(gate489inter1));
  and2  gate605(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate606(.a(s_8), .O(gate489inter3));
  inv1  gate607(.a(s_9), .O(gate489inter4));
  nand2 gate608(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate609(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate610(.a(G1240), .O(gate489inter7));
  inv1  gate611(.a(G1241), .O(gate489inter8));
  nand2 gate612(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate613(.a(s_9), .b(gate489inter3), .O(gate489inter10));
  nor2  gate614(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate615(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate616(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1065(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1066(.a(gate491inter0), .b(s_74), .O(gate491inter1));
  and2  gate1067(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1068(.a(s_74), .O(gate491inter3));
  inv1  gate1069(.a(s_75), .O(gate491inter4));
  nand2 gate1070(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1071(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1072(.a(G1244), .O(gate491inter7));
  inv1  gate1073(.a(G1245), .O(gate491inter8));
  nand2 gate1074(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1075(.a(s_75), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1076(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1077(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1078(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1303(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1304(.a(gate501inter0), .b(s_108), .O(gate501inter1));
  and2  gate1305(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1306(.a(s_108), .O(gate501inter3));
  inv1  gate1307(.a(s_109), .O(gate501inter4));
  nand2 gate1308(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1309(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1310(.a(G1264), .O(gate501inter7));
  inv1  gate1311(.a(G1265), .O(gate501inter8));
  nand2 gate1312(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1313(.a(s_109), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1314(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1315(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1316(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1471(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1472(.a(gate508inter0), .b(s_132), .O(gate508inter1));
  and2  gate1473(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1474(.a(s_132), .O(gate508inter3));
  inv1  gate1475(.a(s_133), .O(gate508inter4));
  nand2 gate1476(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1477(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1478(.a(G1278), .O(gate508inter7));
  inv1  gate1479(.a(G1279), .O(gate508inter8));
  nand2 gate1480(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1481(.a(s_133), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1482(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1483(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1484(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule