module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );

  xor2  gate273(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate274(.a(gate20inter0), .b(s_16), .O(gate20inter1));
  and2  gate275(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate276(.a(s_16), .O(gate20inter3));
  inv1  gate277(.a(s_17), .O(gate20inter4));
  nand2 gate278(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate279(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate280(.a(N8), .O(gate20inter7));
  inv1  gate281(.a(N119), .O(gate20inter8));
  nand2 gate282(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate283(.a(s_17), .b(gate20inter3), .O(gate20inter10));
  nor2  gate284(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate285(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate286(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );

  xor2  gate329(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate330(.a(gate22inter0), .b(s_24), .O(gate22inter1));
  and2  gate331(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate332(.a(s_24), .O(gate22inter3));
  inv1  gate333(.a(s_25), .O(gate22inter4));
  nand2 gate334(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate335(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate336(.a(N122), .O(gate22inter7));
  inv1  gate337(.a(N17), .O(gate22inter8));
  nand2 gate338(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate339(.a(s_25), .b(gate22inter3), .O(gate22inter10));
  nor2  gate340(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate341(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate342(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );

  xor2  gate203(.a(N56), .b(N134), .O(gate25inter0));
  nand2 gate204(.a(gate25inter0), .b(s_6), .O(gate25inter1));
  and2  gate205(.a(N56), .b(N134), .O(gate25inter2));
  inv1  gate206(.a(s_6), .O(gate25inter3));
  inv1  gate207(.a(s_7), .O(gate25inter4));
  nand2 gate208(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate209(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate210(.a(N134), .O(gate25inter7));
  inv1  gate211(.a(N56), .O(gate25inter8));
  nand2 gate212(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate213(.a(s_7), .b(gate25inter3), .O(gate25inter10));
  nor2  gate214(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate215(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate216(.a(gate25inter12), .b(gate25inter1), .O(N168));
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate217(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate218(.a(gate29inter0), .b(s_8), .O(gate29inter1));
  and2  gate219(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate220(.a(s_8), .O(gate29inter3));
  inv1  gate221(.a(s_9), .O(gate29inter4));
  nand2 gate222(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate223(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate224(.a(N150), .O(gate29inter7));
  inv1  gate225(.a(N108), .O(gate29inter8));
  nand2 gate226(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate227(.a(s_9), .b(gate29inter3), .O(gate29inter10));
  nor2  gate228(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate229(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate230(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );

  xor2  gate259(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate260(.a(gate31inter0), .b(s_14), .O(gate31inter1));
  and2  gate261(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate262(.a(s_14), .O(gate31inter3));
  inv1  gate263(.a(s_15), .O(gate31inter4));
  nand2 gate264(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate265(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate266(.a(N27), .O(gate31inter7));
  inv1  gate267(.a(N123), .O(gate31inter8));
  nand2 gate268(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate269(.a(s_15), .b(gate31inter3), .O(gate31inter10));
  nor2  gate270(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate271(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate272(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate371(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate372(.a(gate40inter0), .b(s_30), .O(gate40inter1));
  and2  gate373(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate374(.a(s_30), .O(gate40inter3));
  inv1  gate375(.a(s_31), .O(gate40inter4));
  nand2 gate376(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate377(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate378(.a(N86), .O(gate40inter7));
  inv1  gate379(.a(N143), .O(gate40inter8));
  nand2 gate380(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate381(.a(s_31), .b(gate40inter3), .O(gate40inter10));
  nor2  gate382(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate383(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate384(.a(gate40inter12), .b(gate40inter1), .O(N193));
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );

  xor2  gate231(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate232(.a(gate51inter0), .b(s_10), .O(gate51inter1));
  and2  gate233(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate234(.a(s_10), .O(gate51inter3));
  inv1  gate235(.a(s_11), .O(gate51inter4));
  nand2 gate236(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate237(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate238(.a(N203), .O(gate51inter7));
  inv1  gate239(.a(N159), .O(gate51inter8));
  nand2 gate240(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate241(.a(s_11), .b(gate51inter3), .O(gate51inter10));
  nor2  gate242(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate243(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate244(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );

  xor2  gate301(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate302(.a(gate53inter0), .b(s_20), .O(gate53inter1));
  and2  gate303(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate304(.a(s_20), .O(gate53inter3));
  inv1  gate305(.a(s_21), .O(gate53inter4));
  nand2 gate306(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate307(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate308(.a(N203), .O(gate53inter7));
  inv1  gate309(.a(N165), .O(gate53inter8));
  nand2 gate310(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate311(.a(s_21), .b(gate53inter3), .O(gate53inter10));
  nor2  gate312(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate313(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate314(.a(gate53inter12), .b(gate53inter1), .O(N233));
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );

  xor2  gate189(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate190(.a(gate56inter0), .b(s_4), .O(gate56inter1));
  and2  gate191(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate192(.a(s_4), .O(gate56inter3));
  inv1  gate193(.a(s_5), .O(gate56inter4));
  nand2 gate194(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate195(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate196(.a(N1), .O(gate56inter7));
  inv1  gate197(.a(N213), .O(gate56inter8));
  nand2 gate198(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate199(.a(s_5), .b(gate56inter3), .O(gate56inter10));
  nor2  gate200(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate201(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate202(.a(gate56inter12), .b(gate56inter1), .O(N242));

  xor2  gate175(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate176(.a(gate57inter0), .b(s_2), .O(gate57inter1));
  and2  gate177(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate178(.a(s_2), .O(gate57inter3));
  inv1  gate179(.a(s_3), .O(gate57inter4));
  nand2 gate180(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate181(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate182(.a(N203), .O(gate57inter7));
  inv1  gate183(.a(N174), .O(gate57inter8));
  nand2 gate184(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate185(.a(s_3), .b(gate57inter3), .O(gate57inter10));
  nor2  gate186(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate187(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate188(.a(gate57inter12), .b(gate57inter1), .O(N243));
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );

  xor2  gate287(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate288(.a(gate76inter0), .b(s_18), .O(gate76inter1));
  and2  gate289(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate290(.a(s_18), .O(gate76inter3));
  inv1  gate291(.a(s_19), .O(gate76inter4));
  nand2 gate292(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate293(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate294(.a(N247), .O(gate76inter7));
  inv1  gate295(.a(N195), .O(gate76inter8));
  nand2 gate296(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate297(.a(s_19), .b(gate76inter3), .O(gate76inter10));
  nor2  gate298(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate299(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate300(.a(gate76inter12), .b(gate76inter1), .O(N282));
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );

  xor2  gate343(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate344(.a(gate84inter0), .b(s_26), .O(gate84inter1));
  and2  gate345(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate346(.a(s_26), .O(gate84inter3));
  inv1  gate347(.a(s_27), .O(gate84inter4));
  nand2 gate348(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate349(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate350(.a(N247), .O(gate84inter7));
  inv1  gate351(.a(N196), .O(gate84inter8));
  nand2 gate352(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate353(.a(s_27), .b(gate84inter3), .O(gate84inter10));
  nor2  gate354(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate355(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate356(.a(gate84inter12), .b(gate84inter1), .O(N294));
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate245(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate246(.a(gate105inter0), .b(s_12), .O(gate105inter1));
  and2  gate247(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate248(.a(s_12), .O(gate105inter3));
  inv1  gate249(.a(s_13), .O(gate105inter4));
  nand2 gate250(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate251(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate252(.a(N319), .O(gate105inter7));
  inv1  gate253(.a(N21), .O(gate105inter8));
  nand2 gate254(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate255(.a(s_13), .b(gate105inter3), .O(gate105inter10));
  nor2  gate256(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate257(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate258(.a(gate105inter12), .b(gate105inter1), .O(N336));
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate357(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate358(.a(gate115inter0), .b(s_28), .O(gate115inter1));
  and2  gate359(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate360(.a(s_28), .O(gate115inter3));
  inv1  gate361(.a(s_29), .O(gate115inter4));
  nand2 gate362(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate363(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate364(.a(N319), .O(gate115inter7));
  inv1  gate365(.a(N99), .O(gate115inter8));
  nand2 gate366(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate367(.a(s_29), .b(gate115inter3), .O(gate115inter10));
  nor2  gate368(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate369(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate370(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );

  xor2  gate315(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate316(.a(gate124inter0), .b(s_22), .O(gate124inter1));
  and2  gate317(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate318(.a(s_22), .O(gate124inter3));
  inv1  gate319(.a(s_23), .O(gate124inter4));
  nand2 gate320(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate321(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate322(.a(N341), .O(gate124inter7));
  inv1  gate323(.a(N307), .O(gate124inter8));
  nand2 gate324(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate325(.a(s_23), .b(gate124inter3), .O(gate124inter10));
  nor2  gate326(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate327(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate328(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate161(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate162(.a(gate132inter0), .b(s_0), .O(gate132inter1));
  and2  gate163(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate164(.a(s_0), .O(gate132inter3));
  inv1  gate165(.a(s_1), .O(gate132inter4));
  nand2 gate166(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate167(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate168(.a(N360), .O(gate132inter7));
  inv1  gate169(.a(N53), .O(gate132inter8));
  nand2 gate170(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate171(.a(s_1), .b(gate132inter3), .O(gate132inter10));
  nor2  gate172(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate173(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate174(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule