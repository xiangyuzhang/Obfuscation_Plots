module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate785(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate786(.a(gate9inter0), .b(s_34), .O(gate9inter1));
  and2  gate787(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate788(.a(s_34), .O(gate9inter3));
  inv1  gate789(.a(s_35), .O(gate9inter4));
  nand2 gate790(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate791(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate792(.a(G1), .O(gate9inter7));
  inv1  gate793(.a(G2), .O(gate9inter8));
  nand2 gate794(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate795(.a(s_35), .b(gate9inter3), .O(gate9inter10));
  nor2  gate796(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate797(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate798(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2283(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2284(.a(gate14inter0), .b(s_248), .O(gate14inter1));
  and2  gate2285(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2286(.a(s_248), .O(gate14inter3));
  inv1  gate2287(.a(s_249), .O(gate14inter4));
  nand2 gate2288(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2289(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2290(.a(G11), .O(gate14inter7));
  inv1  gate2291(.a(G12), .O(gate14inter8));
  nand2 gate2292(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2293(.a(s_249), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2294(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2295(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2296(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate687(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate688(.a(gate16inter0), .b(s_20), .O(gate16inter1));
  and2  gate689(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate690(.a(s_20), .O(gate16inter3));
  inv1  gate691(.a(s_21), .O(gate16inter4));
  nand2 gate692(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate693(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate694(.a(G15), .O(gate16inter7));
  inv1  gate695(.a(G16), .O(gate16inter8));
  nand2 gate696(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate697(.a(s_21), .b(gate16inter3), .O(gate16inter10));
  nor2  gate698(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate699(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate700(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1163(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1164(.a(gate17inter0), .b(s_88), .O(gate17inter1));
  and2  gate1165(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1166(.a(s_88), .O(gate17inter3));
  inv1  gate1167(.a(s_89), .O(gate17inter4));
  nand2 gate1168(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1169(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1170(.a(G17), .O(gate17inter7));
  inv1  gate1171(.a(G18), .O(gate17inter8));
  nand2 gate1172(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1173(.a(s_89), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1174(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1175(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1176(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1191(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1192(.a(gate18inter0), .b(s_92), .O(gate18inter1));
  and2  gate1193(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1194(.a(s_92), .O(gate18inter3));
  inv1  gate1195(.a(s_93), .O(gate18inter4));
  nand2 gate1196(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1197(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1198(.a(G19), .O(gate18inter7));
  inv1  gate1199(.a(G20), .O(gate18inter8));
  nand2 gate1200(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1201(.a(s_93), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1202(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1203(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1204(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate939(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate940(.a(gate19inter0), .b(s_56), .O(gate19inter1));
  and2  gate941(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate942(.a(s_56), .O(gate19inter3));
  inv1  gate943(.a(s_57), .O(gate19inter4));
  nand2 gate944(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate945(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate946(.a(G21), .O(gate19inter7));
  inv1  gate947(.a(G22), .O(gate19inter8));
  nand2 gate948(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate949(.a(s_57), .b(gate19inter3), .O(gate19inter10));
  nor2  gate950(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate951(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate952(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1219(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1220(.a(gate21inter0), .b(s_96), .O(gate21inter1));
  and2  gate1221(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1222(.a(s_96), .O(gate21inter3));
  inv1  gate1223(.a(s_97), .O(gate21inter4));
  nand2 gate1224(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1225(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1226(.a(G25), .O(gate21inter7));
  inv1  gate1227(.a(G26), .O(gate21inter8));
  nand2 gate1228(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1229(.a(s_97), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1230(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1231(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1232(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate617(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate618(.a(gate23inter0), .b(s_10), .O(gate23inter1));
  and2  gate619(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate620(.a(s_10), .O(gate23inter3));
  inv1  gate621(.a(s_11), .O(gate23inter4));
  nand2 gate622(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate623(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate624(.a(G29), .O(gate23inter7));
  inv1  gate625(.a(G30), .O(gate23inter8));
  nand2 gate626(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate627(.a(s_11), .b(gate23inter3), .O(gate23inter10));
  nor2  gate628(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate629(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate630(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1415(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1416(.a(gate24inter0), .b(s_124), .O(gate24inter1));
  and2  gate1417(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1418(.a(s_124), .O(gate24inter3));
  inv1  gate1419(.a(s_125), .O(gate24inter4));
  nand2 gate1420(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1421(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1422(.a(G31), .O(gate24inter7));
  inv1  gate1423(.a(G32), .O(gate24inter8));
  nand2 gate1424(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1425(.a(s_125), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1426(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1427(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1428(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2325(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2326(.a(gate28inter0), .b(s_254), .O(gate28inter1));
  and2  gate2327(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2328(.a(s_254), .O(gate28inter3));
  inv1  gate2329(.a(s_255), .O(gate28inter4));
  nand2 gate2330(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2331(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2332(.a(G10), .O(gate28inter7));
  inv1  gate2333(.a(G14), .O(gate28inter8));
  nand2 gate2334(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2335(.a(s_255), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2336(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2337(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2338(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1737(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1738(.a(gate29inter0), .b(s_170), .O(gate29inter1));
  and2  gate1739(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1740(.a(s_170), .O(gate29inter3));
  inv1  gate1741(.a(s_171), .O(gate29inter4));
  nand2 gate1742(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1743(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1744(.a(G3), .O(gate29inter7));
  inv1  gate1745(.a(G7), .O(gate29inter8));
  nand2 gate1746(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1747(.a(s_171), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1748(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1749(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1750(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2675(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2676(.a(gate38inter0), .b(s_304), .O(gate38inter1));
  and2  gate2677(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2678(.a(s_304), .O(gate38inter3));
  inv1  gate2679(.a(s_305), .O(gate38inter4));
  nand2 gate2680(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2681(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2682(.a(G27), .O(gate38inter7));
  inv1  gate2683(.a(G31), .O(gate38inter8));
  nand2 gate2684(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2685(.a(s_305), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2686(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2687(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2688(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1779(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1780(.a(gate39inter0), .b(s_176), .O(gate39inter1));
  and2  gate1781(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1782(.a(s_176), .O(gate39inter3));
  inv1  gate1783(.a(s_177), .O(gate39inter4));
  nand2 gate1784(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1785(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1786(.a(G20), .O(gate39inter7));
  inv1  gate1787(.a(G24), .O(gate39inter8));
  nand2 gate1788(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1789(.a(s_177), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1790(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1791(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1792(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2465(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2466(.a(gate41inter0), .b(s_274), .O(gate41inter1));
  and2  gate2467(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2468(.a(s_274), .O(gate41inter3));
  inv1  gate2469(.a(s_275), .O(gate41inter4));
  nand2 gate2470(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2471(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2472(.a(G1), .O(gate41inter7));
  inv1  gate2473(.a(G266), .O(gate41inter8));
  nand2 gate2474(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2475(.a(s_275), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2476(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2477(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2478(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1569(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1570(.a(gate42inter0), .b(s_146), .O(gate42inter1));
  and2  gate1571(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1572(.a(s_146), .O(gate42inter3));
  inv1  gate1573(.a(s_147), .O(gate42inter4));
  nand2 gate1574(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1575(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1576(.a(G2), .O(gate42inter7));
  inv1  gate1577(.a(G266), .O(gate42inter8));
  nand2 gate1578(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1579(.a(s_147), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1580(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1581(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1582(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate3053(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate3054(.a(gate43inter0), .b(s_358), .O(gate43inter1));
  and2  gate3055(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate3056(.a(s_358), .O(gate43inter3));
  inv1  gate3057(.a(s_359), .O(gate43inter4));
  nand2 gate3058(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate3059(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate3060(.a(G3), .O(gate43inter7));
  inv1  gate3061(.a(G269), .O(gate43inter8));
  nand2 gate3062(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate3063(.a(s_359), .b(gate43inter3), .O(gate43inter10));
  nor2  gate3064(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate3065(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate3066(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1023(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1024(.a(gate44inter0), .b(s_68), .O(gate44inter1));
  and2  gate1025(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1026(.a(s_68), .O(gate44inter3));
  inv1  gate1027(.a(s_69), .O(gate44inter4));
  nand2 gate1028(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1029(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1030(.a(G4), .O(gate44inter7));
  inv1  gate1031(.a(G269), .O(gate44inter8));
  nand2 gate1032(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1033(.a(s_69), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1034(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1035(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1036(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate897(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate898(.a(gate47inter0), .b(s_50), .O(gate47inter1));
  and2  gate899(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate900(.a(s_50), .O(gate47inter3));
  inv1  gate901(.a(s_51), .O(gate47inter4));
  nand2 gate902(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate903(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate904(.a(G7), .O(gate47inter7));
  inv1  gate905(.a(G275), .O(gate47inter8));
  nand2 gate906(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate907(.a(s_51), .b(gate47inter3), .O(gate47inter10));
  nor2  gate908(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate909(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate910(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2647(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2648(.a(gate49inter0), .b(s_300), .O(gate49inter1));
  and2  gate2649(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2650(.a(s_300), .O(gate49inter3));
  inv1  gate2651(.a(s_301), .O(gate49inter4));
  nand2 gate2652(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2653(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2654(.a(G9), .O(gate49inter7));
  inv1  gate2655(.a(G278), .O(gate49inter8));
  nand2 gate2656(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2657(.a(s_301), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2658(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2659(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2660(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1527(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1528(.a(gate55inter0), .b(s_140), .O(gate55inter1));
  and2  gate1529(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1530(.a(s_140), .O(gate55inter3));
  inv1  gate1531(.a(s_141), .O(gate55inter4));
  nand2 gate1532(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1533(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1534(.a(G15), .O(gate55inter7));
  inv1  gate1535(.a(G287), .O(gate55inter8));
  nand2 gate1536(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1537(.a(s_141), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1538(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1539(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1540(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1331(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1332(.a(gate60inter0), .b(s_112), .O(gate60inter1));
  and2  gate1333(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1334(.a(s_112), .O(gate60inter3));
  inv1  gate1335(.a(s_113), .O(gate60inter4));
  nand2 gate1336(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1337(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1338(.a(G20), .O(gate60inter7));
  inv1  gate1339(.a(G293), .O(gate60inter8));
  nand2 gate1340(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1341(.a(s_113), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1342(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1343(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1344(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1149(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1150(.a(gate61inter0), .b(s_86), .O(gate61inter1));
  and2  gate1151(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1152(.a(s_86), .O(gate61inter3));
  inv1  gate1153(.a(s_87), .O(gate61inter4));
  nand2 gate1154(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1155(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1156(.a(G21), .O(gate61inter7));
  inv1  gate1157(.a(G296), .O(gate61inter8));
  nand2 gate1158(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1159(.a(s_87), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1160(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1161(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1162(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1429(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1430(.a(gate64inter0), .b(s_126), .O(gate64inter1));
  and2  gate1431(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1432(.a(s_126), .O(gate64inter3));
  inv1  gate1433(.a(s_127), .O(gate64inter4));
  nand2 gate1434(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1435(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1436(.a(G24), .O(gate64inter7));
  inv1  gate1437(.a(G299), .O(gate64inter8));
  nand2 gate1438(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1439(.a(s_127), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1440(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1441(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1442(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1821(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1822(.a(gate65inter0), .b(s_182), .O(gate65inter1));
  and2  gate1823(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1824(.a(s_182), .O(gate65inter3));
  inv1  gate1825(.a(s_183), .O(gate65inter4));
  nand2 gate1826(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1827(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1828(.a(G25), .O(gate65inter7));
  inv1  gate1829(.a(G302), .O(gate65inter8));
  nand2 gate1830(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1831(.a(s_183), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1832(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1833(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1834(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1177(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1178(.a(gate68inter0), .b(s_90), .O(gate68inter1));
  and2  gate1179(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1180(.a(s_90), .O(gate68inter3));
  inv1  gate1181(.a(s_91), .O(gate68inter4));
  nand2 gate1182(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1183(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1184(.a(G28), .O(gate68inter7));
  inv1  gate1185(.a(G305), .O(gate68inter8));
  nand2 gate1186(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1187(.a(s_91), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1188(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1189(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1190(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate1891(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1892(.a(gate69inter0), .b(s_192), .O(gate69inter1));
  and2  gate1893(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1894(.a(s_192), .O(gate69inter3));
  inv1  gate1895(.a(s_193), .O(gate69inter4));
  nand2 gate1896(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1897(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1898(.a(G29), .O(gate69inter7));
  inv1  gate1899(.a(G308), .O(gate69inter8));
  nand2 gate1900(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1901(.a(s_193), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1902(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1903(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1904(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2367(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2368(.a(gate72inter0), .b(s_260), .O(gate72inter1));
  and2  gate2369(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2370(.a(s_260), .O(gate72inter3));
  inv1  gate2371(.a(s_261), .O(gate72inter4));
  nand2 gate2372(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2373(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2374(.a(G32), .O(gate72inter7));
  inv1  gate2375(.a(G311), .O(gate72inter8));
  nand2 gate2376(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2377(.a(s_261), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2378(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2379(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2380(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2297(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2298(.a(gate76inter0), .b(s_250), .O(gate76inter1));
  and2  gate2299(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2300(.a(s_250), .O(gate76inter3));
  inv1  gate2301(.a(s_251), .O(gate76inter4));
  nand2 gate2302(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2303(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2304(.a(G13), .O(gate76inter7));
  inv1  gate2305(.a(G317), .O(gate76inter8));
  nand2 gate2306(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2307(.a(s_251), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2308(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2309(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2310(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1457(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1458(.a(gate77inter0), .b(s_130), .O(gate77inter1));
  and2  gate1459(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1460(.a(s_130), .O(gate77inter3));
  inv1  gate1461(.a(s_131), .O(gate77inter4));
  nand2 gate1462(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1463(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1464(.a(G2), .O(gate77inter7));
  inv1  gate1465(.a(G320), .O(gate77inter8));
  nand2 gate1466(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1467(.a(s_131), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1468(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1469(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1470(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1625(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1626(.a(gate84inter0), .b(s_154), .O(gate84inter1));
  and2  gate1627(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1628(.a(s_154), .O(gate84inter3));
  inv1  gate1629(.a(s_155), .O(gate84inter4));
  nand2 gate1630(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1631(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1632(.a(G15), .O(gate84inter7));
  inv1  gate1633(.a(G329), .O(gate84inter8));
  nand2 gate1634(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1635(.a(s_155), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1636(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1637(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1638(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1653(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1654(.a(gate85inter0), .b(s_158), .O(gate85inter1));
  and2  gate1655(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1656(.a(s_158), .O(gate85inter3));
  inv1  gate1657(.a(s_159), .O(gate85inter4));
  nand2 gate1658(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1659(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1660(.a(G4), .O(gate85inter7));
  inv1  gate1661(.a(G332), .O(gate85inter8));
  nand2 gate1662(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1663(.a(s_159), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1664(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1665(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1666(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate2815(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2816(.a(gate86inter0), .b(s_324), .O(gate86inter1));
  and2  gate2817(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2818(.a(s_324), .O(gate86inter3));
  inv1  gate2819(.a(s_325), .O(gate86inter4));
  nand2 gate2820(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2821(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2822(.a(G8), .O(gate86inter7));
  inv1  gate2823(.a(G332), .O(gate86inter8));
  nand2 gate2824(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2825(.a(s_325), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2826(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2827(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2828(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1765(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1766(.a(gate87inter0), .b(s_174), .O(gate87inter1));
  and2  gate1767(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1768(.a(s_174), .O(gate87inter3));
  inv1  gate1769(.a(s_175), .O(gate87inter4));
  nand2 gate1770(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1771(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1772(.a(G12), .O(gate87inter7));
  inv1  gate1773(.a(G335), .O(gate87inter8));
  nand2 gate1774(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1775(.a(s_175), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1776(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1777(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1778(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2073(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2074(.a(gate90inter0), .b(s_218), .O(gate90inter1));
  and2  gate2075(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2076(.a(s_218), .O(gate90inter3));
  inv1  gate2077(.a(s_219), .O(gate90inter4));
  nand2 gate2078(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2079(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2080(.a(G21), .O(gate90inter7));
  inv1  gate2081(.a(G338), .O(gate90inter8));
  nand2 gate2082(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2083(.a(s_219), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2084(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2085(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2086(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate673(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate674(.a(gate94inter0), .b(s_18), .O(gate94inter1));
  and2  gate675(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate676(.a(s_18), .O(gate94inter3));
  inv1  gate677(.a(s_19), .O(gate94inter4));
  nand2 gate678(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate679(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate680(.a(G22), .O(gate94inter7));
  inv1  gate681(.a(G344), .O(gate94inter8));
  nand2 gate682(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate683(.a(s_19), .b(gate94inter3), .O(gate94inter10));
  nor2  gate684(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate685(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate686(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2969(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2970(.a(gate96inter0), .b(s_346), .O(gate96inter1));
  and2  gate2971(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2972(.a(s_346), .O(gate96inter3));
  inv1  gate2973(.a(s_347), .O(gate96inter4));
  nand2 gate2974(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2975(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2976(.a(G30), .O(gate96inter7));
  inv1  gate2977(.a(G347), .O(gate96inter8));
  nand2 gate2978(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2979(.a(s_347), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2980(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2981(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2982(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate659(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate660(.a(gate97inter0), .b(s_16), .O(gate97inter1));
  and2  gate661(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate662(.a(s_16), .O(gate97inter3));
  inv1  gate663(.a(s_17), .O(gate97inter4));
  nand2 gate664(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate665(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate666(.a(G19), .O(gate97inter7));
  inv1  gate667(.a(G350), .O(gate97inter8));
  nand2 gate668(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate669(.a(s_17), .b(gate97inter3), .O(gate97inter10));
  nor2  gate670(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate671(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate672(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1499(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1500(.a(gate98inter0), .b(s_136), .O(gate98inter1));
  and2  gate1501(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1502(.a(s_136), .O(gate98inter3));
  inv1  gate1503(.a(s_137), .O(gate98inter4));
  nand2 gate1504(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1505(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1506(.a(G23), .O(gate98inter7));
  inv1  gate1507(.a(G350), .O(gate98inter8));
  nand2 gate1508(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1509(.a(s_137), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1510(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1511(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1512(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate2899(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2900(.a(gate99inter0), .b(s_336), .O(gate99inter1));
  and2  gate2901(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2902(.a(s_336), .O(gate99inter3));
  inv1  gate2903(.a(s_337), .O(gate99inter4));
  nand2 gate2904(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2905(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2906(.a(G27), .O(gate99inter7));
  inv1  gate2907(.a(G353), .O(gate99inter8));
  nand2 gate2908(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2909(.a(s_337), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2910(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2911(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2912(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1051(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1052(.a(gate100inter0), .b(s_72), .O(gate100inter1));
  and2  gate1053(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1054(.a(s_72), .O(gate100inter3));
  inv1  gate1055(.a(s_73), .O(gate100inter4));
  nand2 gate1056(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1057(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1058(.a(G31), .O(gate100inter7));
  inv1  gate1059(.a(G353), .O(gate100inter8));
  nand2 gate1060(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1061(.a(s_73), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1062(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1063(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1064(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1233(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1234(.a(gate102inter0), .b(s_98), .O(gate102inter1));
  and2  gate1235(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1236(.a(s_98), .O(gate102inter3));
  inv1  gate1237(.a(s_99), .O(gate102inter4));
  nand2 gate1238(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1239(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1240(.a(G24), .O(gate102inter7));
  inv1  gate1241(.a(G356), .O(gate102inter8));
  nand2 gate1242(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1243(.a(s_99), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1244(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1245(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1246(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2409(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2410(.a(gate108inter0), .b(s_266), .O(gate108inter1));
  and2  gate2411(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2412(.a(s_266), .O(gate108inter3));
  inv1  gate2413(.a(s_267), .O(gate108inter4));
  nand2 gate2414(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2415(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2416(.a(G368), .O(gate108inter7));
  inv1  gate2417(.a(G369), .O(gate108inter8));
  nand2 gate2418(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2419(.a(s_267), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2420(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2421(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2422(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate841(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate842(.a(gate110inter0), .b(s_42), .O(gate110inter1));
  and2  gate843(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate844(.a(s_42), .O(gate110inter3));
  inv1  gate845(.a(s_43), .O(gate110inter4));
  nand2 gate846(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate847(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate848(.a(G372), .O(gate110inter7));
  inv1  gate849(.a(G373), .O(gate110inter8));
  nand2 gate850(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate851(.a(s_43), .b(gate110inter3), .O(gate110inter10));
  nor2  gate852(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate853(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate854(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate799(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate800(.a(gate111inter0), .b(s_36), .O(gate111inter1));
  and2  gate801(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate802(.a(s_36), .O(gate111inter3));
  inv1  gate803(.a(s_37), .O(gate111inter4));
  nand2 gate804(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate805(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate806(.a(G374), .O(gate111inter7));
  inv1  gate807(.a(G375), .O(gate111inter8));
  nand2 gate808(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate809(.a(s_37), .b(gate111inter3), .O(gate111inter10));
  nor2  gate810(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate811(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate812(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2717(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2718(.a(gate117inter0), .b(s_310), .O(gate117inter1));
  and2  gate2719(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2720(.a(s_310), .O(gate117inter3));
  inv1  gate2721(.a(s_311), .O(gate117inter4));
  nand2 gate2722(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2723(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2724(.a(G386), .O(gate117inter7));
  inv1  gate2725(.a(G387), .O(gate117inter8));
  nand2 gate2726(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2727(.a(s_311), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2728(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2729(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2730(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate1485(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1486(.a(gate118inter0), .b(s_134), .O(gate118inter1));
  and2  gate1487(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1488(.a(s_134), .O(gate118inter3));
  inv1  gate1489(.a(s_135), .O(gate118inter4));
  nand2 gate1490(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1491(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1492(.a(G388), .O(gate118inter7));
  inv1  gate1493(.a(G389), .O(gate118inter8));
  nand2 gate1494(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1495(.a(s_135), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1496(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1497(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1498(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2983(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2984(.a(gate121inter0), .b(s_348), .O(gate121inter1));
  and2  gate2985(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2986(.a(s_348), .O(gate121inter3));
  inv1  gate2987(.a(s_349), .O(gate121inter4));
  nand2 gate2988(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2989(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2990(.a(G394), .O(gate121inter7));
  inv1  gate2991(.a(G395), .O(gate121inter8));
  nand2 gate2992(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2993(.a(s_349), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2994(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2995(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2996(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate701(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate702(.a(gate125inter0), .b(s_22), .O(gate125inter1));
  and2  gate703(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate704(.a(s_22), .O(gate125inter3));
  inv1  gate705(.a(s_23), .O(gate125inter4));
  nand2 gate706(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate707(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate708(.a(G402), .O(gate125inter7));
  inv1  gate709(.a(G403), .O(gate125inter8));
  nand2 gate710(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate711(.a(s_23), .b(gate125inter3), .O(gate125inter10));
  nor2  gate712(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate713(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate714(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate827(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate828(.a(gate127inter0), .b(s_40), .O(gate127inter1));
  and2  gate829(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate830(.a(s_40), .O(gate127inter3));
  inv1  gate831(.a(s_41), .O(gate127inter4));
  nand2 gate832(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate833(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate834(.a(G406), .O(gate127inter7));
  inv1  gate835(.a(G407), .O(gate127inter8));
  nand2 gate836(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate837(.a(s_41), .b(gate127inter3), .O(gate127inter10));
  nor2  gate838(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate839(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate840(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2017(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2018(.a(gate131inter0), .b(s_210), .O(gate131inter1));
  and2  gate2019(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2020(.a(s_210), .O(gate131inter3));
  inv1  gate2021(.a(s_211), .O(gate131inter4));
  nand2 gate2022(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2023(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2024(.a(G414), .O(gate131inter7));
  inv1  gate2025(.a(G415), .O(gate131inter8));
  nand2 gate2026(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2027(.a(s_211), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2028(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2029(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2030(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2591(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2592(.a(gate134inter0), .b(s_292), .O(gate134inter1));
  and2  gate2593(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2594(.a(s_292), .O(gate134inter3));
  inv1  gate2595(.a(s_293), .O(gate134inter4));
  nand2 gate2596(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2597(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2598(.a(G420), .O(gate134inter7));
  inv1  gate2599(.a(G421), .O(gate134inter8));
  nand2 gate2600(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2601(.a(s_293), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2602(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2603(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2604(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1345(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1346(.a(gate136inter0), .b(s_114), .O(gate136inter1));
  and2  gate1347(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1348(.a(s_114), .O(gate136inter3));
  inv1  gate1349(.a(s_115), .O(gate136inter4));
  nand2 gate1350(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1351(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1352(.a(G424), .O(gate136inter7));
  inv1  gate1353(.a(G425), .O(gate136inter8));
  nand2 gate1354(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1355(.a(s_115), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1356(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1357(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1358(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2871(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2872(.a(gate137inter0), .b(s_332), .O(gate137inter1));
  and2  gate2873(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2874(.a(s_332), .O(gate137inter3));
  inv1  gate2875(.a(s_333), .O(gate137inter4));
  nand2 gate2876(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2877(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2878(.a(G426), .O(gate137inter7));
  inv1  gate2879(.a(G429), .O(gate137inter8));
  nand2 gate2880(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2881(.a(s_333), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2882(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2883(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2884(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate911(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate912(.a(gate138inter0), .b(s_52), .O(gate138inter1));
  and2  gate913(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate914(.a(s_52), .O(gate138inter3));
  inv1  gate915(.a(s_53), .O(gate138inter4));
  nand2 gate916(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate917(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate918(.a(G432), .O(gate138inter7));
  inv1  gate919(.a(G435), .O(gate138inter8));
  nand2 gate920(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate921(.a(s_53), .b(gate138inter3), .O(gate138inter10));
  nor2  gate922(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate923(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate924(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1681(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1682(.a(gate142inter0), .b(s_162), .O(gate142inter1));
  and2  gate1683(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1684(.a(s_162), .O(gate142inter3));
  inv1  gate1685(.a(s_163), .O(gate142inter4));
  nand2 gate1686(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1687(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1688(.a(G456), .O(gate142inter7));
  inv1  gate1689(.a(G459), .O(gate142inter8));
  nand2 gate1690(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1691(.a(s_163), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1692(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1693(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1694(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1373(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1374(.a(gate144inter0), .b(s_118), .O(gate144inter1));
  and2  gate1375(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1376(.a(s_118), .O(gate144inter3));
  inv1  gate1377(.a(s_119), .O(gate144inter4));
  nand2 gate1378(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1379(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1380(.a(G468), .O(gate144inter7));
  inv1  gate1381(.a(G471), .O(gate144inter8));
  nand2 gate1382(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1383(.a(s_119), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1384(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1385(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1386(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2829(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2830(.a(gate145inter0), .b(s_326), .O(gate145inter1));
  and2  gate2831(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2832(.a(s_326), .O(gate145inter3));
  inv1  gate2833(.a(s_327), .O(gate145inter4));
  nand2 gate2834(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2835(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2836(.a(G474), .O(gate145inter7));
  inv1  gate2837(.a(G477), .O(gate145inter8));
  nand2 gate2838(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2839(.a(s_327), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2840(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2841(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2842(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate2577(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2578(.a(gate146inter0), .b(s_290), .O(gate146inter1));
  and2  gate2579(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2580(.a(s_290), .O(gate146inter3));
  inv1  gate2581(.a(s_291), .O(gate146inter4));
  nand2 gate2582(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2583(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2584(.a(G480), .O(gate146inter7));
  inv1  gate2585(.a(G483), .O(gate146inter8));
  nand2 gate2586(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2587(.a(s_291), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2588(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2589(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2590(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1541(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1542(.a(gate148inter0), .b(s_142), .O(gate148inter1));
  and2  gate1543(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1544(.a(s_142), .O(gate148inter3));
  inv1  gate1545(.a(s_143), .O(gate148inter4));
  nand2 gate1546(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1547(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1548(.a(G492), .O(gate148inter7));
  inv1  gate1549(.a(G495), .O(gate148inter8));
  nand2 gate1550(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1551(.a(s_143), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1552(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1553(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1554(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate2619(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2620(.a(gate149inter0), .b(s_296), .O(gate149inter1));
  and2  gate2621(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2622(.a(s_296), .O(gate149inter3));
  inv1  gate2623(.a(s_297), .O(gate149inter4));
  nand2 gate2624(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2625(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2626(.a(G498), .O(gate149inter7));
  inv1  gate2627(.a(G501), .O(gate149inter8));
  nand2 gate2628(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2629(.a(s_297), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2630(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2631(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2632(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2731(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2732(.a(gate152inter0), .b(s_312), .O(gate152inter1));
  and2  gate2733(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2734(.a(s_312), .O(gate152inter3));
  inv1  gate2735(.a(s_313), .O(gate152inter4));
  nand2 gate2736(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2737(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2738(.a(G516), .O(gate152inter7));
  inv1  gate2739(.a(G519), .O(gate152inter8));
  nand2 gate2740(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2741(.a(s_313), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2742(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2743(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2744(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2549(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2550(.a(gate154inter0), .b(s_286), .O(gate154inter1));
  and2  gate2551(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2552(.a(s_286), .O(gate154inter3));
  inv1  gate2553(.a(s_287), .O(gate154inter4));
  nand2 gate2554(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2555(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2556(.a(G429), .O(gate154inter7));
  inv1  gate2557(.a(G522), .O(gate154inter8));
  nand2 gate2558(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2559(.a(s_287), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2560(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2561(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2562(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1905(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1906(.a(gate155inter0), .b(s_194), .O(gate155inter1));
  and2  gate1907(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1908(.a(s_194), .O(gate155inter3));
  inv1  gate1909(.a(s_195), .O(gate155inter4));
  nand2 gate1910(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1911(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1912(.a(G432), .O(gate155inter7));
  inv1  gate1913(.a(G525), .O(gate155inter8));
  nand2 gate1914(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1915(.a(s_195), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1916(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1917(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1918(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate729(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate730(.a(gate157inter0), .b(s_26), .O(gate157inter1));
  and2  gate731(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate732(.a(s_26), .O(gate157inter3));
  inv1  gate733(.a(s_27), .O(gate157inter4));
  nand2 gate734(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate735(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate736(.a(G438), .O(gate157inter7));
  inv1  gate737(.a(G528), .O(gate157inter8));
  nand2 gate738(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate739(.a(s_27), .b(gate157inter3), .O(gate157inter10));
  nor2  gate740(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate741(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate742(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1555(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1556(.a(gate158inter0), .b(s_144), .O(gate158inter1));
  and2  gate1557(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1558(.a(s_144), .O(gate158inter3));
  inv1  gate1559(.a(s_145), .O(gate158inter4));
  nand2 gate1560(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1561(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1562(.a(G441), .O(gate158inter7));
  inv1  gate1563(.a(G528), .O(gate158inter8));
  nand2 gate1564(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1565(.a(s_145), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1566(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1567(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1568(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate3067(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate3068(.a(gate159inter0), .b(s_360), .O(gate159inter1));
  and2  gate3069(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate3070(.a(s_360), .O(gate159inter3));
  inv1  gate3071(.a(s_361), .O(gate159inter4));
  nand2 gate3072(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate3073(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate3074(.a(G444), .O(gate159inter7));
  inv1  gate3075(.a(G531), .O(gate159inter8));
  nand2 gate3076(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate3077(.a(s_361), .b(gate159inter3), .O(gate159inter10));
  nor2  gate3078(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate3079(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate3080(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2745(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2746(.a(gate161inter0), .b(s_314), .O(gate161inter1));
  and2  gate2747(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2748(.a(s_314), .O(gate161inter3));
  inv1  gate2749(.a(s_315), .O(gate161inter4));
  nand2 gate2750(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2751(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2752(.a(G450), .O(gate161inter7));
  inv1  gate2753(.a(G534), .O(gate161inter8));
  nand2 gate2754(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2755(.a(s_315), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2756(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2757(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2758(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1835(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1836(.a(gate162inter0), .b(s_184), .O(gate162inter1));
  and2  gate1837(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1838(.a(s_184), .O(gate162inter3));
  inv1  gate1839(.a(s_185), .O(gate162inter4));
  nand2 gate1840(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1841(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1842(.a(G453), .O(gate162inter7));
  inv1  gate1843(.a(G534), .O(gate162inter8));
  nand2 gate1844(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1845(.a(s_185), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1846(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1847(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1848(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate967(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate968(.a(gate169inter0), .b(s_60), .O(gate169inter1));
  and2  gate969(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate970(.a(s_60), .O(gate169inter3));
  inv1  gate971(.a(s_61), .O(gate169inter4));
  nand2 gate972(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate973(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate974(.a(G474), .O(gate169inter7));
  inv1  gate975(.a(G546), .O(gate169inter8));
  nand2 gate976(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate977(.a(s_61), .b(gate169inter3), .O(gate169inter10));
  nor2  gate978(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate979(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate980(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2339(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2340(.a(gate170inter0), .b(s_256), .O(gate170inter1));
  and2  gate2341(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2342(.a(s_256), .O(gate170inter3));
  inv1  gate2343(.a(s_257), .O(gate170inter4));
  nand2 gate2344(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2345(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2346(.a(G477), .O(gate170inter7));
  inv1  gate2347(.a(G546), .O(gate170inter8));
  nand2 gate2348(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2349(.a(s_257), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2350(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2351(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2352(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1093(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1094(.a(gate172inter0), .b(s_78), .O(gate172inter1));
  and2  gate1095(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1096(.a(s_78), .O(gate172inter3));
  inv1  gate1097(.a(s_79), .O(gate172inter4));
  nand2 gate1098(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1099(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1100(.a(G483), .O(gate172inter7));
  inv1  gate1101(.a(G549), .O(gate172inter8));
  nand2 gate1102(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1103(.a(s_79), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1104(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1105(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1106(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1135(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1136(.a(gate186inter0), .b(s_84), .O(gate186inter1));
  and2  gate1137(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1138(.a(s_84), .O(gate186inter3));
  inv1  gate1139(.a(s_85), .O(gate186inter4));
  nand2 gate1140(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1141(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1142(.a(G572), .O(gate186inter7));
  inv1  gate1143(.a(G573), .O(gate186inter8));
  nand2 gate1144(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1145(.a(s_85), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1146(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1147(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1148(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2269(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2270(.a(gate188inter0), .b(s_246), .O(gate188inter1));
  and2  gate2271(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2272(.a(s_246), .O(gate188inter3));
  inv1  gate2273(.a(s_247), .O(gate188inter4));
  nand2 gate2274(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2275(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2276(.a(G576), .O(gate188inter7));
  inv1  gate2277(.a(G577), .O(gate188inter8));
  nand2 gate2278(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2279(.a(s_247), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2280(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2281(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2282(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate589(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate590(.a(gate191inter0), .b(s_6), .O(gate191inter1));
  and2  gate591(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate592(.a(s_6), .O(gate191inter3));
  inv1  gate593(.a(s_7), .O(gate191inter4));
  nand2 gate594(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate595(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate596(.a(G582), .O(gate191inter7));
  inv1  gate597(.a(G583), .O(gate191inter8));
  nand2 gate598(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate599(.a(s_7), .b(gate191inter3), .O(gate191inter10));
  nor2  gate600(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate601(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate602(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2255(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2256(.a(gate192inter0), .b(s_244), .O(gate192inter1));
  and2  gate2257(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2258(.a(s_244), .O(gate192inter3));
  inv1  gate2259(.a(s_245), .O(gate192inter4));
  nand2 gate2260(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2261(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2262(.a(G584), .O(gate192inter7));
  inv1  gate2263(.a(G585), .O(gate192inter8));
  nand2 gate2264(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2265(.a(s_245), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2266(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2267(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2268(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1709(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1710(.a(gate196inter0), .b(s_166), .O(gate196inter1));
  and2  gate1711(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1712(.a(s_166), .O(gate196inter3));
  inv1  gate1713(.a(s_167), .O(gate196inter4));
  nand2 gate1714(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1715(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1716(.a(G592), .O(gate196inter7));
  inv1  gate1717(.a(G593), .O(gate196inter8));
  nand2 gate1718(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1719(.a(s_167), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1720(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1721(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1722(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2787(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2788(.a(gate198inter0), .b(s_320), .O(gate198inter1));
  and2  gate2789(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2790(.a(s_320), .O(gate198inter3));
  inv1  gate2791(.a(s_321), .O(gate198inter4));
  nand2 gate2792(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2793(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2794(.a(G596), .O(gate198inter7));
  inv1  gate2795(.a(G597), .O(gate198inter8));
  nand2 gate2796(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2797(.a(s_321), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2798(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2799(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2800(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2129(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2130(.a(gate200inter0), .b(s_226), .O(gate200inter1));
  and2  gate2131(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2132(.a(s_226), .O(gate200inter3));
  inv1  gate2133(.a(s_227), .O(gate200inter4));
  nand2 gate2134(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2135(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2136(.a(G600), .O(gate200inter7));
  inv1  gate2137(.a(G601), .O(gate200inter8));
  nand2 gate2138(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2139(.a(s_227), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2140(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2141(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2142(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate3011(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate3012(.a(gate203inter0), .b(s_352), .O(gate203inter1));
  and2  gate3013(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate3014(.a(s_352), .O(gate203inter3));
  inv1  gate3015(.a(s_353), .O(gate203inter4));
  nand2 gate3016(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate3017(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate3018(.a(G602), .O(gate203inter7));
  inv1  gate3019(.a(G612), .O(gate203inter8));
  nand2 gate3020(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate3021(.a(s_353), .b(gate203inter3), .O(gate203inter10));
  nor2  gate3022(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate3023(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate3024(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1317(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1318(.a(gate204inter0), .b(s_110), .O(gate204inter1));
  and2  gate1319(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1320(.a(s_110), .O(gate204inter3));
  inv1  gate1321(.a(s_111), .O(gate204inter4));
  nand2 gate1322(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1323(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1324(.a(G607), .O(gate204inter7));
  inv1  gate1325(.a(G617), .O(gate204inter8));
  nand2 gate1326(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1327(.a(s_111), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1328(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1329(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1330(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1513(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1514(.a(gate207inter0), .b(s_138), .O(gate207inter1));
  and2  gate1515(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1516(.a(s_138), .O(gate207inter3));
  inv1  gate1517(.a(s_139), .O(gate207inter4));
  nand2 gate1518(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1519(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1520(.a(G622), .O(gate207inter7));
  inv1  gate1521(.a(G632), .O(gate207inter8));
  nand2 gate1522(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1523(.a(s_139), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1524(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1525(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1526(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate995(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate996(.a(gate209inter0), .b(s_64), .O(gate209inter1));
  and2  gate997(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate998(.a(s_64), .O(gate209inter3));
  inv1  gate999(.a(s_65), .O(gate209inter4));
  nand2 gate1000(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1001(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1002(.a(G602), .O(gate209inter7));
  inv1  gate1003(.a(G666), .O(gate209inter8));
  nand2 gate1004(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1005(.a(s_65), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1006(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1007(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1008(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate603(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate604(.a(gate213inter0), .b(s_8), .O(gate213inter1));
  and2  gate605(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate606(.a(s_8), .O(gate213inter3));
  inv1  gate607(.a(s_9), .O(gate213inter4));
  nand2 gate608(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate609(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate610(.a(G602), .O(gate213inter7));
  inv1  gate611(.a(G672), .O(gate213inter8));
  nand2 gate612(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate613(.a(s_9), .b(gate213inter3), .O(gate213inter10));
  nor2  gate614(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate615(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate616(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2115(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2116(.a(gate215inter0), .b(s_224), .O(gate215inter1));
  and2  gate2117(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2118(.a(s_224), .O(gate215inter3));
  inv1  gate2119(.a(s_225), .O(gate215inter4));
  nand2 gate2120(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2121(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2122(.a(G607), .O(gate215inter7));
  inv1  gate2123(.a(G675), .O(gate215inter8));
  nand2 gate2124(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2125(.a(s_225), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2126(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2127(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2128(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2003(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2004(.a(gate218inter0), .b(s_208), .O(gate218inter1));
  and2  gate2005(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2006(.a(s_208), .O(gate218inter3));
  inv1  gate2007(.a(s_209), .O(gate218inter4));
  nand2 gate2008(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2009(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2010(.a(G627), .O(gate218inter7));
  inv1  gate2011(.a(G678), .O(gate218inter8));
  nand2 gate2012(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2013(.a(s_209), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2014(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2015(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2016(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate925(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate926(.a(gate223inter0), .b(s_54), .O(gate223inter1));
  and2  gate927(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate928(.a(s_54), .O(gate223inter3));
  inv1  gate929(.a(s_55), .O(gate223inter4));
  nand2 gate930(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate931(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate932(.a(G627), .O(gate223inter7));
  inv1  gate933(.a(G687), .O(gate223inter8));
  nand2 gate934(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate935(.a(s_55), .b(gate223inter3), .O(gate223inter10));
  nor2  gate936(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate937(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate938(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1667(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1668(.a(gate224inter0), .b(s_160), .O(gate224inter1));
  and2  gate1669(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1670(.a(s_160), .O(gate224inter3));
  inv1  gate1671(.a(s_161), .O(gate224inter4));
  nand2 gate1672(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1673(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1674(.a(G637), .O(gate224inter7));
  inv1  gate1675(.a(G687), .O(gate224inter8));
  nand2 gate1676(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1677(.a(s_161), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1678(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1679(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1680(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate2857(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2858(.a(gate225inter0), .b(s_330), .O(gate225inter1));
  and2  gate2859(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2860(.a(s_330), .O(gate225inter3));
  inv1  gate2861(.a(s_331), .O(gate225inter4));
  nand2 gate2862(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2863(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2864(.a(G690), .O(gate225inter7));
  inv1  gate2865(.a(G691), .O(gate225inter8));
  nand2 gate2866(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2867(.a(s_331), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2868(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2869(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2870(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1289(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1290(.a(gate227inter0), .b(s_106), .O(gate227inter1));
  and2  gate1291(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1292(.a(s_106), .O(gate227inter3));
  inv1  gate1293(.a(s_107), .O(gate227inter4));
  nand2 gate1294(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1295(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1296(.a(G694), .O(gate227inter7));
  inv1  gate1297(.a(G695), .O(gate227inter8));
  nand2 gate1298(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1299(.a(s_107), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1300(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1301(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1302(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2087(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2088(.a(gate229inter0), .b(s_220), .O(gate229inter1));
  and2  gate2089(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2090(.a(s_220), .O(gate229inter3));
  inv1  gate2091(.a(s_221), .O(gate229inter4));
  nand2 gate2092(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2093(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2094(.a(G698), .O(gate229inter7));
  inv1  gate2095(.a(G699), .O(gate229inter8));
  nand2 gate2096(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2097(.a(s_221), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2098(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2099(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2100(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate2395(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2396(.a(gate230inter0), .b(s_264), .O(gate230inter1));
  and2  gate2397(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2398(.a(s_264), .O(gate230inter3));
  inv1  gate2399(.a(s_265), .O(gate230inter4));
  nand2 gate2400(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2401(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2402(.a(G700), .O(gate230inter7));
  inv1  gate2403(.a(G701), .O(gate230inter8));
  nand2 gate2404(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2405(.a(s_265), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2406(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2407(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2408(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate2843(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2844(.a(gate231inter0), .b(s_328), .O(gate231inter1));
  and2  gate2845(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2846(.a(s_328), .O(gate231inter3));
  inv1  gate2847(.a(s_329), .O(gate231inter4));
  nand2 gate2848(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2849(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2850(.a(G702), .O(gate231inter7));
  inv1  gate2851(.a(G703), .O(gate231inter8));
  nand2 gate2852(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2853(.a(s_329), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2854(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2855(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2856(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1037(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1038(.a(gate233inter0), .b(s_70), .O(gate233inter1));
  and2  gate1039(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1040(.a(s_70), .O(gate233inter3));
  inv1  gate1041(.a(s_71), .O(gate233inter4));
  nand2 gate1042(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1043(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1044(.a(G242), .O(gate233inter7));
  inv1  gate1045(.a(G718), .O(gate233inter8));
  nand2 gate1046(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1047(.a(s_71), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1048(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1049(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1050(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2437(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2438(.a(gate234inter0), .b(s_270), .O(gate234inter1));
  and2  gate2439(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2440(.a(s_270), .O(gate234inter3));
  inv1  gate2441(.a(s_271), .O(gate234inter4));
  nand2 gate2442(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2443(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2444(.a(G245), .O(gate234inter7));
  inv1  gate2445(.a(G721), .O(gate234inter8));
  nand2 gate2446(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2447(.a(s_271), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2448(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2449(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2450(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2941(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2942(.a(gate235inter0), .b(s_342), .O(gate235inter1));
  and2  gate2943(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2944(.a(s_342), .O(gate235inter3));
  inv1  gate2945(.a(s_343), .O(gate235inter4));
  nand2 gate2946(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2947(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2948(.a(G248), .O(gate235inter7));
  inv1  gate2949(.a(G724), .O(gate235inter8));
  nand2 gate2950(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2951(.a(s_343), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2952(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2953(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2954(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate2955(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2956(.a(gate242inter0), .b(s_344), .O(gate242inter1));
  and2  gate2957(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2958(.a(s_344), .O(gate242inter3));
  inv1  gate2959(.a(s_345), .O(gate242inter4));
  nand2 gate2960(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2961(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2962(.a(G718), .O(gate242inter7));
  inv1  gate2963(.a(G730), .O(gate242inter8));
  nand2 gate2964(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2965(.a(s_345), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2966(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2967(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2968(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2479(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2480(.a(gate244inter0), .b(s_276), .O(gate244inter1));
  and2  gate2481(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2482(.a(s_276), .O(gate244inter3));
  inv1  gate2483(.a(s_277), .O(gate244inter4));
  nand2 gate2484(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2485(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2486(.a(G721), .O(gate244inter7));
  inv1  gate2487(.a(G733), .O(gate244inter8));
  nand2 gate2488(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2489(.a(s_277), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2490(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2491(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2492(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2171(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2172(.a(gate246inter0), .b(s_232), .O(gate246inter1));
  and2  gate2173(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2174(.a(s_232), .O(gate246inter3));
  inv1  gate2175(.a(s_233), .O(gate246inter4));
  nand2 gate2176(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2177(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2178(.a(G724), .O(gate246inter7));
  inv1  gate2179(.a(G736), .O(gate246inter8));
  nand2 gate2180(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2181(.a(s_233), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2182(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2183(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2184(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate2199(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate2200(.a(gate247inter0), .b(s_236), .O(gate247inter1));
  and2  gate2201(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate2202(.a(s_236), .O(gate247inter3));
  inv1  gate2203(.a(s_237), .O(gate247inter4));
  nand2 gate2204(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate2205(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate2206(.a(G251), .O(gate247inter7));
  inv1  gate2207(.a(G739), .O(gate247inter8));
  nand2 gate2208(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate2209(.a(s_237), .b(gate247inter3), .O(gate247inter10));
  nor2  gate2210(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate2211(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate2212(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1989(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1990(.a(gate249inter0), .b(s_206), .O(gate249inter1));
  and2  gate1991(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1992(.a(s_206), .O(gate249inter3));
  inv1  gate1993(.a(s_207), .O(gate249inter4));
  nand2 gate1994(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1995(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1996(.a(G254), .O(gate249inter7));
  inv1  gate1997(.a(G742), .O(gate249inter8));
  nand2 gate1998(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1999(.a(s_207), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2000(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2001(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2002(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1597(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1598(.a(gate253inter0), .b(s_150), .O(gate253inter1));
  and2  gate1599(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1600(.a(s_150), .O(gate253inter3));
  inv1  gate1601(.a(s_151), .O(gate253inter4));
  nand2 gate1602(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1603(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1604(.a(G260), .O(gate253inter7));
  inv1  gate1605(.a(G748), .O(gate253inter8));
  nand2 gate1606(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1607(.a(s_151), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1608(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1609(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1610(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2311(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2312(.a(gate256inter0), .b(s_252), .O(gate256inter1));
  and2  gate2313(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2314(.a(s_252), .O(gate256inter3));
  inv1  gate2315(.a(s_253), .O(gate256inter4));
  nand2 gate2316(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2317(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2318(.a(G715), .O(gate256inter7));
  inv1  gate2319(.a(G751), .O(gate256inter8));
  nand2 gate2320(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2321(.a(s_253), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2322(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2323(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2324(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate869(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate870(.a(gate257inter0), .b(s_46), .O(gate257inter1));
  and2  gate871(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate872(.a(s_46), .O(gate257inter3));
  inv1  gate873(.a(s_47), .O(gate257inter4));
  nand2 gate874(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate875(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate876(.a(G754), .O(gate257inter7));
  inv1  gate877(.a(G755), .O(gate257inter8));
  nand2 gate878(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate879(.a(s_47), .b(gate257inter3), .O(gate257inter10));
  nor2  gate880(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate881(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate882(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1261(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1262(.a(gate259inter0), .b(s_102), .O(gate259inter1));
  and2  gate1263(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1264(.a(s_102), .O(gate259inter3));
  inv1  gate1265(.a(s_103), .O(gate259inter4));
  nand2 gate1266(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1267(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1268(.a(G758), .O(gate259inter7));
  inv1  gate1269(.a(G759), .O(gate259inter8));
  nand2 gate1270(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1271(.a(s_103), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1272(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1273(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1274(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2885(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2886(.a(gate261inter0), .b(s_334), .O(gate261inter1));
  and2  gate2887(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2888(.a(s_334), .O(gate261inter3));
  inv1  gate2889(.a(s_335), .O(gate261inter4));
  nand2 gate2890(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2891(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2892(.a(G762), .O(gate261inter7));
  inv1  gate2893(.a(G763), .O(gate261inter8));
  nand2 gate2894(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2895(.a(s_335), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2896(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2897(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2898(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1107(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1108(.a(gate262inter0), .b(s_80), .O(gate262inter1));
  and2  gate1109(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1110(.a(s_80), .O(gate262inter3));
  inv1  gate1111(.a(s_81), .O(gate262inter4));
  nand2 gate1112(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1113(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1114(.a(G764), .O(gate262inter7));
  inv1  gate1115(.a(G765), .O(gate262inter8));
  nand2 gate1116(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1117(.a(s_81), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1118(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1119(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1120(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate645(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate646(.a(gate263inter0), .b(s_14), .O(gate263inter1));
  and2  gate647(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate648(.a(s_14), .O(gate263inter3));
  inv1  gate649(.a(s_15), .O(gate263inter4));
  nand2 gate650(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate651(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate652(.a(G766), .O(gate263inter7));
  inv1  gate653(.a(G767), .O(gate263inter8));
  nand2 gate654(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate655(.a(s_15), .b(gate263inter3), .O(gate263inter10));
  nor2  gate656(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate657(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate658(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1275(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1276(.a(gate264inter0), .b(s_104), .O(gate264inter1));
  and2  gate1277(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1278(.a(s_104), .O(gate264inter3));
  inv1  gate1279(.a(s_105), .O(gate264inter4));
  nand2 gate1280(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1281(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1282(.a(G768), .O(gate264inter7));
  inv1  gate1283(.a(G769), .O(gate264inter8));
  nand2 gate1284(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1285(.a(s_105), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1286(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1287(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1288(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate771(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate772(.a(gate265inter0), .b(s_32), .O(gate265inter1));
  and2  gate773(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate774(.a(s_32), .O(gate265inter3));
  inv1  gate775(.a(s_33), .O(gate265inter4));
  nand2 gate776(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate777(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate778(.a(G642), .O(gate265inter7));
  inv1  gate779(.a(G770), .O(gate265inter8));
  nand2 gate780(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate781(.a(s_33), .b(gate265inter3), .O(gate265inter10));
  nor2  gate782(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate783(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate784(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2353(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2354(.a(gate267inter0), .b(s_258), .O(gate267inter1));
  and2  gate2355(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2356(.a(s_258), .O(gate267inter3));
  inv1  gate2357(.a(s_259), .O(gate267inter4));
  nand2 gate2358(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2359(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2360(.a(G648), .O(gate267inter7));
  inv1  gate2361(.a(G776), .O(gate267inter8));
  nand2 gate2362(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2363(.a(s_259), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2364(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2365(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2366(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1065(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1066(.a(gate272inter0), .b(s_74), .O(gate272inter1));
  and2  gate1067(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1068(.a(s_74), .O(gate272inter3));
  inv1  gate1069(.a(s_75), .O(gate272inter4));
  nand2 gate1070(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1071(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1072(.a(G663), .O(gate272inter7));
  inv1  gate1073(.a(G791), .O(gate272inter8));
  nand2 gate1074(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1075(.a(s_75), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1076(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1077(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1078(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1793(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1794(.a(gate275inter0), .b(s_178), .O(gate275inter1));
  and2  gate1795(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1796(.a(s_178), .O(gate275inter3));
  inv1  gate1797(.a(s_179), .O(gate275inter4));
  nand2 gate1798(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1799(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1800(.a(G645), .O(gate275inter7));
  inv1  gate1801(.a(G797), .O(gate275inter8));
  nand2 gate1802(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1803(.a(s_179), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1804(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1805(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1806(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate953(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate954(.a(gate278inter0), .b(s_58), .O(gate278inter1));
  and2  gate955(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate956(.a(s_58), .O(gate278inter3));
  inv1  gate957(.a(s_59), .O(gate278inter4));
  nand2 gate958(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate959(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate960(.a(G776), .O(gate278inter7));
  inv1  gate961(.a(G800), .O(gate278inter8));
  nand2 gate962(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate963(.a(s_59), .b(gate278inter3), .O(gate278inter10));
  nor2  gate964(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate965(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate966(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1079(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1080(.a(gate280inter0), .b(s_76), .O(gate280inter1));
  and2  gate1081(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1082(.a(s_76), .O(gate280inter3));
  inv1  gate1083(.a(s_77), .O(gate280inter4));
  nand2 gate1084(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1085(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1086(.a(G779), .O(gate280inter7));
  inv1  gate1087(.a(G803), .O(gate280inter8));
  nand2 gate1088(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1089(.a(s_77), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1090(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1091(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1092(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate631(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate632(.a(gate281inter0), .b(s_12), .O(gate281inter1));
  and2  gate633(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate634(.a(s_12), .O(gate281inter3));
  inv1  gate635(.a(s_13), .O(gate281inter4));
  nand2 gate636(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate637(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate638(.a(G654), .O(gate281inter7));
  inv1  gate639(.a(G806), .O(gate281inter8));
  nand2 gate640(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate641(.a(s_13), .b(gate281inter3), .O(gate281inter10));
  nor2  gate642(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate643(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate644(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2535(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2536(.a(gate285inter0), .b(s_284), .O(gate285inter1));
  and2  gate2537(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2538(.a(s_284), .O(gate285inter3));
  inv1  gate2539(.a(s_285), .O(gate285inter4));
  nand2 gate2540(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2541(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2542(.a(G660), .O(gate285inter7));
  inv1  gate2543(.a(G812), .O(gate285inter8));
  nand2 gate2544(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2545(.a(s_285), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2546(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2547(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2548(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2927(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2928(.a(gate288inter0), .b(s_340), .O(gate288inter1));
  and2  gate2929(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2930(.a(s_340), .O(gate288inter3));
  inv1  gate2931(.a(s_341), .O(gate288inter4));
  nand2 gate2932(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2933(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2934(.a(G791), .O(gate288inter7));
  inv1  gate2935(.a(G815), .O(gate288inter8));
  nand2 gate2936(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2937(.a(s_341), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2938(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2939(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2940(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate855(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate856(.a(gate291inter0), .b(s_44), .O(gate291inter1));
  and2  gate857(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate858(.a(s_44), .O(gate291inter3));
  inv1  gate859(.a(s_45), .O(gate291inter4));
  nand2 gate860(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate861(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate862(.a(G822), .O(gate291inter7));
  inv1  gate863(.a(G823), .O(gate291inter8));
  nand2 gate864(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate865(.a(s_45), .b(gate291inter3), .O(gate291inter10));
  nor2  gate866(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate867(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate868(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1247(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1248(.a(gate294inter0), .b(s_100), .O(gate294inter1));
  and2  gate1249(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1250(.a(s_100), .O(gate294inter3));
  inv1  gate1251(.a(s_101), .O(gate294inter4));
  nand2 gate1252(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1253(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1254(.a(G832), .O(gate294inter7));
  inv1  gate1255(.a(G833), .O(gate294inter8));
  nand2 gate1256(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1257(.a(s_101), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1258(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1259(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1260(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1443(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1444(.a(gate296inter0), .b(s_128), .O(gate296inter1));
  and2  gate1445(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1446(.a(s_128), .O(gate296inter3));
  inv1  gate1447(.a(s_129), .O(gate296inter4));
  nand2 gate1448(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1449(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1450(.a(G826), .O(gate296inter7));
  inv1  gate1451(.a(G827), .O(gate296inter8));
  nand2 gate1452(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1453(.a(s_129), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1454(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1455(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1456(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2689(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2690(.a(gate387inter0), .b(s_306), .O(gate387inter1));
  and2  gate2691(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2692(.a(s_306), .O(gate387inter3));
  inv1  gate2693(.a(s_307), .O(gate387inter4));
  nand2 gate2694(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2695(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2696(.a(G1), .O(gate387inter7));
  inv1  gate2697(.a(G1036), .O(gate387inter8));
  nand2 gate2698(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2699(.a(s_307), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2700(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2701(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2702(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1751(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1752(.a(gate389inter0), .b(s_172), .O(gate389inter1));
  and2  gate1753(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1754(.a(s_172), .O(gate389inter3));
  inv1  gate1755(.a(s_173), .O(gate389inter4));
  nand2 gate1756(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1757(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1758(.a(G3), .O(gate389inter7));
  inv1  gate1759(.a(G1042), .O(gate389inter8));
  nand2 gate1760(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1761(.a(s_173), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1762(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1763(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1764(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate2661(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2662(.a(gate390inter0), .b(s_302), .O(gate390inter1));
  and2  gate2663(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2664(.a(s_302), .O(gate390inter3));
  inv1  gate2665(.a(s_303), .O(gate390inter4));
  nand2 gate2666(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2667(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2668(.a(G4), .O(gate390inter7));
  inv1  gate2669(.a(G1045), .O(gate390inter8));
  nand2 gate2670(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2671(.a(s_303), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2672(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2673(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2674(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate715(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate716(.a(gate391inter0), .b(s_24), .O(gate391inter1));
  and2  gate717(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate718(.a(s_24), .O(gate391inter3));
  inv1  gate719(.a(s_25), .O(gate391inter4));
  nand2 gate720(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate721(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate722(.a(G5), .O(gate391inter7));
  inv1  gate723(.a(G1048), .O(gate391inter8));
  nand2 gate724(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate725(.a(s_25), .b(gate391inter3), .O(gate391inter10));
  nor2  gate726(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate727(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate728(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1205(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1206(.a(gate392inter0), .b(s_94), .O(gate392inter1));
  and2  gate1207(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1208(.a(s_94), .O(gate392inter3));
  inv1  gate1209(.a(s_95), .O(gate392inter4));
  nand2 gate1210(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1211(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1212(.a(G6), .O(gate392inter7));
  inv1  gate1213(.a(G1051), .O(gate392inter8));
  nand2 gate1214(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1215(.a(s_95), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1216(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1217(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1218(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1933(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1934(.a(gate394inter0), .b(s_198), .O(gate394inter1));
  and2  gate1935(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1936(.a(s_198), .O(gate394inter3));
  inv1  gate1937(.a(s_199), .O(gate394inter4));
  nand2 gate1938(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1939(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1940(.a(G8), .O(gate394inter7));
  inv1  gate1941(.a(G1057), .O(gate394inter8));
  nand2 gate1942(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1943(.a(s_199), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1944(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1945(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1946(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2801(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2802(.a(gate397inter0), .b(s_322), .O(gate397inter1));
  and2  gate2803(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2804(.a(s_322), .O(gate397inter3));
  inv1  gate2805(.a(s_323), .O(gate397inter4));
  nand2 gate2806(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2807(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2808(.a(G11), .O(gate397inter7));
  inv1  gate2809(.a(G1066), .O(gate397inter8));
  nand2 gate2810(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2811(.a(s_323), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2812(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2813(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2814(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate2227(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2228(.a(gate398inter0), .b(s_240), .O(gate398inter1));
  and2  gate2229(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2230(.a(s_240), .O(gate398inter3));
  inv1  gate2231(.a(s_241), .O(gate398inter4));
  nand2 gate2232(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2233(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2234(.a(G12), .O(gate398inter7));
  inv1  gate2235(.a(G1069), .O(gate398inter8));
  nand2 gate2236(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2237(.a(s_241), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2238(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2239(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2240(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1401(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1402(.a(gate400inter0), .b(s_122), .O(gate400inter1));
  and2  gate1403(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1404(.a(s_122), .O(gate400inter3));
  inv1  gate1405(.a(s_123), .O(gate400inter4));
  nand2 gate1406(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1407(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1408(.a(G14), .O(gate400inter7));
  inv1  gate1409(.a(G1075), .O(gate400inter8));
  nand2 gate1410(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1411(.a(s_123), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1412(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1413(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1414(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2563(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2564(.a(gate401inter0), .b(s_288), .O(gate401inter1));
  and2  gate2565(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2566(.a(s_288), .O(gate401inter3));
  inv1  gate2567(.a(s_289), .O(gate401inter4));
  nand2 gate2568(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2569(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2570(.a(G15), .O(gate401inter7));
  inv1  gate2571(.a(G1078), .O(gate401inter8));
  nand2 gate2572(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2573(.a(s_289), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2574(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2575(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2576(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2521(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2522(.a(gate408inter0), .b(s_282), .O(gate408inter1));
  and2  gate2523(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2524(.a(s_282), .O(gate408inter3));
  inv1  gate2525(.a(s_283), .O(gate408inter4));
  nand2 gate2526(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2527(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2528(.a(G22), .O(gate408inter7));
  inv1  gate2529(.a(G1099), .O(gate408inter8));
  nand2 gate2530(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2531(.a(s_283), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2532(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2533(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2534(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2493(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2494(.a(gate411inter0), .b(s_278), .O(gate411inter1));
  and2  gate2495(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2496(.a(s_278), .O(gate411inter3));
  inv1  gate2497(.a(s_279), .O(gate411inter4));
  nand2 gate2498(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2499(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2500(.a(G25), .O(gate411inter7));
  inv1  gate2501(.a(G1108), .O(gate411inter8));
  nand2 gate2502(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2503(.a(s_279), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2504(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2505(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2506(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate883(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate884(.a(gate412inter0), .b(s_48), .O(gate412inter1));
  and2  gate885(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate886(.a(s_48), .O(gate412inter3));
  inv1  gate887(.a(s_49), .O(gate412inter4));
  nand2 gate888(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate889(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate890(.a(G26), .O(gate412inter7));
  inv1  gate891(.a(G1111), .O(gate412inter8));
  nand2 gate892(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate893(.a(s_49), .b(gate412inter3), .O(gate412inter10));
  nor2  gate894(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate895(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate896(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate3039(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate3040(.a(gate414inter0), .b(s_356), .O(gate414inter1));
  and2  gate3041(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate3042(.a(s_356), .O(gate414inter3));
  inv1  gate3043(.a(s_357), .O(gate414inter4));
  nand2 gate3044(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate3045(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate3046(.a(G28), .O(gate414inter7));
  inv1  gate3047(.a(G1117), .O(gate414inter8));
  nand2 gate3048(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate3049(.a(s_357), .b(gate414inter3), .O(gate414inter10));
  nor2  gate3050(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate3051(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate3052(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1961(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1962(.a(gate415inter0), .b(s_202), .O(gate415inter1));
  and2  gate1963(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1964(.a(s_202), .O(gate415inter3));
  inv1  gate1965(.a(s_203), .O(gate415inter4));
  nand2 gate1966(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1967(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1968(.a(G29), .O(gate415inter7));
  inv1  gate1969(.a(G1120), .O(gate415inter8));
  nand2 gate1970(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1971(.a(s_203), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1972(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1973(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1974(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate547(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate548(.a(gate416inter0), .b(s_0), .O(gate416inter1));
  and2  gate549(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate550(.a(s_0), .O(gate416inter3));
  inv1  gate551(.a(s_1), .O(gate416inter4));
  nand2 gate552(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate553(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate554(.a(G30), .O(gate416inter7));
  inv1  gate555(.a(G1123), .O(gate416inter8));
  nand2 gate556(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate557(.a(s_1), .b(gate416inter3), .O(gate416inter10));
  nor2  gate558(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate559(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate560(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2185(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2186(.a(gate418inter0), .b(s_234), .O(gate418inter1));
  and2  gate2187(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2188(.a(s_234), .O(gate418inter3));
  inv1  gate2189(.a(s_235), .O(gate418inter4));
  nand2 gate2190(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2191(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2192(.a(G32), .O(gate418inter7));
  inv1  gate2193(.a(G1129), .O(gate418inter8));
  nand2 gate2194(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2195(.a(s_235), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2196(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2197(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2198(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2605(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2606(.a(gate419inter0), .b(s_294), .O(gate419inter1));
  and2  gate2607(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2608(.a(s_294), .O(gate419inter3));
  inv1  gate2609(.a(s_295), .O(gate419inter4));
  nand2 gate2610(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2611(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2612(.a(G1), .O(gate419inter7));
  inv1  gate2613(.a(G1132), .O(gate419inter8));
  nand2 gate2614(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2615(.a(s_295), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2616(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2617(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2618(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate3025(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate3026(.a(gate420inter0), .b(s_354), .O(gate420inter1));
  and2  gate3027(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate3028(.a(s_354), .O(gate420inter3));
  inv1  gate3029(.a(s_355), .O(gate420inter4));
  nand2 gate3030(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate3031(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate3032(.a(G1036), .O(gate420inter7));
  inv1  gate3033(.a(G1132), .O(gate420inter8));
  nand2 gate3034(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate3035(.a(s_355), .b(gate420inter3), .O(gate420inter10));
  nor2  gate3036(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate3037(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate3038(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate2423(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2424(.a(gate421inter0), .b(s_268), .O(gate421inter1));
  and2  gate2425(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2426(.a(s_268), .O(gate421inter3));
  inv1  gate2427(.a(s_269), .O(gate421inter4));
  nand2 gate2428(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2429(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2430(.a(G2), .O(gate421inter7));
  inv1  gate2431(.a(G1135), .O(gate421inter8));
  nand2 gate2432(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2433(.a(s_269), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2434(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2435(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2436(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2507(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2508(.a(gate422inter0), .b(s_280), .O(gate422inter1));
  and2  gate2509(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2510(.a(s_280), .O(gate422inter3));
  inv1  gate2511(.a(s_281), .O(gate422inter4));
  nand2 gate2512(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2513(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2514(.a(G1039), .O(gate422inter7));
  inv1  gate2515(.a(G1135), .O(gate422inter8));
  nand2 gate2516(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2517(.a(s_281), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2518(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2519(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2520(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2241(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2242(.a(gate425inter0), .b(s_242), .O(gate425inter1));
  and2  gate2243(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2244(.a(s_242), .O(gate425inter3));
  inv1  gate2245(.a(s_243), .O(gate425inter4));
  nand2 gate2246(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2247(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2248(.a(G4), .O(gate425inter7));
  inv1  gate2249(.a(G1141), .O(gate425inter8));
  nand2 gate2250(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2251(.a(s_243), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2252(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2253(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2254(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1723(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1724(.a(gate426inter0), .b(s_168), .O(gate426inter1));
  and2  gate1725(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1726(.a(s_168), .O(gate426inter3));
  inv1  gate1727(.a(s_169), .O(gate426inter4));
  nand2 gate1728(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1729(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1730(.a(G1045), .O(gate426inter7));
  inv1  gate1731(.a(G1141), .O(gate426inter8));
  nand2 gate1732(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1733(.a(s_169), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1734(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1735(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1736(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1863(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1864(.a(gate427inter0), .b(s_188), .O(gate427inter1));
  and2  gate1865(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1866(.a(s_188), .O(gate427inter3));
  inv1  gate1867(.a(s_189), .O(gate427inter4));
  nand2 gate1868(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1869(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1870(.a(G5), .O(gate427inter7));
  inv1  gate1871(.a(G1144), .O(gate427inter8));
  nand2 gate1872(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1873(.a(s_189), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1874(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1875(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1876(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2773(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2774(.a(gate429inter0), .b(s_318), .O(gate429inter1));
  and2  gate2775(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2776(.a(s_318), .O(gate429inter3));
  inv1  gate2777(.a(s_319), .O(gate429inter4));
  nand2 gate2778(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2779(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2780(.a(G6), .O(gate429inter7));
  inv1  gate2781(.a(G1147), .O(gate429inter8));
  nand2 gate2782(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2783(.a(s_319), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2784(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2785(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2786(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate575(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate576(.a(gate430inter0), .b(s_4), .O(gate430inter1));
  and2  gate577(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate578(.a(s_4), .O(gate430inter3));
  inv1  gate579(.a(s_5), .O(gate430inter4));
  nand2 gate580(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate581(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate582(.a(G1051), .O(gate430inter7));
  inv1  gate583(.a(G1147), .O(gate430inter8));
  nand2 gate584(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate585(.a(s_5), .b(gate430inter3), .O(gate430inter10));
  nor2  gate586(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate587(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate588(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2045(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2046(.a(gate432inter0), .b(s_214), .O(gate432inter1));
  and2  gate2047(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2048(.a(s_214), .O(gate432inter3));
  inv1  gate2049(.a(s_215), .O(gate432inter4));
  nand2 gate2050(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2051(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2052(.a(G1054), .O(gate432inter7));
  inv1  gate2053(.a(G1150), .O(gate432inter8));
  nand2 gate2054(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2055(.a(s_215), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2056(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2057(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2058(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2997(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2998(.a(gate434inter0), .b(s_350), .O(gate434inter1));
  and2  gate2999(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate3000(.a(s_350), .O(gate434inter3));
  inv1  gate3001(.a(s_351), .O(gate434inter4));
  nand2 gate3002(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate3003(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate3004(.a(G1057), .O(gate434inter7));
  inv1  gate3005(.a(G1153), .O(gate434inter8));
  nand2 gate3006(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate3007(.a(s_351), .b(gate434inter3), .O(gate434inter10));
  nor2  gate3008(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate3009(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate3010(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2381(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2382(.a(gate435inter0), .b(s_262), .O(gate435inter1));
  and2  gate2383(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2384(.a(s_262), .O(gate435inter3));
  inv1  gate2385(.a(s_263), .O(gate435inter4));
  nand2 gate2386(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2387(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2388(.a(G9), .O(gate435inter7));
  inv1  gate2389(.a(G1156), .O(gate435inter8));
  nand2 gate2390(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2391(.a(s_263), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2392(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2393(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2394(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1919(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1920(.a(gate437inter0), .b(s_196), .O(gate437inter1));
  and2  gate1921(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1922(.a(s_196), .O(gate437inter3));
  inv1  gate1923(.a(s_197), .O(gate437inter4));
  nand2 gate1924(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1925(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1926(.a(G10), .O(gate437inter7));
  inv1  gate1927(.a(G1159), .O(gate437inter8));
  nand2 gate1928(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1929(.a(s_197), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1930(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1931(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1932(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2759(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2760(.a(gate438inter0), .b(s_316), .O(gate438inter1));
  and2  gate2761(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2762(.a(s_316), .O(gate438inter3));
  inv1  gate2763(.a(s_317), .O(gate438inter4));
  nand2 gate2764(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2765(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2766(.a(G1063), .O(gate438inter7));
  inv1  gate2767(.a(G1159), .O(gate438inter8));
  nand2 gate2768(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2769(.a(s_317), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2770(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2771(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2772(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1009(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1010(.a(gate440inter0), .b(s_66), .O(gate440inter1));
  and2  gate1011(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1012(.a(s_66), .O(gate440inter3));
  inv1  gate1013(.a(s_67), .O(gate440inter4));
  nand2 gate1014(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1015(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1016(.a(G1066), .O(gate440inter7));
  inv1  gate1017(.a(G1162), .O(gate440inter8));
  nand2 gate1018(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1019(.a(s_67), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1020(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1021(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1022(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2059(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2060(.a(gate443inter0), .b(s_216), .O(gate443inter1));
  and2  gate2061(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2062(.a(s_216), .O(gate443inter3));
  inv1  gate2063(.a(s_217), .O(gate443inter4));
  nand2 gate2064(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2065(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2066(.a(G13), .O(gate443inter7));
  inv1  gate2067(.a(G1168), .O(gate443inter8));
  nand2 gate2068(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2069(.a(s_217), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2070(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2071(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2072(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate743(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate744(.a(gate444inter0), .b(s_28), .O(gate444inter1));
  and2  gate745(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate746(.a(s_28), .O(gate444inter3));
  inv1  gate747(.a(s_29), .O(gate444inter4));
  nand2 gate748(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate749(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate750(.a(G1072), .O(gate444inter7));
  inv1  gate751(.a(G1168), .O(gate444inter8));
  nand2 gate752(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate753(.a(s_29), .b(gate444inter3), .O(gate444inter10));
  nor2  gate754(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate755(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate756(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1849(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1850(.a(gate445inter0), .b(s_186), .O(gate445inter1));
  and2  gate1851(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1852(.a(s_186), .O(gate445inter3));
  inv1  gate1853(.a(s_187), .O(gate445inter4));
  nand2 gate1854(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1855(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1856(.a(G14), .O(gate445inter7));
  inv1  gate1857(.a(G1171), .O(gate445inter8));
  nand2 gate1858(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1859(.a(s_187), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1860(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1861(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1862(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1583(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1584(.a(gate448inter0), .b(s_148), .O(gate448inter1));
  and2  gate1585(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1586(.a(s_148), .O(gate448inter3));
  inv1  gate1587(.a(s_149), .O(gate448inter4));
  nand2 gate1588(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1589(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1590(.a(G1078), .O(gate448inter7));
  inv1  gate1591(.a(G1174), .O(gate448inter8));
  nand2 gate1592(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1593(.a(s_149), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1594(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1595(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1596(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2213(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2214(.a(gate450inter0), .b(s_238), .O(gate450inter1));
  and2  gate2215(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2216(.a(s_238), .O(gate450inter3));
  inv1  gate2217(.a(s_239), .O(gate450inter4));
  nand2 gate2218(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2219(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2220(.a(G1081), .O(gate450inter7));
  inv1  gate2221(.a(G1177), .O(gate450inter8));
  nand2 gate2222(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2223(.a(s_239), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2224(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2225(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2226(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate561(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate562(.a(gate454inter0), .b(s_2), .O(gate454inter1));
  and2  gate563(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate564(.a(s_2), .O(gate454inter3));
  inv1  gate565(.a(s_3), .O(gate454inter4));
  nand2 gate566(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate567(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate568(.a(G1087), .O(gate454inter7));
  inv1  gate569(.a(G1183), .O(gate454inter8));
  nand2 gate570(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate571(.a(s_3), .b(gate454inter3), .O(gate454inter10));
  nor2  gate572(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate573(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate574(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1877(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1878(.a(gate455inter0), .b(s_190), .O(gate455inter1));
  and2  gate1879(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1880(.a(s_190), .O(gate455inter3));
  inv1  gate1881(.a(s_191), .O(gate455inter4));
  nand2 gate1882(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1883(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1884(.a(G19), .O(gate455inter7));
  inv1  gate1885(.a(G1186), .O(gate455inter8));
  nand2 gate1886(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1887(.a(s_191), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1888(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1889(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1890(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2633(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2634(.a(gate458inter0), .b(s_298), .O(gate458inter1));
  and2  gate2635(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2636(.a(s_298), .O(gate458inter3));
  inv1  gate2637(.a(s_299), .O(gate458inter4));
  nand2 gate2638(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2639(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2640(.a(G1093), .O(gate458inter7));
  inv1  gate2641(.a(G1189), .O(gate458inter8));
  nand2 gate2642(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2643(.a(s_299), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2644(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2645(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2646(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1359(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1360(.a(gate459inter0), .b(s_116), .O(gate459inter1));
  and2  gate1361(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1362(.a(s_116), .O(gate459inter3));
  inv1  gate1363(.a(s_117), .O(gate459inter4));
  nand2 gate1364(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1365(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1366(.a(G21), .O(gate459inter7));
  inv1  gate1367(.a(G1192), .O(gate459inter8));
  nand2 gate1368(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1369(.a(s_117), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1370(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1371(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1372(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2451(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2452(.a(gate462inter0), .b(s_272), .O(gate462inter1));
  and2  gate2453(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2454(.a(s_272), .O(gate462inter3));
  inv1  gate2455(.a(s_273), .O(gate462inter4));
  nand2 gate2456(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2457(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2458(.a(G1099), .O(gate462inter7));
  inv1  gate2459(.a(G1195), .O(gate462inter8));
  nand2 gate2460(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2461(.a(s_273), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2462(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2463(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2464(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate2101(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2102(.a(gate464inter0), .b(s_222), .O(gate464inter1));
  and2  gate2103(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2104(.a(s_222), .O(gate464inter3));
  inv1  gate2105(.a(s_223), .O(gate464inter4));
  nand2 gate2106(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2107(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2108(.a(G1102), .O(gate464inter7));
  inv1  gate2109(.a(G1198), .O(gate464inter8));
  nand2 gate2110(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2111(.a(s_223), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2112(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2113(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2114(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1639(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1640(.a(gate465inter0), .b(s_156), .O(gate465inter1));
  and2  gate1641(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1642(.a(s_156), .O(gate465inter3));
  inv1  gate1643(.a(s_157), .O(gate465inter4));
  nand2 gate1644(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1645(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1646(.a(G24), .O(gate465inter7));
  inv1  gate1647(.a(G1201), .O(gate465inter8));
  nand2 gate1648(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1649(.a(s_157), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1650(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1651(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1652(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2143(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2144(.a(gate466inter0), .b(s_228), .O(gate466inter1));
  and2  gate2145(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2146(.a(s_228), .O(gate466inter3));
  inv1  gate2147(.a(s_229), .O(gate466inter4));
  nand2 gate2148(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2149(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2150(.a(G1105), .O(gate466inter7));
  inv1  gate2151(.a(G1201), .O(gate466inter8));
  nand2 gate2152(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2153(.a(s_229), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2154(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2155(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2156(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1947(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1948(.a(gate467inter0), .b(s_200), .O(gate467inter1));
  and2  gate1949(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1950(.a(s_200), .O(gate467inter3));
  inv1  gate1951(.a(s_201), .O(gate467inter4));
  nand2 gate1952(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1953(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1954(.a(G25), .O(gate467inter7));
  inv1  gate1955(.a(G1204), .O(gate467inter8));
  nand2 gate1956(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1957(.a(s_201), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1958(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1959(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1960(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2157(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2158(.a(gate471inter0), .b(s_230), .O(gate471inter1));
  and2  gate2159(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2160(.a(s_230), .O(gate471inter3));
  inv1  gate2161(.a(s_231), .O(gate471inter4));
  nand2 gate2162(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2163(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2164(.a(G27), .O(gate471inter7));
  inv1  gate2165(.a(G1210), .O(gate471inter8));
  nand2 gate2166(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2167(.a(s_231), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2168(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2169(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2170(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2913(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2914(.a(gate477inter0), .b(s_338), .O(gate477inter1));
  and2  gate2915(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2916(.a(s_338), .O(gate477inter3));
  inv1  gate2917(.a(s_339), .O(gate477inter4));
  nand2 gate2918(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2919(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2920(.a(G30), .O(gate477inter7));
  inv1  gate2921(.a(G1219), .O(gate477inter8));
  nand2 gate2922(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2923(.a(s_339), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2924(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2925(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2926(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2031(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2032(.a(gate486inter0), .b(s_212), .O(gate486inter1));
  and2  gate2033(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2034(.a(s_212), .O(gate486inter3));
  inv1  gate2035(.a(s_213), .O(gate486inter4));
  nand2 gate2036(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2037(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2038(.a(G1234), .O(gate486inter7));
  inv1  gate2039(.a(G1235), .O(gate486inter8));
  nand2 gate2040(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2041(.a(s_213), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2042(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2043(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2044(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate1695(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1696(.a(gate487inter0), .b(s_164), .O(gate487inter1));
  and2  gate1697(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1698(.a(s_164), .O(gate487inter3));
  inv1  gate1699(.a(s_165), .O(gate487inter4));
  nand2 gate1700(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1701(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1702(.a(G1236), .O(gate487inter7));
  inv1  gate1703(.a(G1237), .O(gate487inter8));
  nand2 gate1704(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1705(.a(s_165), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1706(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1707(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1708(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1303(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1304(.a(gate489inter0), .b(s_108), .O(gate489inter1));
  and2  gate1305(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1306(.a(s_108), .O(gate489inter3));
  inv1  gate1307(.a(s_109), .O(gate489inter4));
  nand2 gate1308(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1309(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1310(.a(G1240), .O(gate489inter7));
  inv1  gate1311(.a(G1241), .O(gate489inter8));
  nand2 gate1312(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1313(.a(s_109), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1314(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1315(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1316(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1975(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1976(.a(gate491inter0), .b(s_204), .O(gate491inter1));
  and2  gate1977(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1978(.a(s_204), .O(gate491inter3));
  inv1  gate1979(.a(s_205), .O(gate491inter4));
  nand2 gate1980(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1981(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1982(.a(G1244), .O(gate491inter7));
  inv1  gate1983(.a(G1245), .O(gate491inter8));
  nand2 gate1984(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1985(.a(s_205), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1986(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1987(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1988(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate813(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate814(.a(gate492inter0), .b(s_38), .O(gate492inter1));
  and2  gate815(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate816(.a(s_38), .O(gate492inter3));
  inv1  gate817(.a(s_39), .O(gate492inter4));
  nand2 gate818(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate819(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate820(.a(G1246), .O(gate492inter7));
  inv1  gate821(.a(G1247), .O(gate492inter8));
  nand2 gate822(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate823(.a(s_39), .b(gate492inter3), .O(gate492inter10));
  nor2  gate824(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate825(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate826(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2703(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2704(.a(gate497inter0), .b(s_308), .O(gate497inter1));
  and2  gate2705(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2706(.a(s_308), .O(gate497inter3));
  inv1  gate2707(.a(s_309), .O(gate497inter4));
  nand2 gate2708(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2709(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2710(.a(G1256), .O(gate497inter7));
  inv1  gate2711(.a(G1257), .O(gate497inter8));
  nand2 gate2712(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2713(.a(s_309), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2714(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2715(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2716(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1471(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1472(.a(gate498inter0), .b(s_132), .O(gate498inter1));
  and2  gate1473(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1474(.a(s_132), .O(gate498inter3));
  inv1  gate1475(.a(s_133), .O(gate498inter4));
  nand2 gate1476(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1477(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1478(.a(G1258), .O(gate498inter7));
  inv1  gate1479(.a(G1259), .O(gate498inter8));
  nand2 gate1480(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1481(.a(s_133), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1482(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1483(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1484(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1387(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1388(.a(gate500inter0), .b(s_120), .O(gate500inter1));
  and2  gate1389(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1390(.a(s_120), .O(gate500inter3));
  inv1  gate1391(.a(s_121), .O(gate500inter4));
  nand2 gate1392(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1393(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1394(.a(G1262), .O(gate500inter7));
  inv1  gate1395(.a(G1263), .O(gate500inter8));
  nand2 gate1396(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1397(.a(s_121), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1398(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1399(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1400(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1611(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1612(.a(gate503inter0), .b(s_152), .O(gate503inter1));
  and2  gate1613(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1614(.a(s_152), .O(gate503inter3));
  inv1  gate1615(.a(s_153), .O(gate503inter4));
  nand2 gate1616(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1617(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1618(.a(G1268), .O(gate503inter7));
  inv1  gate1619(.a(G1269), .O(gate503inter8));
  nand2 gate1620(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1621(.a(s_153), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1622(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1623(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1624(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate757(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate758(.a(gate504inter0), .b(s_30), .O(gate504inter1));
  and2  gate759(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate760(.a(s_30), .O(gate504inter3));
  inv1  gate761(.a(s_31), .O(gate504inter4));
  nand2 gate762(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate763(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate764(.a(G1270), .O(gate504inter7));
  inv1  gate765(.a(G1271), .O(gate504inter8));
  nand2 gate766(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate767(.a(s_31), .b(gate504inter3), .O(gate504inter10));
  nor2  gate768(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate769(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate770(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1121(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1122(.a(gate506inter0), .b(s_82), .O(gate506inter1));
  and2  gate1123(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1124(.a(s_82), .O(gate506inter3));
  inv1  gate1125(.a(s_83), .O(gate506inter4));
  nand2 gate1126(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1127(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1128(.a(G1274), .O(gate506inter7));
  inv1  gate1129(.a(G1275), .O(gate506inter8));
  nand2 gate1130(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1131(.a(s_83), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1132(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1133(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1134(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate981(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate982(.a(gate509inter0), .b(s_62), .O(gate509inter1));
  and2  gate983(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate984(.a(s_62), .O(gate509inter3));
  inv1  gate985(.a(s_63), .O(gate509inter4));
  nand2 gate986(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate987(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate988(.a(G1280), .O(gate509inter7));
  inv1  gate989(.a(G1281), .O(gate509inter8));
  nand2 gate990(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate991(.a(s_63), .b(gate509inter3), .O(gate509inter10));
  nor2  gate992(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate993(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate994(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1807(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1808(.a(gate512inter0), .b(s_180), .O(gate512inter1));
  and2  gate1809(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1810(.a(s_180), .O(gate512inter3));
  inv1  gate1811(.a(s_181), .O(gate512inter4));
  nand2 gate1812(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1813(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1814(.a(G1286), .O(gate512inter7));
  inv1  gate1815(.a(G1287), .O(gate512inter8));
  nand2 gate1816(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1817(.a(s_181), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1818(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1819(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1820(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule