module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1499(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1500(.a(gate11inter0), .b(s_136), .O(gate11inter1));
  and2  gate1501(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1502(.a(s_136), .O(gate11inter3));
  inv1  gate1503(.a(s_137), .O(gate11inter4));
  nand2 gate1504(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1505(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1506(.a(G5), .O(gate11inter7));
  inv1  gate1507(.a(G6), .O(gate11inter8));
  nand2 gate1508(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1509(.a(s_137), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1510(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1511(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1512(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2045(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2046(.a(gate12inter0), .b(s_214), .O(gate12inter1));
  and2  gate2047(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2048(.a(s_214), .O(gate12inter3));
  inv1  gate2049(.a(s_215), .O(gate12inter4));
  nand2 gate2050(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2051(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2052(.a(G7), .O(gate12inter7));
  inv1  gate2053(.a(G8), .O(gate12inter8));
  nand2 gate2054(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2055(.a(s_215), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2056(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2057(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2058(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2255(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2256(.a(gate16inter0), .b(s_244), .O(gate16inter1));
  and2  gate2257(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2258(.a(s_244), .O(gate16inter3));
  inv1  gate2259(.a(s_245), .O(gate16inter4));
  nand2 gate2260(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2261(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2262(.a(G15), .O(gate16inter7));
  inv1  gate2263(.a(G16), .O(gate16inter8));
  nand2 gate2264(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2265(.a(s_245), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2266(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2267(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2268(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2031(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2032(.a(gate19inter0), .b(s_212), .O(gate19inter1));
  and2  gate2033(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2034(.a(s_212), .O(gate19inter3));
  inv1  gate2035(.a(s_213), .O(gate19inter4));
  nand2 gate2036(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2037(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2038(.a(G21), .O(gate19inter7));
  inv1  gate2039(.a(G22), .O(gate19inter8));
  nand2 gate2040(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2041(.a(s_213), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2042(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2043(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2044(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1429(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1430(.a(gate20inter0), .b(s_126), .O(gate20inter1));
  and2  gate1431(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1432(.a(s_126), .O(gate20inter3));
  inv1  gate1433(.a(s_127), .O(gate20inter4));
  nand2 gate1434(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1435(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1436(.a(G23), .O(gate20inter7));
  inv1  gate1437(.a(G24), .O(gate20inter8));
  nand2 gate1438(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1439(.a(s_127), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1440(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1441(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1442(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1191(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1192(.a(gate26inter0), .b(s_92), .O(gate26inter1));
  and2  gate1193(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1194(.a(s_92), .O(gate26inter3));
  inv1  gate1195(.a(s_93), .O(gate26inter4));
  nand2 gate1196(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1197(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1198(.a(G9), .O(gate26inter7));
  inv1  gate1199(.a(G13), .O(gate26inter8));
  nand2 gate1200(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1201(.a(s_93), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1202(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1203(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1204(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1793(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1794(.a(gate30inter0), .b(s_178), .O(gate30inter1));
  and2  gate1795(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1796(.a(s_178), .O(gate30inter3));
  inv1  gate1797(.a(s_179), .O(gate30inter4));
  nand2 gate1798(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1799(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1800(.a(G11), .O(gate30inter7));
  inv1  gate1801(.a(G15), .O(gate30inter8));
  nand2 gate1802(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1803(.a(s_179), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1804(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1805(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1806(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate813(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate814(.a(gate31inter0), .b(s_38), .O(gate31inter1));
  and2  gate815(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate816(.a(s_38), .O(gate31inter3));
  inv1  gate817(.a(s_39), .O(gate31inter4));
  nand2 gate818(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate819(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate820(.a(G4), .O(gate31inter7));
  inv1  gate821(.a(G8), .O(gate31inter8));
  nand2 gate822(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate823(.a(s_39), .b(gate31inter3), .O(gate31inter10));
  nor2  gate824(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate825(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate826(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate827(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate828(.a(gate34inter0), .b(s_40), .O(gate34inter1));
  and2  gate829(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate830(.a(s_40), .O(gate34inter3));
  inv1  gate831(.a(s_41), .O(gate34inter4));
  nand2 gate832(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate833(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate834(.a(G25), .O(gate34inter7));
  inv1  gate835(.a(G29), .O(gate34inter8));
  nand2 gate836(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate837(.a(s_41), .b(gate34inter3), .O(gate34inter10));
  nor2  gate838(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate839(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate840(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate2059(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2060(.a(gate35inter0), .b(s_216), .O(gate35inter1));
  and2  gate2061(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2062(.a(s_216), .O(gate35inter3));
  inv1  gate2063(.a(s_217), .O(gate35inter4));
  nand2 gate2064(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2065(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2066(.a(G18), .O(gate35inter7));
  inv1  gate2067(.a(G22), .O(gate35inter8));
  nand2 gate2068(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2069(.a(s_217), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2070(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2071(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2072(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1443(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1444(.a(gate37inter0), .b(s_128), .O(gate37inter1));
  and2  gate1445(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1446(.a(s_128), .O(gate37inter3));
  inv1  gate1447(.a(s_129), .O(gate37inter4));
  nand2 gate1448(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1449(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1450(.a(G19), .O(gate37inter7));
  inv1  gate1451(.a(G23), .O(gate37inter8));
  nand2 gate1452(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1453(.a(s_129), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1454(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1455(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1456(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate785(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate786(.a(gate39inter0), .b(s_34), .O(gate39inter1));
  and2  gate787(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate788(.a(s_34), .O(gate39inter3));
  inv1  gate789(.a(s_35), .O(gate39inter4));
  nand2 gate790(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate791(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate792(.a(G20), .O(gate39inter7));
  inv1  gate793(.a(G24), .O(gate39inter8));
  nand2 gate794(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate795(.a(s_35), .b(gate39inter3), .O(gate39inter10));
  nor2  gate796(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate797(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate798(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2213(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2214(.a(gate42inter0), .b(s_238), .O(gate42inter1));
  and2  gate2215(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2216(.a(s_238), .O(gate42inter3));
  inv1  gate2217(.a(s_239), .O(gate42inter4));
  nand2 gate2218(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2219(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2220(.a(G2), .O(gate42inter7));
  inv1  gate2221(.a(G266), .O(gate42inter8));
  nand2 gate2222(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2223(.a(s_239), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2224(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2225(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2226(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate645(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate646(.a(gate43inter0), .b(s_14), .O(gate43inter1));
  and2  gate647(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate648(.a(s_14), .O(gate43inter3));
  inv1  gate649(.a(s_15), .O(gate43inter4));
  nand2 gate650(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate651(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate652(.a(G3), .O(gate43inter7));
  inv1  gate653(.a(G269), .O(gate43inter8));
  nand2 gate654(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate655(.a(s_15), .b(gate43inter3), .O(gate43inter10));
  nor2  gate656(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate657(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate658(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2171(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2172(.a(gate44inter0), .b(s_232), .O(gate44inter1));
  and2  gate2173(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2174(.a(s_232), .O(gate44inter3));
  inv1  gate2175(.a(s_233), .O(gate44inter4));
  nand2 gate2176(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2177(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2178(.a(G4), .O(gate44inter7));
  inv1  gate2179(.a(G269), .O(gate44inter8));
  nand2 gate2180(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2181(.a(s_233), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2182(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2183(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2184(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2101(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2102(.a(gate45inter0), .b(s_222), .O(gate45inter1));
  and2  gate2103(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2104(.a(s_222), .O(gate45inter3));
  inv1  gate2105(.a(s_223), .O(gate45inter4));
  nand2 gate2106(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2107(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2108(.a(G5), .O(gate45inter7));
  inv1  gate2109(.a(G272), .O(gate45inter8));
  nand2 gate2110(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2111(.a(s_223), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2112(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2113(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2114(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1331(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1332(.a(gate49inter0), .b(s_112), .O(gate49inter1));
  and2  gate1333(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1334(.a(s_112), .O(gate49inter3));
  inv1  gate1335(.a(s_113), .O(gate49inter4));
  nand2 gate1336(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1337(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1338(.a(G9), .O(gate49inter7));
  inv1  gate1339(.a(G278), .O(gate49inter8));
  nand2 gate1340(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1341(.a(s_113), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1342(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1343(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1344(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1345(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1346(.a(gate66inter0), .b(s_114), .O(gate66inter1));
  and2  gate1347(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1348(.a(s_114), .O(gate66inter3));
  inv1  gate1349(.a(s_115), .O(gate66inter4));
  nand2 gate1350(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1351(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1352(.a(G26), .O(gate66inter7));
  inv1  gate1353(.a(G302), .O(gate66inter8));
  nand2 gate1354(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1355(.a(s_115), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1356(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1357(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1358(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate743(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate744(.a(gate72inter0), .b(s_28), .O(gate72inter1));
  and2  gate745(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate746(.a(s_28), .O(gate72inter3));
  inv1  gate747(.a(s_29), .O(gate72inter4));
  nand2 gate748(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate749(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate750(.a(G32), .O(gate72inter7));
  inv1  gate751(.a(G311), .O(gate72inter8));
  nand2 gate752(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate753(.a(s_29), .b(gate72inter3), .O(gate72inter10));
  nor2  gate754(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate755(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate756(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1373(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1374(.a(gate75inter0), .b(s_118), .O(gate75inter1));
  and2  gate1375(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1376(.a(s_118), .O(gate75inter3));
  inv1  gate1377(.a(s_119), .O(gate75inter4));
  nand2 gate1378(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1379(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1380(.a(G9), .O(gate75inter7));
  inv1  gate1381(.a(G317), .O(gate75inter8));
  nand2 gate1382(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1383(.a(s_119), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1384(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1385(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1386(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate603(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate604(.a(gate76inter0), .b(s_8), .O(gate76inter1));
  and2  gate605(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate606(.a(s_8), .O(gate76inter3));
  inv1  gate607(.a(s_9), .O(gate76inter4));
  nand2 gate608(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate609(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate610(.a(G13), .O(gate76inter7));
  inv1  gate611(.a(G317), .O(gate76inter8));
  nand2 gate612(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate613(.a(s_9), .b(gate76inter3), .O(gate76inter10));
  nor2  gate614(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate615(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate616(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1765(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1766(.a(gate77inter0), .b(s_174), .O(gate77inter1));
  and2  gate1767(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1768(.a(s_174), .O(gate77inter3));
  inv1  gate1769(.a(s_175), .O(gate77inter4));
  nand2 gate1770(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1771(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1772(.a(G2), .O(gate77inter7));
  inv1  gate1773(.a(G320), .O(gate77inter8));
  nand2 gate1774(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1775(.a(s_175), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1776(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1777(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1778(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1359(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1360(.a(gate78inter0), .b(s_116), .O(gate78inter1));
  and2  gate1361(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1362(.a(s_116), .O(gate78inter3));
  inv1  gate1363(.a(s_117), .O(gate78inter4));
  nand2 gate1364(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1365(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1366(.a(G6), .O(gate78inter7));
  inv1  gate1367(.a(G320), .O(gate78inter8));
  nand2 gate1368(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1369(.a(s_117), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1370(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1371(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1372(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate883(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate884(.a(gate79inter0), .b(s_48), .O(gate79inter1));
  and2  gate885(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate886(.a(s_48), .O(gate79inter3));
  inv1  gate887(.a(s_49), .O(gate79inter4));
  nand2 gate888(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate889(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate890(.a(G10), .O(gate79inter7));
  inv1  gate891(.a(G323), .O(gate79inter8));
  nand2 gate892(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate893(.a(s_49), .b(gate79inter3), .O(gate79inter10));
  nor2  gate894(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate895(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate896(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1135(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1136(.a(gate80inter0), .b(s_84), .O(gate80inter1));
  and2  gate1137(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1138(.a(s_84), .O(gate80inter3));
  inv1  gate1139(.a(s_85), .O(gate80inter4));
  nand2 gate1140(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1141(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1142(.a(G14), .O(gate80inter7));
  inv1  gate1143(.a(G323), .O(gate80inter8));
  nand2 gate1144(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1145(.a(s_85), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1146(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1147(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1148(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1079(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1080(.a(gate81inter0), .b(s_76), .O(gate81inter1));
  and2  gate1081(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1082(.a(s_76), .O(gate81inter3));
  inv1  gate1083(.a(s_77), .O(gate81inter4));
  nand2 gate1084(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1085(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1086(.a(G3), .O(gate81inter7));
  inv1  gate1087(.a(G326), .O(gate81inter8));
  nand2 gate1088(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1089(.a(s_77), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1090(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1091(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1092(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate2325(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2326(.a(gate83inter0), .b(s_254), .O(gate83inter1));
  and2  gate2327(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2328(.a(s_254), .O(gate83inter3));
  inv1  gate2329(.a(s_255), .O(gate83inter4));
  nand2 gate2330(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2331(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2332(.a(G11), .O(gate83inter7));
  inv1  gate2333(.a(G329), .O(gate83inter8));
  nand2 gate2334(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2335(.a(s_255), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2336(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2337(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2338(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate715(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate716(.a(gate88inter0), .b(s_24), .O(gate88inter1));
  and2  gate717(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate718(.a(s_24), .O(gate88inter3));
  inv1  gate719(.a(s_25), .O(gate88inter4));
  nand2 gate720(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate721(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate722(.a(G16), .O(gate88inter7));
  inv1  gate723(.a(G335), .O(gate88inter8));
  nand2 gate724(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate725(.a(s_25), .b(gate88inter3), .O(gate88inter10));
  nor2  gate726(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate727(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate728(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1667(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1668(.a(gate90inter0), .b(s_160), .O(gate90inter1));
  and2  gate1669(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1670(.a(s_160), .O(gate90inter3));
  inv1  gate1671(.a(s_161), .O(gate90inter4));
  nand2 gate1672(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1673(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1674(.a(G21), .O(gate90inter7));
  inv1  gate1675(.a(G338), .O(gate90inter8));
  nand2 gate1676(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1677(.a(s_161), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1678(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1679(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1680(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1275(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1276(.a(gate97inter0), .b(s_104), .O(gate97inter1));
  and2  gate1277(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1278(.a(s_104), .O(gate97inter3));
  inv1  gate1279(.a(s_105), .O(gate97inter4));
  nand2 gate1280(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1281(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1282(.a(G19), .O(gate97inter7));
  inv1  gate1283(.a(G350), .O(gate97inter8));
  nand2 gate1284(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1285(.a(s_105), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1286(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1287(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1288(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1387(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1388(.a(gate100inter0), .b(s_120), .O(gate100inter1));
  and2  gate1389(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1390(.a(s_120), .O(gate100inter3));
  inv1  gate1391(.a(s_121), .O(gate100inter4));
  nand2 gate1392(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1393(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1394(.a(G31), .O(gate100inter7));
  inv1  gate1395(.a(G353), .O(gate100inter8));
  nand2 gate1396(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1397(.a(s_121), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1398(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1399(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1400(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1891(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1892(.a(gate102inter0), .b(s_192), .O(gate102inter1));
  and2  gate1893(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1894(.a(s_192), .O(gate102inter3));
  inv1  gate1895(.a(s_193), .O(gate102inter4));
  nand2 gate1896(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1897(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1898(.a(G24), .O(gate102inter7));
  inv1  gate1899(.a(G356), .O(gate102inter8));
  nand2 gate1900(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1901(.a(s_193), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1902(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1903(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1904(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate771(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate772(.a(gate105inter0), .b(s_32), .O(gate105inter1));
  and2  gate773(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate774(.a(s_32), .O(gate105inter3));
  inv1  gate775(.a(s_33), .O(gate105inter4));
  nand2 gate776(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate777(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate778(.a(G362), .O(gate105inter7));
  inv1  gate779(.a(G363), .O(gate105inter8));
  nand2 gate780(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate781(.a(s_33), .b(gate105inter3), .O(gate105inter10));
  nor2  gate782(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate783(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate784(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate673(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate674(.a(gate106inter0), .b(s_18), .O(gate106inter1));
  and2  gate675(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate676(.a(s_18), .O(gate106inter3));
  inv1  gate677(.a(s_19), .O(gate106inter4));
  nand2 gate678(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate679(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate680(.a(G364), .O(gate106inter7));
  inv1  gate681(.a(G365), .O(gate106inter8));
  nand2 gate682(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate683(.a(s_19), .b(gate106inter3), .O(gate106inter10));
  nor2  gate684(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate685(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate686(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1639(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1640(.a(gate107inter0), .b(s_156), .O(gate107inter1));
  and2  gate1641(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1642(.a(s_156), .O(gate107inter3));
  inv1  gate1643(.a(s_157), .O(gate107inter4));
  nand2 gate1644(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1645(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1646(.a(G366), .O(gate107inter7));
  inv1  gate1647(.a(G367), .O(gate107inter8));
  nand2 gate1648(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1649(.a(s_157), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1650(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1651(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1652(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate2073(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2074(.a(gate112inter0), .b(s_218), .O(gate112inter1));
  and2  gate2075(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2076(.a(s_218), .O(gate112inter3));
  inv1  gate2077(.a(s_219), .O(gate112inter4));
  nand2 gate2078(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2079(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2080(.a(G376), .O(gate112inter7));
  inv1  gate2081(.a(G377), .O(gate112inter8));
  nand2 gate2082(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2083(.a(s_219), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2084(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2085(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2086(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2283(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2284(.a(gate115inter0), .b(s_248), .O(gate115inter1));
  and2  gate2285(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2286(.a(s_248), .O(gate115inter3));
  inv1  gate2287(.a(s_249), .O(gate115inter4));
  nand2 gate2288(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2289(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2290(.a(G382), .O(gate115inter7));
  inv1  gate2291(.a(G383), .O(gate115inter8));
  nand2 gate2292(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2293(.a(s_249), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2294(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2295(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2296(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate589(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate590(.a(gate117inter0), .b(s_6), .O(gate117inter1));
  and2  gate591(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate592(.a(s_6), .O(gate117inter3));
  inv1  gate593(.a(s_7), .O(gate117inter4));
  nand2 gate594(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate595(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate596(.a(G386), .O(gate117inter7));
  inv1  gate597(.a(G387), .O(gate117inter8));
  nand2 gate598(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate599(.a(s_7), .b(gate117inter3), .O(gate117inter10));
  nor2  gate600(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate601(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate602(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1107(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1108(.a(gate124inter0), .b(s_80), .O(gate124inter1));
  and2  gate1109(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1110(.a(s_80), .O(gate124inter3));
  inv1  gate1111(.a(s_81), .O(gate124inter4));
  nand2 gate1112(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1113(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1114(.a(G400), .O(gate124inter7));
  inv1  gate1115(.a(G401), .O(gate124inter8));
  nand2 gate1116(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1117(.a(s_81), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1118(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1119(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1120(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1023(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1024(.a(gate125inter0), .b(s_68), .O(gate125inter1));
  and2  gate1025(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1026(.a(s_68), .O(gate125inter3));
  inv1  gate1027(.a(s_69), .O(gate125inter4));
  nand2 gate1028(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1029(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1030(.a(G402), .O(gate125inter7));
  inv1  gate1031(.a(G403), .O(gate125inter8));
  nand2 gate1032(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1033(.a(s_69), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1034(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1035(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1036(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate701(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate702(.a(gate135inter0), .b(s_22), .O(gate135inter1));
  and2  gate703(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate704(.a(s_22), .O(gate135inter3));
  inv1  gate705(.a(s_23), .O(gate135inter4));
  nand2 gate706(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate707(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate708(.a(G422), .O(gate135inter7));
  inv1  gate709(.a(G423), .O(gate135inter8));
  nand2 gate710(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate711(.a(s_23), .b(gate135inter3), .O(gate135inter10));
  nor2  gate712(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate713(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate714(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1163(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1164(.a(gate136inter0), .b(s_88), .O(gate136inter1));
  and2  gate1165(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1166(.a(s_88), .O(gate136inter3));
  inv1  gate1167(.a(s_89), .O(gate136inter4));
  nand2 gate1168(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1169(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1170(.a(G424), .O(gate136inter7));
  inv1  gate1171(.a(G425), .O(gate136inter8));
  nand2 gate1172(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1173(.a(s_89), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1174(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1175(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1176(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate561(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate562(.a(gate139inter0), .b(s_2), .O(gate139inter1));
  and2  gate563(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate564(.a(s_2), .O(gate139inter3));
  inv1  gate565(.a(s_3), .O(gate139inter4));
  nand2 gate566(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate567(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate568(.a(G438), .O(gate139inter7));
  inv1  gate569(.a(G441), .O(gate139inter8));
  nand2 gate570(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate571(.a(s_3), .b(gate139inter3), .O(gate139inter10));
  nor2  gate572(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate573(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate574(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate631(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate632(.a(gate142inter0), .b(s_12), .O(gate142inter1));
  and2  gate633(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate634(.a(s_12), .O(gate142inter3));
  inv1  gate635(.a(s_13), .O(gate142inter4));
  nand2 gate636(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate637(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate638(.a(G456), .O(gate142inter7));
  inv1  gate639(.a(G459), .O(gate142inter8));
  nand2 gate640(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate641(.a(s_13), .b(gate142inter3), .O(gate142inter10));
  nor2  gate642(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate643(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate644(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1051(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1052(.a(gate150inter0), .b(s_72), .O(gate150inter1));
  and2  gate1053(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1054(.a(s_72), .O(gate150inter3));
  inv1  gate1055(.a(s_73), .O(gate150inter4));
  nand2 gate1056(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1057(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1058(.a(G504), .O(gate150inter7));
  inv1  gate1059(.a(G507), .O(gate150inter8));
  nand2 gate1060(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1061(.a(s_73), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1062(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1063(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1064(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1065(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1066(.a(gate154inter0), .b(s_74), .O(gate154inter1));
  and2  gate1067(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1068(.a(s_74), .O(gate154inter3));
  inv1  gate1069(.a(s_75), .O(gate154inter4));
  nand2 gate1070(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1071(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1072(.a(G429), .O(gate154inter7));
  inv1  gate1073(.a(G522), .O(gate154inter8));
  nand2 gate1074(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1075(.a(s_75), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1076(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1077(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1078(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate981(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate982(.a(gate155inter0), .b(s_62), .O(gate155inter1));
  and2  gate983(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate984(.a(s_62), .O(gate155inter3));
  inv1  gate985(.a(s_63), .O(gate155inter4));
  nand2 gate986(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate987(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate988(.a(G432), .O(gate155inter7));
  inv1  gate989(.a(G525), .O(gate155inter8));
  nand2 gate990(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate991(.a(s_63), .b(gate155inter3), .O(gate155inter10));
  nor2  gate992(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate993(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate994(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1037(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1038(.a(gate160inter0), .b(s_70), .O(gate160inter1));
  and2  gate1039(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1040(.a(s_70), .O(gate160inter3));
  inv1  gate1041(.a(s_71), .O(gate160inter4));
  nand2 gate1042(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1043(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1044(.a(G447), .O(gate160inter7));
  inv1  gate1045(.a(G531), .O(gate160inter8));
  nand2 gate1046(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1047(.a(s_71), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1048(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1049(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1050(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2269(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2270(.a(gate170inter0), .b(s_246), .O(gate170inter1));
  and2  gate2271(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2272(.a(s_246), .O(gate170inter3));
  inv1  gate2273(.a(s_247), .O(gate170inter4));
  nand2 gate2274(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2275(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2276(.a(G477), .O(gate170inter7));
  inv1  gate2277(.a(G546), .O(gate170inter8));
  nand2 gate2278(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2279(.a(s_247), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2280(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2281(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2282(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1751(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1752(.a(gate180inter0), .b(s_172), .O(gate180inter1));
  and2  gate1753(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1754(.a(s_172), .O(gate180inter3));
  inv1  gate1755(.a(s_173), .O(gate180inter4));
  nand2 gate1756(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1757(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1758(.a(G507), .O(gate180inter7));
  inv1  gate1759(.a(G561), .O(gate180inter8));
  nand2 gate1760(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1761(.a(s_173), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1762(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1763(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1764(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1737(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1738(.a(gate182inter0), .b(s_170), .O(gate182inter1));
  and2  gate1739(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1740(.a(s_170), .O(gate182inter3));
  inv1  gate1741(.a(s_171), .O(gate182inter4));
  nand2 gate1742(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1743(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1744(.a(G513), .O(gate182inter7));
  inv1  gate1745(.a(G564), .O(gate182inter8));
  nand2 gate1746(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1747(.a(s_171), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1748(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1749(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1750(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate659(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate660(.a(gate188inter0), .b(s_16), .O(gate188inter1));
  and2  gate661(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate662(.a(s_16), .O(gate188inter3));
  inv1  gate663(.a(s_17), .O(gate188inter4));
  nand2 gate664(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate665(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate666(.a(G576), .O(gate188inter7));
  inv1  gate667(.a(G577), .O(gate188inter8));
  nand2 gate668(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate669(.a(s_17), .b(gate188inter3), .O(gate188inter10));
  nor2  gate670(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate671(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate672(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1877(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1878(.a(gate192inter0), .b(s_190), .O(gate192inter1));
  and2  gate1879(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1880(.a(s_190), .O(gate192inter3));
  inv1  gate1881(.a(s_191), .O(gate192inter4));
  nand2 gate1882(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1883(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1884(.a(G584), .O(gate192inter7));
  inv1  gate1885(.a(G585), .O(gate192inter8));
  nand2 gate1886(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1887(.a(s_191), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1888(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1889(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1890(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2115(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2116(.a(gate193inter0), .b(s_224), .O(gate193inter1));
  and2  gate2117(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2118(.a(s_224), .O(gate193inter3));
  inv1  gate2119(.a(s_225), .O(gate193inter4));
  nand2 gate2120(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2121(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2122(.a(G586), .O(gate193inter7));
  inv1  gate2123(.a(G587), .O(gate193inter8));
  nand2 gate2124(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2125(.a(s_225), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2126(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2127(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2128(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate2199(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2200(.a(gate196inter0), .b(s_236), .O(gate196inter1));
  and2  gate2201(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2202(.a(s_236), .O(gate196inter3));
  inv1  gate2203(.a(s_237), .O(gate196inter4));
  nand2 gate2204(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2205(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2206(.a(G592), .O(gate196inter7));
  inv1  gate2207(.a(G593), .O(gate196inter8));
  nand2 gate2208(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2209(.a(s_237), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2210(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2211(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2212(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1849(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1850(.a(gate199inter0), .b(s_186), .O(gate199inter1));
  and2  gate1851(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1852(.a(s_186), .O(gate199inter3));
  inv1  gate1853(.a(s_187), .O(gate199inter4));
  nand2 gate1854(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1855(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1856(.a(G598), .O(gate199inter7));
  inv1  gate1857(.a(G599), .O(gate199inter8));
  nand2 gate1858(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1859(.a(s_187), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1860(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1861(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1862(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1219(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1220(.a(gate200inter0), .b(s_96), .O(gate200inter1));
  and2  gate1221(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1222(.a(s_96), .O(gate200inter3));
  inv1  gate1223(.a(s_97), .O(gate200inter4));
  nand2 gate1224(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1225(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1226(.a(G600), .O(gate200inter7));
  inv1  gate1227(.a(G601), .O(gate200inter8));
  nand2 gate1228(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1229(.a(s_97), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1230(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1231(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1232(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate967(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate968(.a(gate202inter0), .b(s_60), .O(gate202inter1));
  and2  gate969(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate970(.a(s_60), .O(gate202inter3));
  inv1  gate971(.a(s_61), .O(gate202inter4));
  nand2 gate972(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate973(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate974(.a(G612), .O(gate202inter7));
  inv1  gate975(.a(G617), .O(gate202inter8));
  nand2 gate976(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate977(.a(s_61), .b(gate202inter3), .O(gate202inter10));
  nor2  gate978(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate979(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate980(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1695(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1696(.a(gate203inter0), .b(s_164), .O(gate203inter1));
  and2  gate1697(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1698(.a(s_164), .O(gate203inter3));
  inv1  gate1699(.a(s_165), .O(gate203inter4));
  nand2 gate1700(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1701(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1702(.a(G602), .O(gate203inter7));
  inv1  gate1703(.a(G612), .O(gate203inter8));
  nand2 gate1704(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1705(.a(s_165), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1706(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1707(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1708(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1555(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1556(.a(gate206inter0), .b(s_144), .O(gate206inter1));
  and2  gate1557(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1558(.a(s_144), .O(gate206inter3));
  inv1  gate1559(.a(s_145), .O(gate206inter4));
  nand2 gate1560(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1561(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1562(.a(G632), .O(gate206inter7));
  inv1  gate1563(.a(G637), .O(gate206inter8));
  nand2 gate1564(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1565(.a(s_145), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1566(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1567(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1568(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1835(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1836(.a(gate207inter0), .b(s_184), .O(gate207inter1));
  and2  gate1837(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1838(.a(s_184), .O(gate207inter3));
  inv1  gate1839(.a(s_185), .O(gate207inter4));
  nand2 gate1840(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1841(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1842(.a(G622), .O(gate207inter7));
  inv1  gate1843(.a(G632), .O(gate207inter8));
  nand2 gate1844(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1845(.a(s_185), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1846(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1847(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1848(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1905(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1906(.a(gate211inter0), .b(s_194), .O(gate211inter1));
  and2  gate1907(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1908(.a(s_194), .O(gate211inter3));
  inv1  gate1909(.a(s_195), .O(gate211inter4));
  nand2 gate1910(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1911(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1912(.a(G612), .O(gate211inter7));
  inv1  gate1913(.a(G669), .O(gate211inter8));
  nand2 gate1914(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1915(.a(s_195), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1916(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1917(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1918(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2367(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2368(.a(gate216inter0), .b(s_260), .O(gate216inter1));
  and2  gate2369(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2370(.a(s_260), .O(gate216inter3));
  inv1  gate2371(.a(s_261), .O(gate216inter4));
  nand2 gate2372(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2373(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2374(.a(G617), .O(gate216inter7));
  inv1  gate2375(.a(G675), .O(gate216inter8));
  nand2 gate2376(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2377(.a(s_261), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2378(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2379(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2380(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate729(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate730(.a(gate219inter0), .b(s_26), .O(gate219inter1));
  and2  gate731(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate732(.a(s_26), .O(gate219inter3));
  inv1  gate733(.a(s_27), .O(gate219inter4));
  nand2 gate734(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate735(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate736(.a(G632), .O(gate219inter7));
  inv1  gate737(.a(G681), .O(gate219inter8));
  nand2 gate738(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate739(.a(s_27), .b(gate219inter3), .O(gate219inter10));
  nor2  gate740(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate741(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate742(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate687(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate688(.a(gate220inter0), .b(s_20), .O(gate220inter1));
  and2  gate689(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate690(.a(s_20), .O(gate220inter3));
  inv1  gate691(.a(s_21), .O(gate220inter4));
  nand2 gate692(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate693(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate694(.a(G637), .O(gate220inter7));
  inv1  gate695(.a(G681), .O(gate220inter8));
  nand2 gate696(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate697(.a(s_21), .b(gate220inter3), .O(gate220inter10));
  nor2  gate698(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate699(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate700(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate617(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate618(.a(gate222inter0), .b(s_10), .O(gate222inter1));
  and2  gate619(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate620(.a(s_10), .O(gate222inter3));
  inv1  gate621(.a(s_11), .O(gate222inter4));
  nand2 gate622(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate623(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate624(.a(G632), .O(gate222inter7));
  inv1  gate625(.a(G684), .O(gate222inter8));
  nand2 gate626(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate627(.a(s_11), .b(gate222inter3), .O(gate222inter10));
  nor2  gate628(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate629(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate630(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1807(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1808(.a(gate229inter0), .b(s_180), .O(gate229inter1));
  and2  gate1809(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1810(.a(s_180), .O(gate229inter3));
  inv1  gate1811(.a(s_181), .O(gate229inter4));
  nand2 gate1812(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1813(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1814(.a(G698), .O(gate229inter7));
  inv1  gate1815(.a(G699), .O(gate229inter8));
  nand2 gate1816(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1817(.a(s_181), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1818(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1819(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1820(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1989(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1990(.a(gate236inter0), .b(s_206), .O(gate236inter1));
  and2  gate1991(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1992(.a(s_206), .O(gate236inter3));
  inv1  gate1993(.a(s_207), .O(gate236inter4));
  nand2 gate1994(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1995(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1996(.a(G251), .O(gate236inter7));
  inv1  gate1997(.a(G727), .O(gate236inter8));
  nand2 gate1998(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1999(.a(s_207), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2000(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2001(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2002(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1583(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1584(.a(gate240inter0), .b(s_148), .O(gate240inter1));
  and2  gate1585(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1586(.a(s_148), .O(gate240inter3));
  inv1  gate1587(.a(s_149), .O(gate240inter4));
  nand2 gate1588(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1589(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1590(.a(G263), .O(gate240inter7));
  inv1  gate1591(.a(G715), .O(gate240inter8));
  nand2 gate1592(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1593(.a(s_149), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1594(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1595(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1596(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate953(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate954(.a(gate243inter0), .b(s_58), .O(gate243inter1));
  and2  gate955(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate956(.a(s_58), .O(gate243inter3));
  inv1  gate957(.a(s_59), .O(gate243inter4));
  nand2 gate958(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate959(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate960(.a(G245), .O(gate243inter7));
  inv1  gate961(.a(G733), .O(gate243inter8));
  nand2 gate962(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate963(.a(s_59), .b(gate243inter3), .O(gate243inter10));
  nor2  gate964(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate965(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate966(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate897(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate898(.a(gate244inter0), .b(s_50), .O(gate244inter1));
  and2  gate899(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate900(.a(s_50), .O(gate244inter3));
  inv1  gate901(.a(s_51), .O(gate244inter4));
  nand2 gate902(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate903(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate904(.a(G721), .O(gate244inter7));
  inv1  gate905(.a(G733), .O(gate244inter8));
  nand2 gate906(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate907(.a(s_51), .b(gate244inter3), .O(gate244inter10));
  nor2  gate908(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate909(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate910(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1541(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1542(.a(gate246inter0), .b(s_142), .O(gate246inter1));
  and2  gate1543(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1544(.a(s_142), .O(gate246inter3));
  inv1  gate1545(.a(s_143), .O(gate246inter4));
  nand2 gate1546(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1547(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1548(.a(G724), .O(gate246inter7));
  inv1  gate1549(.a(G736), .O(gate246inter8));
  nand2 gate1550(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1551(.a(s_143), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1552(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1553(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1554(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2003(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2004(.a(gate249inter0), .b(s_208), .O(gate249inter1));
  and2  gate2005(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2006(.a(s_208), .O(gate249inter3));
  inv1  gate2007(.a(s_209), .O(gate249inter4));
  nand2 gate2008(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2009(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2010(.a(G254), .O(gate249inter7));
  inv1  gate2011(.a(G742), .O(gate249inter8));
  nand2 gate2012(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2013(.a(s_209), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2014(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2015(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2016(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1933(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1934(.a(gate250inter0), .b(s_198), .O(gate250inter1));
  and2  gate1935(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1936(.a(s_198), .O(gate250inter3));
  inv1  gate1937(.a(s_199), .O(gate250inter4));
  nand2 gate1938(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1939(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1940(.a(G706), .O(gate250inter7));
  inv1  gate1941(.a(G742), .O(gate250inter8));
  nand2 gate1942(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1943(.a(s_199), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1944(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1945(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1946(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1709(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1710(.a(gate252inter0), .b(s_166), .O(gate252inter1));
  and2  gate1711(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1712(.a(s_166), .O(gate252inter3));
  inv1  gate1713(.a(s_167), .O(gate252inter4));
  nand2 gate1714(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1715(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1716(.a(G709), .O(gate252inter7));
  inv1  gate1717(.a(G745), .O(gate252inter8));
  nand2 gate1718(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1719(.a(s_167), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1720(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1721(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1722(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1975(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1976(.a(gate257inter0), .b(s_204), .O(gate257inter1));
  and2  gate1977(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1978(.a(s_204), .O(gate257inter3));
  inv1  gate1979(.a(s_205), .O(gate257inter4));
  nand2 gate1980(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1981(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1982(.a(G754), .O(gate257inter7));
  inv1  gate1983(.a(G755), .O(gate257inter8));
  nand2 gate1984(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1985(.a(s_205), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1986(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1987(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1988(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate2339(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2340(.a(gate260inter0), .b(s_256), .O(gate260inter1));
  and2  gate2341(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2342(.a(s_256), .O(gate260inter3));
  inv1  gate2343(.a(s_257), .O(gate260inter4));
  nand2 gate2344(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2345(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2346(.a(G760), .O(gate260inter7));
  inv1  gate2347(.a(G761), .O(gate260inter8));
  nand2 gate2348(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2349(.a(s_257), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2350(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2351(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2352(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2157(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2158(.a(gate263inter0), .b(s_230), .O(gate263inter1));
  and2  gate2159(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2160(.a(s_230), .O(gate263inter3));
  inv1  gate2161(.a(s_231), .O(gate263inter4));
  nand2 gate2162(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2163(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2164(.a(G766), .O(gate263inter7));
  inv1  gate2165(.a(G767), .O(gate263inter8));
  nand2 gate2166(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2167(.a(s_231), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2168(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2169(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2170(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1149(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1150(.a(gate264inter0), .b(s_86), .O(gate264inter1));
  and2  gate1151(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1152(.a(s_86), .O(gate264inter3));
  inv1  gate1153(.a(s_87), .O(gate264inter4));
  nand2 gate1154(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1155(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1156(.a(G768), .O(gate264inter7));
  inv1  gate1157(.a(G769), .O(gate264inter8));
  nand2 gate1158(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1159(.a(s_87), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1160(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1161(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1162(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1317(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1318(.a(gate265inter0), .b(s_110), .O(gate265inter1));
  and2  gate1319(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1320(.a(s_110), .O(gate265inter3));
  inv1  gate1321(.a(s_111), .O(gate265inter4));
  nand2 gate1322(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1323(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1324(.a(G642), .O(gate265inter7));
  inv1  gate1325(.a(G770), .O(gate265inter8));
  nand2 gate1326(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1327(.a(s_111), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1328(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1329(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1330(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1681(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1682(.a(gate269inter0), .b(s_162), .O(gate269inter1));
  and2  gate1683(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1684(.a(s_162), .O(gate269inter3));
  inv1  gate1685(.a(s_163), .O(gate269inter4));
  nand2 gate1686(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1687(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1688(.a(G654), .O(gate269inter7));
  inv1  gate1689(.a(G782), .O(gate269inter8));
  nand2 gate1690(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1691(.a(s_163), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1692(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1693(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1694(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2311(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2312(.a(gate271inter0), .b(s_252), .O(gate271inter1));
  and2  gate2313(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2314(.a(s_252), .O(gate271inter3));
  inv1  gate2315(.a(s_253), .O(gate271inter4));
  nand2 gate2316(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2317(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2318(.a(G660), .O(gate271inter7));
  inv1  gate2319(.a(G788), .O(gate271inter8));
  nand2 gate2320(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2321(.a(s_253), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2322(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2323(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2324(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1653(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1654(.a(gate274inter0), .b(s_158), .O(gate274inter1));
  and2  gate1655(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1656(.a(s_158), .O(gate274inter3));
  inv1  gate1657(.a(s_159), .O(gate274inter4));
  nand2 gate1658(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1659(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1660(.a(G770), .O(gate274inter7));
  inv1  gate1661(.a(G794), .O(gate274inter8));
  nand2 gate1662(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1663(.a(s_159), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1664(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1665(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1666(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2129(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2130(.a(gate278inter0), .b(s_226), .O(gate278inter1));
  and2  gate2131(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2132(.a(s_226), .O(gate278inter3));
  inv1  gate2133(.a(s_227), .O(gate278inter4));
  nand2 gate2134(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2135(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2136(.a(G776), .O(gate278inter7));
  inv1  gate2137(.a(G800), .O(gate278inter8));
  nand2 gate2138(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2139(.a(s_227), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2140(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2141(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2142(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2017(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2018(.a(gate285inter0), .b(s_210), .O(gate285inter1));
  and2  gate2019(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2020(.a(s_210), .O(gate285inter3));
  inv1  gate2021(.a(s_211), .O(gate285inter4));
  nand2 gate2022(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2023(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2024(.a(G660), .O(gate285inter7));
  inv1  gate2025(.a(G812), .O(gate285inter8));
  nand2 gate2026(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2027(.a(s_211), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2028(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2029(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2030(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2353(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2354(.a(gate287inter0), .b(s_258), .O(gate287inter1));
  and2  gate2355(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2356(.a(s_258), .O(gate287inter3));
  inv1  gate2357(.a(s_259), .O(gate287inter4));
  nand2 gate2358(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2359(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2360(.a(G663), .O(gate287inter7));
  inv1  gate2361(.a(G815), .O(gate287inter8));
  nand2 gate2362(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2363(.a(s_259), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2364(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2365(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2366(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2087(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2088(.a(gate292inter0), .b(s_220), .O(gate292inter1));
  and2  gate2089(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2090(.a(s_220), .O(gate292inter3));
  inv1  gate2091(.a(s_221), .O(gate292inter4));
  nand2 gate2092(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2093(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2094(.a(G824), .O(gate292inter7));
  inv1  gate2095(.a(G825), .O(gate292inter8));
  nand2 gate2096(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2097(.a(s_221), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2098(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2099(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2100(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1569(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1570(.a(gate294inter0), .b(s_146), .O(gate294inter1));
  and2  gate1571(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1572(.a(s_146), .O(gate294inter3));
  inv1  gate1573(.a(s_147), .O(gate294inter4));
  nand2 gate1574(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1575(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1576(.a(G832), .O(gate294inter7));
  inv1  gate1577(.a(G833), .O(gate294inter8));
  nand2 gate1578(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1579(.a(s_147), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1580(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1581(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1582(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1779(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1780(.a(gate296inter0), .b(s_176), .O(gate296inter1));
  and2  gate1781(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1782(.a(s_176), .O(gate296inter3));
  inv1  gate1783(.a(s_177), .O(gate296inter4));
  nand2 gate1784(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1785(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1786(.a(G826), .O(gate296inter7));
  inv1  gate1787(.a(G827), .O(gate296inter8));
  nand2 gate1788(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1789(.a(s_177), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1790(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1791(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1792(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1485(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1486(.a(gate387inter0), .b(s_134), .O(gate387inter1));
  and2  gate1487(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1488(.a(s_134), .O(gate387inter3));
  inv1  gate1489(.a(s_135), .O(gate387inter4));
  nand2 gate1490(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1491(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1492(.a(G1), .O(gate387inter7));
  inv1  gate1493(.a(G1036), .O(gate387inter8));
  nand2 gate1494(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1495(.a(s_135), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1496(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1497(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1498(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate799(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate800(.a(gate395inter0), .b(s_36), .O(gate395inter1));
  and2  gate801(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate802(.a(s_36), .O(gate395inter3));
  inv1  gate803(.a(s_37), .O(gate395inter4));
  nand2 gate804(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate805(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate806(.a(G9), .O(gate395inter7));
  inv1  gate807(.a(G1060), .O(gate395inter8));
  nand2 gate808(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate809(.a(s_37), .b(gate395inter3), .O(gate395inter10));
  nor2  gate810(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate811(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate812(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1205(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1206(.a(gate398inter0), .b(s_94), .O(gate398inter1));
  and2  gate1207(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1208(.a(s_94), .O(gate398inter3));
  inv1  gate1209(.a(s_95), .O(gate398inter4));
  nand2 gate1210(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1211(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1212(.a(G12), .O(gate398inter7));
  inv1  gate1213(.a(G1069), .O(gate398inter8));
  nand2 gate1214(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1215(.a(s_95), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1216(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1217(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1218(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate911(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate912(.a(gate401inter0), .b(s_52), .O(gate401inter1));
  and2  gate913(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate914(.a(s_52), .O(gate401inter3));
  inv1  gate915(.a(s_53), .O(gate401inter4));
  nand2 gate916(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate917(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate918(.a(G15), .O(gate401inter7));
  inv1  gate919(.a(G1078), .O(gate401inter8));
  nand2 gate920(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate921(.a(s_53), .b(gate401inter3), .O(gate401inter10));
  nor2  gate922(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate923(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate924(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate1597(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1598(.a(gate402inter0), .b(s_150), .O(gate402inter1));
  and2  gate1599(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1600(.a(s_150), .O(gate402inter3));
  inv1  gate1601(.a(s_151), .O(gate402inter4));
  nand2 gate1602(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1603(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1604(.a(G16), .O(gate402inter7));
  inv1  gate1605(.a(G1081), .O(gate402inter8));
  nand2 gate1606(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1607(.a(s_151), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1608(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1609(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1610(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate547(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate548(.a(gate404inter0), .b(s_0), .O(gate404inter1));
  and2  gate549(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate550(.a(s_0), .O(gate404inter3));
  inv1  gate551(.a(s_1), .O(gate404inter4));
  nand2 gate552(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate553(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate554(.a(G18), .O(gate404inter7));
  inv1  gate555(.a(G1087), .O(gate404inter8));
  nand2 gate556(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate557(.a(s_1), .b(gate404inter3), .O(gate404inter10));
  nor2  gate558(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate559(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate560(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1177(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1178(.a(gate407inter0), .b(s_90), .O(gate407inter1));
  and2  gate1179(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1180(.a(s_90), .O(gate407inter3));
  inv1  gate1181(.a(s_91), .O(gate407inter4));
  nand2 gate1182(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1183(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1184(.a(G21), .O(gate407inter7));
  inv1  gate1185(.a(G1096), .O(gate407inter8));
  nand2 gate1186(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1187(.a(s_91), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1188(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1189(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1190(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1247(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1248(.a(gate411inter0), .b(s_100), .O(gate411inter1));
  and2  gate1249(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1250(.a(s_100), .O(gate411inter3));
  inv1  gate1251(.a(s_101), .O(gate411inter4));
  nand2 gate1252(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1253(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1254(.a(G25), .O(gate411inter7));
  inv1  gate1255(.a(G1108), .O(gate411inter8));
  nand2 gate1256(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1257(.a(s_101), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1258(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1259(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1260(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1233(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1234(.a(gate412inter0), .b(s_98), .O(gate412inter1));
  and2  gate1235(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1236(.a(s_98), .O(gate412inter3));
  inv1  gate1237(.a(s_99), .O(gate412inter4));
  nand2 gate1238(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1239(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1240(.a(G26), .O(gate412inter7));
  inv1  gate1241(.a(G1111), .O(gate412inter8));
  nand2 gate1242(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1243(.a(s_99), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1244(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1245(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1246(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate2241(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2242(.a(gate413inter0), .b(s_242), .O(gate413inter1));
  and2  gate2243(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2244(.a(s_242), .O(gate413inter3));
  inv1  gate2245(.a(s_243), .O(gate413inter4));
  nand2 gate2246(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2247(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2248(.a(G27), .O(gate413inter7));
  inv1  gate2249(.a(G1114), .O(gate413inter8));
  nand2 gate2250(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2251(.a(s_243), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2252(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2253(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2254(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1961(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1962(.a(gate426inter0), .b(s_202), .O(gate426inter1));
  and2  gate1963(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1964(.a(s_202), .O(gate426inter3));
  inv1  gate1965(.a(s_203), .O(gate426inter4));
  nand2 gate1966(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1967(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1968(.a(G1045), .O(gate426inter7));
  inv1  gate1969(.a(G1141), .O(gate426inter8));
  nand2 gate1970(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1971(.a(s_203), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1972(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1973(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1974(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1947(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1948(.a(gate427inter0), .b(s_200), .O(gate427inter1));
  and2  gate1949(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1950(.a(s_200), .O(gate427inter3));
  inv1  gate1951(.a(s_201), .O(gate427inter4));
  nand2 gate1952(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1953(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1954(.a(G5), .O(gate427inter7));
  inv1  gate1955(.a(G1144), .O(gate427inter8));
  nand2 gate1956(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1957(.a(s_201), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1958(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1959(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1960(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1821(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1822(.a(gate429inter0), .b(s_182), .O(gate429inter1));
  and2  gate1823(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1824(.a(s_182), .O(gate429inter3));
  inv1  gate1825(.a(s_183), .O(gate429inter4));
  nand2 gate1826(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1827(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1828(.a(G6), .O(gate429inter7));
  inv1  gate1829(.a(G1147), .O(gate429inter8));
  nand2 gate1830(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1831(.a(s_183), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1832(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1833(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1834(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate757(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate758(.a(gate430inter0), .b(s_30), .O(gate430inter1));
  and2  gate759(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate760(.a(s_30), .O(gate430inter3));
  inv1  gate761(.a(s_31), .O(gate430inter4));
  nand2 gate762(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate763(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate764(.a(G1051), .O(gate430inter7));
  inv1  gate765(.a(G1147), .O(gate430inter8));
  nand2 gate766(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate767(.a(s_31), .b(gate430inter3), .O(gate430inter10));
  nor2  gate768(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate769(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate770(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1303(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1304(.a(gate432inter0), .b(s_108), .O(gate432inter1));
  and2  gate1305(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1306(.a(s_108), .O(gate432inter3));
  inv1  gate1307(.a(s_109), .O(gate432inter4));
  nand2 gate1308(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1309(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1310(.a(G1054), .O(gate432inter7));
  inv1  gate1311(.a(G1150), .O(gate432inter8));
  nand2 gate1312(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1313(.a(s_109), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1314(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1315(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1316(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate925(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate926(.a(gate434inter0), .b(s_54), .O(gate434inter1));
  and2  gate927(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate928(.a(s_54), .O(gate434inter3));
  inv1  gate929(.a(s_55), .O(gate434inter4));
  nand2 gate930(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate931(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate932(.a(G1057), .O(gate434inter7));
  inv1  gate933(.a(G1153), .O(gate434inter8));
  nand2 gate934(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate935(.a(s_55), .b(gate434inter3), .O(gate434inter10));
  nor2  gate936(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate937(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate938(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate575(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate576(.a(gate440inter0), .b(s_4), .O(gate440inter1));
  and2  gate577(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate578(.a(s_4), .O(gate440inter3));
  inv1  gate579(.a(s_5), .O(gate440inter4));
  nand2 gate580(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate581(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate582(.a(G1066), .O(gate440inter7));
  inv1  gate583(.a(G1162), .O(gate440inter8));
  nand2 gate584(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate585(.a(s_5), .b(gate440inter3), .O(gate440inter10));
  nor2  gate586(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate587(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate588(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1415(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1416(.a(gate443inter0), .b(s_124), .O(gate443inter1));
  and2  gate1417(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1418(.a(s_124), .O(gate443inter3));
  inv1  gate1419(.a(s_125), .O(gate443inter4));
  nand2 gate1420(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1421(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1422(.a(G13), .O(gate443inter7));
  inv1  gate1423(.a(G1168), .O(gate443inter8));
  nand2 gate1424(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1425(.a(s_125), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1426(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1427(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1428(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1261(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1262(.a(gate445inter0), .b(s_102), .O(gate445inter1));
  and2  gate1263(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1264(.a(s_102), .O(gate445inter3));
  inv1  gate1265(.a(s_103), .O(gate445inter4));
  nand2 gate1266(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1267(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1268(.a(G14), .O(gate445inter7));
  inv1  gate1269(.a(G1171), .O(gate445inter8));
  nand2 gate1270(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1271(.a(s_103), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1272(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1273(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1274(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1457(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1458(.a(gate446inter0), .b(s_130), .O(gate446inter1));
  and2  gate1459(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1460(.a(s_130), .O(gate446inter3));
  inv1  gate1461(.a(s_131), .O(gate446inter4));
  nand2 gate1462(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1463(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1464(.a(G1075), .O(gate446inter7));
  inv1  gate1465(.a(G1171), .O(gate446inter8));
  nand2 gate1466(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1467(.a(s_131), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1468(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1469(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1470(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate939(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate940(.a(gate447inter0), .b(s_56), .O(gate447inter1));
  and2  gate941(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate942(.a(s_56), .O(gate447inter3));
  inv1  gate943(.a(s_57), .O(gate447inter4));
  nand2 gate944(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate945(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate946(.a(G15), .O(gate447inter7));
  inv1  gate947(.a(G1174), .O(gate447inter8));
  nand2 gate948(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate949(.a(s_57), .b(gate447inter3), .O(gate447inter10));
  nor2  gate950(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate951(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate952(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate841(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate842(.a(gate449inter0), .b(s_42), .O(gate449inter1));
  and2  gate843(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate844(.a(s_42), .O(gate449inter3));
  inv1  gate845(.a(s_43), .O(gate449inter4));
  nand2 gate846(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate847(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate848(.a(G16), .O(gate449inter7));
  inv1  gate849(.a(G1177), .O(gate449inter8));
  nand2 gate850(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate851(.a(s_43), .b(gate449inter3), .O(gate449inter10));
  nor2  gate852(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate853(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate854(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1919(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1920(.a(gate450inter0), .b(s_196), .O(gate450inter1));
  and2  gate1921(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1922(.a(s_196), .O(gate450inter3));
  inv1  gate1923(.a(s_197), .O(gate450inter4));
  nand2 gate1924(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1925(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1926(.a(G1081), .O(gate450inter7));
  inv1  gate1927(.a(G1177), .O(gate450inter8));
  nand2 gate1928(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1929(.a(s_197), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1930(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1931(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1932(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2143(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2144(.a(gate454inter0), .b(s_228), .O(gate454inter1));
  and2  gate2145(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2146(.a(s_228), .O(gate454inter3));
  inv1  gate2147(.a(s_229), .O(gate454inter4));
  nand2 gate2148(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2149(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2150(.a(G1087), .O(gate454inter7));
  inv1  gate2151(.a(G1183), .O(gate454inter8));
  nand2 gate2152(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2153(.a(s_229), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2154(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2155(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2156(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1289(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1290(.a(gate455inter0), .b(s_106), .O(gate455inter1));
  and2  gate1291(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1292(.a(s_106), .O(gate455inter3));
  inv1  gate1293(.a(s_107), .O(gate455inter4));
  nand2 gate1294(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1295(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1296(.a(G19), .O(gate455inter7));
  inv1  gate1297(.a(G1186), .O(gate455inter8));
  nand2 gate1298(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1299(.a(s_107), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1300(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1301(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1302(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2185(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2186(.a(gate458inter0), .b(s_234), .O(gate458inter1));
  and2  gate2187(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2188(.a(s_234), .O(gate458inter3));
  inv1  gate2189(.a(s_235), .O(gate458inter4));
  nand2 gate2190(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2191(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2192(.a(G1093), .O(gate458inter7));
  inv1  gate2193(.a(G1189), .O(gate458inter8));
  nand2 gate2194(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2195(.a(s_235), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2196(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2197(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2198(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1625(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1626(.a(gate459inter0), .b(s_154), .O(gate459inter1));
  and2  gate1627(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1628(.a(s_154), .O(gate459inter3));
  inv1  gate1629(.a(s_155), .O(gate459inter4));
  nand2 gate1630(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1631(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1632(.a(G21), .O(gate459inter7));
  inv1  gate1633(.a(G1192), .O(gate459inter8));
  nand2 gate1634(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1635(.a(s_155), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1636(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1637(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1638(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1093(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1094(.a(gate460inter0), .b(s_78), .O(gate460inter1));
  and2  gate1095(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1096(.a(s_78), .O(gate460inter3));
  inv1  gate1097(.a(s_79), .O(gate460inter4));
  nand2 gate1098(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1099(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1100(.a(G1096), .O(gate460inter7));
  inv1  gate1101(.a(G1192), .O(gate460inter8));
  nand2 gate1102(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1103(.a(s_79), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1104(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1105(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1106(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate869(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate870(.a(gate463inter0), .b(s_46), .O(gate463inter1));
  and2  gate871(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate872(.a(s_46), .O(gate463inter3));
  inv1  gate873(.a(s_47), .O(gate463inter4));
  nand2 gate874(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate875(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate876(.a(G23), .O(gate463inter7));
  inv1  gate877(.a(G1198), .O(gate463inter8));
  nand2 gate878(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate879(.a(s_47), .b(gate463inter3), .O(gate463inter10));
  nor2  gate880(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate881(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate882(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1513(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1514(.a(gate464inter0), .b(s_138), .O(gate464inter1));
  and2  gate1515(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1516(.a(s_138), .O(gate464inter3));
  inv1  gate1517(.a(s_139), .O(gate464inter4));
  nand2 gate1518(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1519(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1520(.a(G1102), .O(gate464inter7));
  inv1  gate1521(.a(G1198), .O(gate464inter8));
  nand2 gate1522(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1523(.a(s_139), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1524(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1525(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1526(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1527(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1528(.a(gate471inter0), .b(s_140), .O(gate471inter1));
  and2  gate1529(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1530(.a(s_140), .O(gate471inter3));
  inv1  gate1531(.a(s_141), .O(gate471inter4));
  nand2 gate1532(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1533(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1534(.a(G27), .O(gate471inter7));
  inv1  gate1535(.a(G1210), .O(gate471inter8));
  nand2 gate1536(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1537(.a(s_141), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1538(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1539(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1540(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1009(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1010(.a(gate472inter0), .b(s_66), .O(gate472inter1));
  and2  gate1011(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1012(.a(s_66), .O(gate472inter3));
  inv1  gate1013(.a(s_67), .O(gate472inter4));
  nand2 gate1014(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1015(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1016(.a(G1114), .O(gate472inter7));
  inv1  gate1017(.a(G1210), .O(gate472inter8));
  nand2 gate1018(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1019(.a(s_67), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1020(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1021(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1022(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate995(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate996(.a(gate483inter0), .b(s_64), .O(gate483inter1));
  and2  gate997(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate998(.a(s_64), .O(gate483inter3));
  inv1  gate999(.a(s_65), .O(gate483inter4));
  nand2 gate1000(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1001(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1002(.a(G1228), .O(gate483inter7));
  inv1  gate1003(.a(G1229), .O(gate483inter8));
  nand2 gate1004(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1005(.a(s_65), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1006(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1007(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1008(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1723(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1724(.a(gate486inter0), .b(s_168), .O(gate486inter1));
  and2  gate1725(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1726(.a(s_168), .O(gate486inter3));
  inv1  gate1727(.a(s_169), .O(gate486inter4));
  nand2 gate1728(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1729(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1730(.a(G1234), .O(gate486inter7));
  inv1  gate1731(.a(G1235), .O(gate486inter8));
  nand2 gate1732(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1733(.a(s_169), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1734(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1735(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1736(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1471(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1472(.a(gate488inter0), .b(s_132), .O(gate488inter1));
  and2  gate1473(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1474(.a(s_132), .O(gate488inter3));
  inv1  gate1475(.a(s_133), .O(gate488inter4));
  nand2 gate1476(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1477(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1478(.a(G1238), .O(gate488inter7));
  inv1  gate1479(.a(G1239), .O(gate488inter8));
  nand2 gate1480(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1481(.a(s_133), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1482(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1483(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1484(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1401(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1402(.a(gate490inter0), .b(s_122), .O(gate490inter1));
  and2  gate1403(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1404(.a(s_122), .O(gate490inter3));
  inv1  gate1405(.a(s_123), .O(gate490inter4));
  nand2 gate1406(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1407(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1408(.a(G1242), .O(gate490inter7));
  inv1  gate1409(.a(G1243), .O(gate490inter8));
  nand2 gate1410(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1411(.a(s_123), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1412(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1413(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1414(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1863(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1864(.a(gate491inter0), .b(s_188), .O(gate491inter1));
  and2  gate1865(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1866(.a(s_188), .O(gate491inter3));
  inv1  gate1867(.a(s_189), .O(gate491inter4));
  nand2 gate1868(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1869(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1870(.a(G1244), .O(gate491inter7));
  inv1  gate1871(.a(G1245), .O(gate491inter8));
  nand2 gate1872(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1873(.a(s_189), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1874(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1875(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1876(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate855(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate856(.a(gate494inter0), .b(s_44), .O(gate494inter1));
  and2  gate857(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate858(.a(s_44), .O(gate494inter3));
  inv1  gate859(.a(s_45), .O(gate494inter4));
  nand2 gate860(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate861(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate862(.a(G1250), .O(gate494inter7));
  inv1  gate863(.a(G1251), .O(gate494inter8));
  nand2 gate864(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate865(.a(s_45), .b(gate494inter3), .O(gate494inter10));
  nor2  gate866(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate867(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate868(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2297(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2298(.a(gate497inter0), .b(s_250), .O(gate497inter1));
  and2  gate2299(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2300(.a(s_250), .O(gate497inter3));
  inv1  gate2301(.a(s_251), .O(gate497inter4));
  nand2 gate2302(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2303(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2304(.a(G1256), .O(gate497inter7));
  inv1  gate2305(.a(G1257), .O(gate497inter8));
  nand2 gate2306(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2307(.a(s_251), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2308(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2309(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2310(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1121(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1122(.a(gate501inter0), .b(s_82), .O(gate501inter1));
  and2  gate1123(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1124(.a(s_82), .O(gate501inter3));
  inv1  gate1125(.a(s_83), .O(gate501inter4));
  nand2 gate1126(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1127(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1128(.a(G1264), .O(gate501inter7));
  inv1  gate1129(.a(G1265), .O(gate501inter8));
  nand2 gate1130(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1131(.a(s_83), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1132(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1133(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1134(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2227(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2228(.a(gate503inter0), .b(s_240), .O(gate503inter1));
  and2  gate2229(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2230(.a(s_240), .O(gate503inter3));
  inv1  gate2231(.a(s_241), .O(gate503inter4));
  nand2 gate2232(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2233(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2234(.a(G1268), .O(gate503inter7));
  inv1  gate2235(.a(G1269), .O(gate503inter8));
  nand2 gate2236(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2237(.a(s_241), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2238(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2239(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2240(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1611(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1612(.a(gate506inter0), .b(s_152), .O(gate506inter1));
  and2  gate1613(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1614(.a(s_152), .O(gate506inter3));
  inv1  gate1615(.a(s_153), .O(gate506inter4));
  nand2 gate1616(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1617(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1618(.a(G1274), .O(gate506inter7));
  inv1  gate1619(.a(G1275), .O(gate506inter8));
  nand2 gate1620(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1621(.a(s_153), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1622(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1623(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1624(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule