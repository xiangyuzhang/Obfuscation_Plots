module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate645(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate646(.a(gate14inter0), .b(s_14), .O(gate14inter1));
  and2  gate647(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate648(.a(s_14), .O(gate14inter3));
  inv1  gate649(.a(s_15), .O(gate14inter4));
  nand2 gate650(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate651(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate652(.a(G11), .O(gate14inter7));
  inv1  gate653(.a(G12), .O(gate14inter8));
  nand2 gate654(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate655(.a(s_15), .b(gate14inter3), .O(gate14inter10));
  nor2  gate656(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate657(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate658(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1093(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1094(.a(gate19inter0), .b(s_78), .O(gate19inter1));
  and2  gate1095(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1096(.a(s_78), .O(gate19inter3));
  inv1  gate1097(.a(s_79), .O(gate19inter4));
  nand2 gate1098(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1099(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1100(.a(G21), .O(gate19inter7));
  inv1  gate1101(.a(G22), .O(gate19inter8));
  nand2 gate1102(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1103(.a(s_79), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1104(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1105(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1106(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate925(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate926(.a(gate48inter0), .b(s_54), .O(gate48inter1));
  and2  gate927(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate928(.a(s_54), .O(gate48inter3));
  inv1  gate929(.a(s_55), .O(gate48inter4));
  nand2 gate930(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate931(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate932(.a(G8), .O(gate48inter7));
  inv1  gate933(.a(G275), .O(gate48inter8));
  nand2 gate934(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate935(.a(s_55), .b(gate48inter3), .O(gate48inter10));
  nor2  gate936(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate937(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate938(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate911(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate912(.a(gate49inter0), .b(s_52), .O(gate49inter1));
  and2  gate913(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate914(.a(s_52), .O(gate49inter3));
  inv1  gate915(.a(s_53), .O(gate49inter4));
  nand2 gate916(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate917(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate918(.a(G9), .O(gate49inter7));
  inv1  gate919(.a(G278), .O(gate49inter8));
  nand2 gate920(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate921(.a(s_53), .b(gate49inter3), .O(gate49inter10));
  nor2  gate922(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate923(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate924(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1191(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1192(.a(gate53inter0), .b(s_92), .O(gate53inter1));
  and2  gate1193(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1194(.a(s_92), .O(gate53inter3));
  inv1  gate1195(.a(s_93), .O(gate53inter4));
  nand2 gate1196(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1197(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1198(.a(G13), .O(gate53inter7));
  inv1  gate1199(.a(G284), .O(gate53inter8));
  nand2 gate1200(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1201(.a(s_93), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1202(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1203(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1204(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate883(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate884(.a(gate60inter0), .b(s_48), .O(gate60inter1));
  and2  gate885(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate886(.a(s_48), .O(gate60inter3));
  inv1  gate887(.a(s_49), .O(gate60inter4));
  nand2 gate888(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate889(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate890(.a(G20), .O(gate60inter7));
  inv1  gate891(.a(G293), .O(gate60inter8));
  nand2 gate892(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate893(.a(s_49), .b(gate60inter3), .O(gate60inter10));
  nor2  gate894(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate895(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate896(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate897(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate898(.a(gate61inter0), .b(s_50), .O(gate61inter1));
  and2  gate899(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate900(.a(s_50), .O(gate61inter3));
  inv1  gate901(.a(s_51), .O(gate61inter4));
  nand2 gate902(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate903(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate904(.a(G21), .O(gate61inter7));
  inv1  gate905(.a(G296), .O(gate61inter8));
  nand2 gate906(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate907(.a(s_51), .b(gate61inter3), .O(gate61inter10));
  nor2  gate908(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate909(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate910(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1009(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1010(.a(gate66inter0), .b(s_66), .O(gate66inter1));
  and2  gate1011(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1012(.a(s_66), .O(gate66inter3));
  inv1  gate1013(.a(s_67), .O(gate66inter4));
  nand2 gate1014(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1015(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1016(.a(G26), .O(gate66inter7));
  inv1  gate1017(.a(G302), .O(gate66inter8));
  nand2 gate1018(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1019(.a(s_67), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1020(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1021(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1022(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate939(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate940(.a(gate67inter0), .b(s_56), .O(gate67inter1));
  and2  gate941(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate942(.a(s_56), .O(gate67inter3));
  inv1  gate943(.a(s_57), .O(gate67inter4));
  nand2 gate944(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate945(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate946(.a(G27), .O(gate67inter7));
  inv1  gate947(.a(G305), .O(gate67inter8));
  nand2 gate948(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate949(.a(s_57), .b(gate67inter3), .O(gate67inter10));
  nor2  gate950(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate951(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate952(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate617(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate618(.a(gate71inter0), .b(s_10), .O(gate71inter1));
  and2  gate619(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate620(.a(s_10), .O(gate71inter3));
  inv1  gate621(.a(s_11), .O(gate71inter4));
  nand2 gate622(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate623(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate624(.a(G31), .O(gate71inter7));
  inv1  gate625(.a(G311), .O(gate71inter8));
  nand2 gate626(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate627(.a(s_11), .b(gate71inter3), .O(gate71inter10));
  nor2  gate628(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate629(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate630(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1177(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1178(.a(gate72inter0), .b(s_90), .O(gate72inter1));
  and2  gate1179(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1180(.a(s_90), .O(gate72inter3));
  inv1  gate1181(.a(s_91), .O(gate72inter4));
  nand2 gate1182(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1183(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1184(.a(G32), .O(gate72inter7));
  inv1  gate1185(.a(G311), .O(gate72inter8));
  nand2 gate1186(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1187(.a(s_91), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1188(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1189(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1190(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate967(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate968(.a(gate77inter0), .b(s_60), .O(gate77inter1));
  and2  gate969(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate970(.a(s_60), .O(gate77inter3));
  inv1  gate971(.a(s_61), .O(gate77inter4));
  nand2 gate972(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate973(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate974(.a(G2), .O(gate77inter7));
  inv1  gate975(.a(G320), .O(gate77inter8));
  nand2 gate976(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate977(.a(s_61), .b(gate77inter3), .O(gate77inter10));
  nor2  gate978(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate979(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate980(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1219(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1220(.a(gate78inter0), .b(s_96), .O(gate78inter1));
  and2  gate1221(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1222(.a(s_96), .O(gate78inter3));
  inv1  gate1223(.a(s_97), .O(gate78inter4));
  nand2 gate1224(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1225(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1226(.a(G6), .O(gate78inter7));
  inv1  gate1227(.a(G320), .O(gate78inter8));
  nand2 gate1228(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1229(.a(s_97), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1230(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1231(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1232(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate659(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate660(.a(gate81inter0), .b(s_16), .O(gate81inter1));
  and2  gate661(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate662(.a(s_16), .O(gate81inter3));
  inv1  gate663(.a(s_17), .O(gate81inter4));
  nand2 gate664(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate665(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate666(.a(G3), .O(gate81inter7));
  inv1  gate667(.a(G326), .O(gate81inter8));
  nand2 gate668(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate669(.a(s_17), .b(gate81inter3), .O(gate81inter10));
  nor2  gate670(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate671(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate672(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1261(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1262(.a(gate83inter0), .b(s_102), .O(gate83inter1));
  and2  gate1263(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1264(.a(s_102), .O(gate83inter3));
  inv1  gate1265(.a(s_103), .O(gate83inter4));
  nand2 gate1266(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1267(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1268(.a(G11), .O(gate83inter7));
  inv1  gate1269(.a(G329), .O(gate83inter8));
  nand2 gate1270(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1271(.a(s_103), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1272(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1273(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1274(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1163(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1164(.a(gate93inter0), .b(s_88), .O(gate93inter1));
  and2  gate1165(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1166(.a(s_88), .O(gate93inter3));
  inv1  gate1167(.a(s_89), .O(gate93inter4));
  nand2 gate1168(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1169(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1170(.a(G18), .O(gate93inter7));
  inv1  gate1171(.a(G344), .O(gate93inter8));
  nand2 gate1172(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1173(.a(s_89), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1174(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1175(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1176(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate575(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate576(.a(gate95inter0), .b(s_4), .O(gate95inter1));
  and2  gate577(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate578(.a(s_4), .O(gate95inter3));
  inv1  gate579(.a(s_5), .O(gate95inter4));
  nand2 gate580(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate581(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate582(.a(G26), .O(gate95inter7));
  inv1  gate583(.a(G347), .O(gate95inter8));
  nand2 gate584(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate585(.a(s_5), .b(gate95inter3), .O(gate95inter10));
  nor2  gate586(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate587(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate588(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate841(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate842(.a(gate118inter0), .b(s_42), .O(gate118inter1));
  and2  gate843(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate844(.a(s_42), .O(gate118inter3));
  inv1  gate845(.a(s_43), .O(gate118inter4));
  nand2 gate846(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate847(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate848(.a(G388), .O(gate118inter7));
  inv1  gate849(.a(G389), .O(gate118inter8));
  nand2 gate850(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate851(.a(s_43), .b(gate118inter3), .O(gate118inter10));
  nor2  gate852(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate853(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate854(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate715(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate716(.a(gate126inter0), .b(s_24), .O(gate126inter1));
  and2  gate717(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate718(.a(s_24), .O(gate126inter3));
  inv1  gate719(.a(s_25), .O(gate126inter4));
  nand2 gate720(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate721(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate722(.a(G404), .O(gate126inter7));
  inv1  gate723(.a(G405), .O(gate126inter8));
  nand2 gate724(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate725(.a(s_25), .b(gate126inter3), .O(gate126inter10));
  nor2  gate726(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate727(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate728(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate953(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate954(.a(gate127inter0), .b(s_58), .O(gate127inter1));
  and2  gate955(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate956(.a(s_58), .O(gate127inter3));
  inv1  gate957(.a(s_59), .O(gate127inter4));
  nand2 gate958(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate959(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate960(.a(G406), .O(gate127inter7));
  inv1  gate961(.a(G407), .O(gate127inter8));
  nand2 gate962(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate963(.a(s_59), .b(gate127inter3), .O(gate127inter10));
  nor2  gate964(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate965(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate966(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate785(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate786(.a(gate132inter0), .b(s_34), .O(gate132inter1));
  and2  gate787(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate788(.a(s_34), .O(gate132inter3));
  inv1  gate789(.a(s_35), .O(gate132inter4));
  nand2 gate790(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate791(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate792(.a(G416), .O(gate132inter7));
  inv1  gate793(.a(G417), .O(gate132inter8));
  nand2 gate794(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate795(.a(s_35), .b(gate132inter3), .O(gate132inter10));
  nor2  gate796(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate797(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate798(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate995(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate996(.a(gate149inter0), .b(s_64), .O(gate149inter1));
  and2  gate997(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate998(.a(s_64), .O(gate149inter3));
  inv1  gate999(.a(s_65), .O(gate149inter4));
  nand2 gate1000(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1001(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1002(.a(G498), .O(gate149inter7));
  inv1  gate1003(.a(G501), .O(gate149inter8));
  nand2 gate1004(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1005(.a(s_65), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1006(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1007(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1008(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate589(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate590(.a(gate151inter0), .b(s_6), .O(gate151inter1));
  and2  gate591(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate592(.a(s_6), .O(gate151inter3));
  inv1  gate593(.a(s_7), .O(gate151inter4));
  nand2 gate594(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate595(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate596(.a(G510), .O(gate151inter7));
  inv1  gate597(.a(G513), .O(gate151inter8));
  nand2 gate598(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate599(.a(s_7), .b(gate151inter3), .O(gate151inter10));
  nor2  gate600(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate601(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate602(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1023(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1024(.a(gate171inter0), .b(s_68), .O(gate171inter1));
  and2  gate1025(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1026(.a(s_68), .O(gate171inter3));
  inv1  gate1027(.a(s_69), .O(gate171inter4));
  nand2 gate1028(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1029(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1030(.a(G480), .O(gate171inter7));
  inv1  gate1031(.a(G549), .O(gate171inter8));
  nand2 gate1032(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1033(.a(s_69), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1034(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1035(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1036(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate869(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate870(.a(gate178inter0), .b(s_46), .O(gate178inter1));
  and2  gate871(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate872(.a(s_46), .O(gate178inter3));
  inv1  gate873(.a(s_47), .O(gate178inter4));
  nand2 gate874(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate875(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate876(.a(G501), .O(gate178inter7));
  inv1  gate877(.a(G558), .O(gate178inter8));
  nand2 gate878(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate879(.a(s_47), .b(gate178inter3), .O(gate178inter10));
  nor2  gate880(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate881(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate882(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate701(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate702(.a(gate179inter0), .b(s_22), .O(gate179inter1));
  and2  gate703(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate704(.a(s_22), .O(gate179inter3));
  inv1  gate705(.a(s_23), .O(gate179inter4));
  nand2 gate706(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate707(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate708(.a(G504), .O(gate179inter7));
  inv1  gate709(.a(G561), .O(gate179inter8));
  nand2 gate710(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate711(.a(s_23), .b(gate179inter3), .O(gate179inter10));
  nor2  gate712(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate713(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate714(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate673(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate674(.a(gate186inter0), .b(s_18), .O(gate186inter1));
  and2  gate675(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate676(.a(s_18), .O(gate186inter3));
  inv1  gate677(.a(s_19), .O(gate186inter4));
  nand2 gate678(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate679(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate680(.a(G572), .O(gate186inter7));
  inv1  gate681(.a(G573), .O(gate186inter8));
  nand2 gate682(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate683(.a(s_19), .b(gate186inter3), .O(gate186inter10));
  nor2  gate684(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate685(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate686(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate981(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate982(.a(gate192inter0), .b(s_62), .O(gate192inter1));
  and2  gate983(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate984(.a(s_62), .O(gate192inter3));
  inv1  gate985(.a(s_63), .O(gate192inter4));
  nand2 gate986(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate987(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate988(.a(G584), .O(gate192inter7));
  inv1  gate989(.a(G585), .O(gate192inter8));
  nand2 gate990(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate991(.a(s_63), .b(gate192inter3), .O(gate192inter10));
  nor2  gate992(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate993(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate994(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1233(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1234(.a(gate200inter0), .b(s_98), .O(gate200inter1));
  and2  gate1235(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1236(.a(s_98), .O(gate200inter3));
  inv1  gate1237(.a(s_99), .O(gate200inter4));
  nand2 gate1238(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1239(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1240(.a(G600), .O(gate200inter7));
  inv1  gate1241(.a(G601), .O(gate200inter8));
  nand2 gate1242(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1243(.a(s_99), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1244(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1245(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1246(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate561(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate562(.a(gate201inter0), .b(s_2), .O(gate201inter1));
  and2  gate563(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate564(.a(s_2), .O(gate201inter3));
  inv1  gate565(.a(s_3), .O(gate201inter4));
  nand2 gate566(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate567(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate568(.a(G602), .O(gate201inter7));
  inv1  gate569(.a(G607), .O(gate201inter8));
  nand2 gate570(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate571(.a(s_3), .b(gate201inter3), .O(gate201inter10));
  nor2  gate572(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate573(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate574(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate799(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate800(.a(gate205inter0), .b(s_36), .O(gate205inter1));
  and2  gate801(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate802(.a(s_36), .O(gate205inter3));
  inv1  gate803(.a(s_37), .O(gate205inter4));
  nand2 gate804(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate805(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate806(.a(G622), .O(gate205inter7));
  inv1  gate807(.a(G627), .O(gate205inter8));
  nand2 gate808(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate809(.a(s_37), .b(gate205inter3), .O(gate205inter10));
  nor2  gate810(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate811(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate812(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate687(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate688(.a(gate206inter0), .b(s_20), .O(gate206inter1));
  and2  gate689(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate690(.a(s_20), .O(gate206inter3));
  inv1  gate691(.a(s_21), .O(gate206inter4));
  nand2 gate692(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate693(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate694(.a(G632), .O(gate206inter7));
  inv1  gate695(.a(G637), .O(gate206inter8));
  nand2 gate696(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate697(.a(s_21), .b(gate206inter3), .O(gate206inter10));
  nor2  gate698(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate699(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate700(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1247(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1248(.a(gate234inter0), .b(s_100), .O(gate234inter1));
  and2  gate1249(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1250(.a(s_100), .O(gate234inter3));
  inv1  gate1251(.a(s_101), .O(gate234inter4));
  nand2 gate1252(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1253(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1254(.a(G245), .O(gate234inter7));
  inv1  gate1255(.a(G721), .O(gate234inter8));
  nand2 gate1256(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1257(.a(s_101), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1258(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1259(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1260(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1317(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1318(.a(gate240inter0), .b(s_110), .O(gate240inter1));
  and2  gate1319(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1320(.a(s_110), .O(gate240inter3));
  inv1  gate1321(.a(s_111), .O(gate240inter4));
  nand2 gate1322(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1323(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1324(.a(G263), .O(gate240inter7));
  inv1  gate1325(.a(G715), .O(gate240inter8));
  nand2 gate1326(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1327(.a(s_111), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1328(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1329(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1330(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1065(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1066(.a(gate243inter0), .b(s_74), .O(gate243inter1));
  and2  gate1067(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1068(.a(s_74), .O(gate243inter3));
  inv1  gate1069(.a(s_75), .O(gate243inter4));
  nand2 gate1070(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1071(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1072(.a(G245), .O(gate243inter7));
  inv1  gate1073(.a(G733), .O(gate243inter8));
  nand2 gate1074(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1075(.a(s_75), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1076(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1077(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1078(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate771(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate772(.a(gate249inter0), .b(s_32), .O(gate249inter1));
  and2  gate773(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate774(.a(s_32), .O(gate249inter3));
  inv1  gate775(.a(s_33), .O(gate249inter4));
  nand2 gate776(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate777(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate778(.a(G254), .O(gate249inter7));
  inv1  gate779(.a(G742), .O(gate249inter8));
  nand2 gate780(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate781(.a(s_33), .b(gate249inter3), .O(gate249inter10));
  nor2  gate782(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate783(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate784(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate743(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate744(.a(gate286inter0), .b(s_28), .O(gate286inter1));
  and2  gate745(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate746(.a(s_28), .O(gate286inter3));
  inv1  gate747(.a(s_29), .O(gate286inter4));
  nand2 gate748(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate749(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate750(.a(G788), .O(gate286inter7));
  inv1  gate751(.a(G812), .O(gate286inter8));
  nand2 gate752(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate753(.a(s_29), .b(gate286inter3), .O(gate286inter10));
  nor2  gate754(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate755(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate756(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1275(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1276(.a(gate390inter0), .b(s_104), .O(gate390inter1));
  and2  gate1277(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1278(.a(s_104), .O(gate390inter3));
  inv1  gate1279(.a(s_105), .O(gate390inter4));
  nand2 gate1280(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1281(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1282(.a(G4), .O(gate390inter7));
  inv1  gate1283(.a(G1045), .O(gate390inter8));
  nand2 gate1284(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1285(.a(s_105), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1286(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1287(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1288(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate547(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate548(.a(gate393inter0), .b(s_0), .O(gate393inter1));
  and2  gate549(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate550(.a(s_0), .O(gate393inter3));
  inv1  gate551(.a(s_1), .O(gate393inter4));
  nand2 gate552(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate553(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate554(.a(G7), .O(gate393inter7));
  inv1  gate555(.a(G1054), .O(gate393inter8));
  nand2 gate556(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate557(.a(s_1), .b(gate393inter3), .O(gate393inter10));
  nor2  gate558(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate559(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate560(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate855(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate856(.a(gate400inter0), .b(s_44), .O(gate400inter1));
  and2  gate857(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate858(.a(s_44), .O(gate400inter3));
  inv1  gate859(.a(s_45), .O(gate400inter4));
  nand2 gate860(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate861(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate862(.a(G14), .O(gate400inter7));
  inv1  gate863(.a(G1075), .O(gate400inter8));
  nand2 gate864(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate865(.a(s_45), .b(gate400inter3), .O(gate400inter10));
  nor2  gate866(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate867(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate868(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1205(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1206(.a(gate413inter0), .b(s_94), .O(gate413inter1));
  and2  gate1207(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1208(.a(s_94), .O(gate413inter3));
  inv1  gate1209(.a(s_95), .O(gate413inter4));
  nand2 gate1210(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1211(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1212(.a(G27), .O(gate413inter7));
  inv1  gate1213(.a(G1114), .O(gate413inter8));
  nand2 gate1214(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1215(.a(s_95), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1216(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1217(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1218(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate757(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate758(.a(gate421inter0), .b(s_30), .O(gate421inter1));
  and2  gate759(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate760(.a(s_30), .O(gate421inter3));
  inv1  gate761(.a(s_31), .O(gate421inter4));
  nand2 gate762(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate763(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate764(.a(G2), .O(gate421inter7));
  inv1  gate765(.a(G1135), .O(gate421inter8));
  nand2 gate766(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate767(.a(s_31), .b(gate421inter3), .O(gate421inter10));
  nor2  gate768(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate769(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate770(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1037(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1038(.a(gate426inter0), .b(s_70), .O(gate426inter1));
  and2  gate1039(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1040(.a(s_70), .O(gate426inter3));
  inv1  gate1041(.a(s_71), .O(gate426inter4));
  nand2 gate1042(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1043(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1044(.a(G1045), .O(gate426inter7));
  inv1  gate1045(.a(G1141), .O(gate426inter8));
  nand2 gate1046(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1047(.a(s_71), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1048(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1049(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1050(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1107(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1108(.a(gate427inter0), .b(s_80), .O(gate427inter1));
  and2  gate1109(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1110(.a(s_80), .O(gate427inter3));
  inv1  gate1111(.a(s_81), .O(gate427inter4));
  nand2 gate1112(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1113(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1114(.a(G5), .O(gate427inter7));
  inv1  gate1115(.a(G1144), .O(gate427inter8));
  nand2 gate1116(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1117(.a(s_81), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1118(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1119(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1120(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1121(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1122(.a(gate431inter0), .b(s_82), .O(gate431inter1));
  and2  gate1123(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1124(.a(s_82), .O(gate431inter3));
  inv1  gate1125(.a(s_83), .O(gate431inter4));
  nand2 gate1126(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1127(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1128(.a(G7), .O(gate431inter7));
  inv1  gate1129(.a(G1150), .O(gate431inter8));
  nand2 gate1130(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1131(.a(s_83), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1132(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1133(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1134(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate813(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate814(.a(gate434inter0), .b(s_38), .O(gate434inter1));
  and2  gate815(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate816(.a(s_38), .O(gate434inter3));
  inv1  gate817(.a(s_39), .O(gate434inter4));
  nand2 gate818(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate819(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate820(.a(G1057), .O(gate434inter7));
  inv1  gate821(.a(G1153), .O(gate434inter8));
  nand2 gate822(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate823(.a(s_39), .b(gate434inter3), .O(gate434inter10));
  nor2  gate824(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate825(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate826(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate729(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate730(.a(gate436inter0), .b(s_26), .O(gate436inter1));
  and2  gate731(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate732(.a(s_26), .O(gate436inter3));
  inv1  gate733(.a(s_27), .O(gate436inter4));
  nand2 gate734(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate735(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate736(.a(G1060), .O(gate436inter7));
  inv1  gate737(.a(G1156), .O(gate436inter8));
  nand2 gate738(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate739(.a(s_27), .b(gate436inter3), .O(gate436inter10));
  nor2  gate740(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate741(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate742(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate631(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate632(.a(gate440inter0), .b(s_12), .O(gate440inter1));
  and2  gate633(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate634(.a(s_12), .O(gate440inter3));
  inv1  gate635(.a(s_13), .O(gate440inter4));
  nand2 gate636(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate637(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate638(.a(G1066), .O(gate440inter7));
  inv1  gate639(.a(G1162), .O(gate440inter8));
  nand2 gate640(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate641(.a(s_13), .b(gate440inter3), .O(gate440inter10));
  nor2  gate642(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate643(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate644(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1149(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1150(.a(gate454inter0), .b(s_86), .O(gate454inter1));
  and2  gate1151(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1152(.a(s_86), .O(gate454inter3));
  inv1  gate1153(.a(s_87), .O(gate454inter4));
  nand2 gate1154(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1155(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1156(.a(G1087), .O(gate454inter7));
  inv1  gate1157(.a(G1183), .O(gate454inter8));
  nand2 gate1158(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1159(.a(s_87), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1160(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1161(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1162(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1079(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1080(.a(gate463inter0), .b(s_76), .O(gate463inter1));
  and2  gate1081(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1082(.a(s_76), .O(gate463inter3));
  inv1  gate1083(.a(s_77), .O(gate463inter4));
  nand2 gate1084(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1085(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1086(.a(G23), .O(gate463inter7));
  inv1  gate1087(.a(G1198), .O(gate463inter8));
  nand2 gate1088(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1089(.a(s_77), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1090(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1091(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1092(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1135(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1136(.a(gate467inter0), .b(s_84), .O(gate467inter1));
  and2  gate1137(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1138(.a(s_84), .O(gate467inter3));
  inv1  gate1139(.a(s_85), .O(gate467inter4));
  nand2 gate1140(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1141(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1142(.a(G25), .O(gate467inter7));
  inv1  gate1143(.a(G1204), .O(gate467inter8));
  nand2 gate1144(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1145(.a(s_85), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1146(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1147(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1148(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1289(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1290(.a(gate480inter0), .b(s_106), .O(gate480inter1));
  and2  gate1291(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1292(.a(s_106), .O(gate480inter3));
  inv1  gate1293(.a(s_107), .O(gate480inter4));
  nand2 gate1294(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1295(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1296(.a(G1126), .O(gate480inter7));
  inv1  gate1297(.a(G1222), .O(gate480inter8));
  nand2 gate1298(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1299(.a(s_107), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1300(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1301(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1302(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate827(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate828(.a(gate483inter0), .b(s_40), .O(gate483inter1));
  and2  gate829(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate830(.a(s_40), .O(gate483inter3));
  inv1  gate831(.a(s_41), .O(gate483inter4));
  nand2 gate832(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate833(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate834(.a(G1228), .O(gate483inter7));
  inv1  gate835(.a(G1229), .O(gate483inter8));
  nand2 gate836(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate837(.a(s_41), .b(gate483inter3), .O(gate483inter10));
  nor2  gate838(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate839(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate840(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1303(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1304(.a(gate491inter0), .b(s_108), .O(gate491inter1));
  and2  gate1305(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1306(.a(s_108), .O(gate491inter3));
  inv1  gate1307(.a(s_109), .O(gate491inter4));
  nand2 gate1308(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1309(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1310(.a(G1244), .O(gate491inter7));
  inv1  gate1311(.a(G1245), .O(gate491inter8));
  nand2 gate1312(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1313(.a(s_109), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1314(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1315(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1316(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate603(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate604(.a(gate501inter0), .b(s_8), .O(gate501inter1));
  and2  gate605(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate606(.a(s_8), .O(gate501inter3));
  inv1  gate607(.a(s_9), .O(gate501inter4));
  nand2 gate608(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate609(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate610(.a(G1264), .O(gate501inter7));
  inv1  gate611(.a(G1265), .O(gate501inter8));
  nand2 gate612(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate613(.a(s_9), .b(gate501inter3), .O(gate501inter10));
  nor2  gate614(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate615(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate616(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1051(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1052(.a(gate505inter0), .b(s_72), .O(gate505inter1));
  and2  gate1053(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1054(.a(s_72), .O(gate505inter3));
  inv1  gate1055(.a(s_73), .O(gate505inter4));
  nand2 gate1056(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1057(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1058(.a(G1272), .O(gate505inter7));
  inv1  gate1059(.a(G1273), .O(gate505inter8));
  nand2 gate1060(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1061(.a(s_73), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1062(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1063(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1064(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule