module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate813(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate814(.a(gate9inter0), .b(s_38), .O(gate9inter1));
  and2  gate815(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate816(.a(s_38), .O(gate9inter3));
  inv1  gate817(.a(s_39), .O(gate9inter4));
  nand2 gate818(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate819(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate820(.a(G1), .O(gate9inter7));
  inv1  gate821(.a(G2), .O(gate9inter8));
  nand2 gate822(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate823(.a(s_39), .b(gate9inter3), .O(gate9inter10));
  nor2  gate824(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate825(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate826(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1303(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1304(.a(gate12inter0), .b(s_108), .O(gate12inter1));
  and2  gate1305(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1306(.a(s_108), .O(gate12inter3));
  inv1  gate1307(.a(s_109), .O(gate12inter4));
  nand2 gate1308(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1309(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1310(.a(G7), .O(gate12inter7));
  inv1  gate1311(.a(G8), .O(gate12inter8));
  nand2 gate1312(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1313(.a(s_109), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1314(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1315(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1316(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate659(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate660(.a(gate14inter0), .b(s_16), .O(gate14inter1));
  and2  gate661(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate662(.a(s_16), .O(gate14inter3));
  inv1  gate663(.a(s_17), .O(gate14inter4));
  nand2 gate664(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate665(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate666(.a(G11), .O(gate14inter7));
  inv1  gate667(.a(G12), .O(gate14inter8));
  nand2 gate668(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate669(.a(s_17), .b(gate14inter3), .O(gate14inter10));
  nor2  gate670(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate671(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate672(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1471(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1472(.a(gate16inter0), .b(s_132), .O(gate16inter1));
  and2  gate1473(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1474(.a(s_132), .O(gate16inter3));
  inv1  gate1475(.a(s_133), .O(gate16inter4));
  nand2 gate1476(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1477(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1478(.a(G15), .O(gate16inter7));
  inv1  gate1479(.a(G16), .O(gate16inter8));
  nand2 gate1480(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1481(.a(s_133), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1482(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1483(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1484(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2157(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2158(.a(gate20inter0), .b(s_230), .O(gate20inter1));
  and2  gate2159(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2160(.a(s_230), .O(gate20inter3));
  inv1  gate2161(.a(s_231), .O(gate20inter4));
  nand2 gate2162(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2163(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2164(.a(G23), .O(gate20inter7));
  inv1  gate2165(.a(G24), .O(gate20inter8));
  nand2 gate2166(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2167(.a(s_231), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2168(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2169(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2170(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2353(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2354(.a(gate22inter0), .b(s_258), .O(gate22inter1));
  and2  gate2355(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2356(.a(s_258), .O(gate22inter3));
  inv1  gate2357(.a(s_259), .O(gate22inter4));
  nand2 gate2358(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2359(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2360(.a(G27), .O(gate22inter7));
  inv1  gate2361(.a(G28), .O(gate22inter8));
  nand2 gate2362(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2363(.a(s_259), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2364(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2365(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2366(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate729(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate730(.a(gate23inter0), .b(s_26), .O(gate23inter1));
  and2  gate731(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate732(.a(s_26), .O(gate23inter3));
  inv1  gate733(.a(s_27), .O(gate23inter4));
  nand2 gate734(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate735(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate736(.a(G29), .O(gate23inter7));
  inv1  gate737(.a(G30), .O(gate23inter8));
  nand2 gate738(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate739(.a(s_27), .b(gate23inter3), .O(gate23inter10));
  nor2  gate740(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate741(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate742(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1289(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1290(.a(gate26inter0), .b(s_106), .O(gate26inter1));
  and2  gate1291(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1292(.a(s_106), .O(gate26inter3));
  inv1  gate1293(.a(s_107), .O(gate26inter4));
  nand2 gate1294(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1295(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1296(.a(G9), .O(gate26inter7));
  inv1  gate1297(.a(G13), .O(gate26inter8));
  nand2 gate1298(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1299(.a(s_107), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1300(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1301(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1302(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1345(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1346(.a(gate29inter0), .b(s_114), .O(gate29inter1));
  and2  gate1347(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1348(.a(s_114), .O(gate29inter3));
  inv1  gate1349(.a(s_115), .O(gate29inter4));
  nand2 gate1350(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1351(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1352(.a(G3), .O(gate29inter7));
  inv1  gate1353(.a(G7), .O(gate29inter8));
  nand2 gate1354(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1355(.a(s_115), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1356(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1357(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1358(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate2689(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate2690(.a(gate38inter0), .b(s_306), .O(gate38inter1));
  and2  gate2691(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate2692(.a(s_306), .O(gate38inter3));
  inv1  gate2693(.a(s_307), .O(gate38inter4));
  nand2 gate2694(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate2695(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate2696(.a(G27), .O(gate38inter7));
  inv1  gate2697(.a(G31), .O(gate38inter8));
  nand2 gate2698(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate2699(.a(s_307), .b(gate38inter3), .O(gate38inter10));
  nor2  gate2700(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate2701(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate2702(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2563(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2564(.a(gate43inter0), .b(s_288), .O(gate43inter1));
  and2  gate2565(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2566(.a(s_288), .O(gate43inter3));
  inv1  gate2567(.a(s_289), .O(gate43inter4));
  nand2 gate2568(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2569(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2570(.a(G3), .O(gate43inter7));
  inv1  gate2571(.a(G269), .O(gate43inter8));
  nand2 gate2572(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2573(.a(s_289), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2574(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2575(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2576(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate2591(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2592(.a(gate48inter0), .b(s_292), .O(gate48inter1));
  and2  gate2593(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2594(.a(s_292), .O(gate48inter3));
  inv1  gate2595(.a(s_293), .O(gate48inter4));
  nand2 gate2596(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2597(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2598(.a(G8), .O(gate48inter7));
  inv1  gate2599(.a(G275), .O(gate48inter8));
  nand2 gate2600(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2601(.a(s_293), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2602(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2603(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2604(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1751(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1752(.a(gate49inter0), .b(s_172), .O(gate49inter1));
  and2  gate1753(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1754(.a(s_172), .O(gate49inter3));
  inv1  gate1755(.a(s_173), .O(gate49inter4));
  nand2 gate1756(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1757(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1758(.a(G9), .O(gate49inter7));
  inv1  gate1759(.a(G278), .O(gate49inter8));
  nand2 gate1760(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1761(.a(s_173), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1762(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1763(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1764(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2493(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2494(.a(gate50inter0), .b(s_278), .O(gate50inter1));
  and2  gate2495(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2496(.a(s_278), .O(gate50inter3));
  inv1  gate2497(.a(s_279), .O(gate50inter4));
  nand2 gate2498(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2499(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2500(.a(G10), .O(gate50inter7));
  inv1  gate2501(.a(G278), .O(gate50inter8));
  nand2 gate2502(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2503(.a(s_279), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2504(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2505(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2506(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1709(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1710(.a(gate53inter0), .b(s_166), .O(gate53inter1));
  and2  gate1711(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1712(.a(s_166), .O(gate53inter3));
  inv1  gate1713(.a(s_167), .O(gate53inter4));
  nand2 gate1714(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1715(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1716(.a(G13), .O(gate53inter7));
  inv1  gate1717(.a(G284), .O(gate53inter8));
  nand2 gate1718(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1719(.a(s_167), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1720(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1721(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1722(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1401(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1402(.a(gate57inter0), .b(s_122), .O(gate57inter1));
  and2  gate1403(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1404(.a(s_122), .O(gate57inter3));
  inv1  gate1405(.a(s_123), .O(gate57inter4));
  nand2 gate1406(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1407(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1408(.a(G17), .O(gate57inter7));
  inv1  gate1409(.a(G290), .O(gate57inter8));
  nand2 gate1410(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1411(.a(s_123), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1412(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1413(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1414(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1233(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1234(.a(gate61inter0), .b(s_98), .O(gate61inter1));
  and2  gate1235(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1236(.a(s_98), .O(gate61inter3));
  inv1  gate1237(.a(s_99), .O(gate61inter4));
  nand2 gate1238(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1239(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1240(.a(G21), .O(gate61inter7));
  inv1  gate1241(.a(G296), .O(gate61inter8));
  nand2 gate1242(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1243(.a(s_99), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1244(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1245(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1246(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2717(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2718(.a(gate66inter0), .b(s_310), .O(gate66inter1));
  and2  gate2719(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2720(.a(s_310), .O(gate66inter3));
  inv1  gate2721(.a(s_311), .O(gate66inter4));
  nand2 gate2722(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2723(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2724(.a(G26), .O(gate66inter7));
  inv1  gate2725(.a(G302), .O(gate66inter8));
  nand2 gate2726(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2727(.a(s_311), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2728(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2729(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2730(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2675(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2676(.a(gate70inter0), .b(s_304), .O(gate70inter1));
  and2  gate2677(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2678(.a(s_304), .O(gate70inter3));
  inv1  gate2679(.a(s_305), .O(gate70inter4));
  nand2 gate2680(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2681(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2682(.a(G30), .O(gate70inter7));
  inv1  gate2683(.a(G308), .O(gate70inter8));
  nand2 gate2684(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2685(.a(s_305), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2686(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2687(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2688(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1261(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1262(.a(gate71inter0), .b(s_102), .O(gate71inter1));
  and2  gate1263(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1264(.a(s_102), .O(gate71inter3));
  inv1  gate1265(.a(s_103), .O(gate71inter4));
  nand2 gate1266(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1267(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1268(.a(G31), .O(gate71inter7));
  inv1  gate1269(.a(G311), .O(gate71inter8));
  nand2 gate1270(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1271(.a(s_103), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1272(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1273(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1274(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2801(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2802(.a(gate72inter0), .b(s_322), .O(gate72inter1));
  and2  gate2803(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2804(.a(s_322), .O(gate72inter3));
  inv1  gate2805(.a(s_323), .O(gate72inter4));
  nand2 gate2806(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2807(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2808(.a(G32), .O(gate72inter7));
  inv1  gate2809(.a(G311), .O(gate72inter8));
  nand2 gate2810(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2811(.a(s_323), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2812(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2813(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2814(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate547(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate548(.a(gate77inter0), .b(s_0), .O(gate77inter1));
  and2  gate549(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate550(.a(s_0), .O(gate77inter3));
  inv1  gate551(.a(s_1), .O(gate77inter4));
  nand2 gate552(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate553(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate554(.a(G2), .O(gate77inter7));
  inv1  gate555(.a(G320), .O(gate77inter8));
  nand2 gate556(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate557(.a(s_1), .b(gate77inter3), .O(gate77inter10));
  nor2  gate558(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate559(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate560(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2283(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2284(.a(gate79inter0), .b(s_248), .O(gate79inter1));
  and2  gate2285(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2286(.a(s_248), .O(gate79inter3));
  inv1  gate2287(.a(s_249), .O(gate79inter4));
  nand2 gate2288(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2289(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2290(.a(G10), .O(gate79inter7));
  inv1  gate2291(.a(G323), .O(gate79inter8));
  nand2 gate2292(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2293(.a(s_249), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2294(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2295(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2296(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1037(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1038(.a(gate81inter0), .b(s_70), .O(gate81inter1));
  and2  gate1039(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1040(.a(s_70), .O(gate81inter3));
  inv1  gate1041(.a(s_71), .O(gate81inter4));
  nand2 gate1042(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1043(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1044(.a(G3), .O(gate81inter7));
  inv1  gate1045(.a(G326), .O(gate81inter8));
  nand2 gate1046(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1047(.a(s_71), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1048(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1049(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1050(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1499(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1500(.a(gate82inter0), .b(s_136), .O(gate82inter1));
  and2  gate1501(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1502(.a(s_136), .O(gate82inter3));
  inv1  gate1503(.a(s_137), .O(gate82inter4));
  nand2 gate1504(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1505(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1506(.a(G7), .O(gate82inter7));
  inv1  gate1507(.a(G326), .O(gate82inter8));
  nand2 gate1508(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1509(.a(s_137), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1510(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1511(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1512(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2367(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2368(.a(gate84inter0), .b(s_260), .O(gate84inter1));
  and2  gate2369(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2370(.a(s_260), .O(gate84inter3));
  inv1  gate2371(.a(s_261), .O(gate84inter4));
  nand2 gate2372(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2373(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2374(.a(G15), .O(gate84inter7));
  inv1  gate2375(.a(G329), .O(gate84inter8));
  nand2 gate2376(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2377(.a(s_261), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2378(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2379(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2380(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1177(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1178(.a(gate88inter0), .b(s_90), .O(gate88inter1));
  and2  gate1179(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1180(.a(s_90), .O(gate88inter3));
  inv1  gate1181(.a(s_91), .O(gate88inter4));
  nand2 gate1182(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1183(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1184(.a(G16), .O(gate88inter7));
  inv1  gate1185(.a(G335), .O(gate88inter8));
  nand2 gate1186(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1187(.a(s_91), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1188(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1189(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1190(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate925(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate926(.a(gate91inter0), .b(s_54), .O(gate91inter1));
  and2  gate927(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate928(.a(s_54), .O(gate91inter3));
  inv1  gate929(.a(s_55), .O(gate91inter4));
  nand2 gate930(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate931(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate932(.a(G25), .O(gate91inter7));
  inv1  gate933(.a(G341), .O(gate91inter8));
  nand2 gate934(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate935(.a(s_55), .b(gate91inter3), .O(gate91inter10));
  nor2  gate936(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate937(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate938(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate757(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate758(.a(gate93inter0), .b(s_30), .O(gate93inter1));
  and2  gate759(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate760(.a(s_30), .O(gate93inter3));
  inv1  gate761(.a(s_31), .O(gate93inter4));
  nand2 gate762(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate763(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate764(.a(G18), .O(gate93inter7));
  inv1  gate765(.a(G344), .O(gate93inter8));
  nand2 gate766(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate767(.a(s_31), .b(gate93inter3), .O(gate93inter10));
  nor2  gate768(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate769(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate770(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1989(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1990(.a(gate94inter0), .b(s_206), .O(gate94inter1));
  and2  gate1991(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1992(.a(s_206), .O(gate94inter3));
  inv1  gate1993(.a(s_207), .O(gate94inter4));
  nand2 gate1994(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1995(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1996(.a(G22), .O(gate94inter7));
  inv1  gate1997(.a(G344), .O(gate94inter8));
  nand2 gate1998(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1999(.a(s_207), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2000(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2001(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2002(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate701(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate702(.a(gate95inter0), .b(s_22), .O(gate95inter1));
  and2  gate703(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate704(.a(s_22), .O(gate95inter3));
  inv1  gate705(.a(s_23), .O(gate95inter4));
  nand2 gate706(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate707(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate708(.a(G26), .O(gate95inter7));
  inv1  gate709(.a(G347), .O(gate95inter8));
  nand2 gate710(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate711(.a(s_23), .b(gate95inter3), .O(gate95inter10));
  nor2  gate712(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate713(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate714(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate2479(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2480(.a(gate97inter0), .b(s_276), .O(gate97inter1));
  and2  gate2481(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2482(.a(s_276), .O(gate97inter3));
  inv1  gate2483(.a(s_277), .O(gate97inter4));
  nand2 gate2484(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2485(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2486(.a(G19), .O(gate97inter7));
  inv1  gate2487(.a(G350), .O(gate97inter8));
  nand2 gate2488(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2489(.a(s_277), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2490(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2491(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2492(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1569(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1570(.a(gate99inter0), .b(s_146), .O(gate99inter1));
  and2  gate1571(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1572(.a(s_146), .O(gate99inter3));
  inv1  gate1573(.a(s_147), .O(gate99inter4));
  nand2 gate1574(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1575(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1576(.a(G27), .O(gate99inter7));
  inv1  gate1577(.a(G353), .O(gate99inter8));
  nand2 gate1578(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1579(.a(s_147), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1580(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1581(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1582(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2787(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2788(.a(gate102inter0), .b(s_320), .O(gate102inter1));
  and2  gate2789(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2790(.a(s_320), .O(gate102inter3));
  inv1  gate2791(.a(s_321), .O(gate102inter4));
  nand2 gate2792(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2793(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2794(.a(G24), .O(gate102inter7));
  inv1  gate2795(.a(G356), .O(gate102inter8));
  nand2 gate2796(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2797(.a(s_321), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2798(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2799(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2800(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1891(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1892(.a(gate112inter0), .b(s_192), .O(gate112inter1));
  and2  gate1893(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1894(.a(s_192), .O(gate112inter3));
  inv1  gate1895(.a(s_193), .O(gate112inter4));
  nand2 gate1896(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1897(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1898(.a(G376), .O(gate112inter7));
  inv1  gate1899(.a(G377), .O(gate112inter8));
  nand2 gate1900(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1901(.a(s_193), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1902(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1903(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1904(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate589(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate590(.a(gate114inter0), .b(s_6), .O(gate114inter1));
  and2  gate591(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate592(.a(s_6), .O(gate114inter3));
  inv1  gate593(.a(s_7), .O(gate114inter4));
  nand2 gate594(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate595(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate596(.a(G380), .O(gate114inter7));
  inv1  gate597(.a(G381), .O(gate114inter8));
  nand2 gate598(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate599(.a(s_7), .b(gate114inter3), .O(gate114inter10));
  nor2  gate600(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate601(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate602(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate2857(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2858(.a(gate115inter0), .b(s_330), .O(gate115inter1));
  and2  gate2859(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2860(.a(s_330), .O(gate115inter3));
  inv1  gate2861(.a(s_331), .O(gate115inter4));
  nand2 gate2862(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2863(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2864(.a(G382), .O(gate115inter7));
  inv1  gate2865(.a(G383), .O(gate115inter8));
  nand2 gate2866(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2867(.a(s_331), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2868(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2869(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2870(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2829(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2830(.a(gate117inter0), .b(s_326), .O(gate117inter1));
  and2  gate2831(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2832(.a(s_326), .O(gate117inter3));
  inv1  gate2833(.a(s_327), .O(gate117inter4));
  nand2 gate2834(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2835(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2836(.a(G386), .O(gate117inter7));
  inv1  gate2837(.a(G387), .O(gate117inter8));
  nand2 gate2838(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2839(.a(s_327), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2840(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2841(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2842(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1051(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1052(.a(gate120inter0), .b(s_72), .O(gate120inter1));
  and2  gate1053(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1054(.a(s_72), .O(gate120inter3));
  inv1  gate1055(.a(s_73), .O(gate120inter4));
  nand2 gate1056(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1057(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1058(.a(G392), .O(gate120inter7));
  inv1  gate1059(.a(G393), .O(gate120inter8));
  nand2 gate1060(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1061(.a(s_73), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1062(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1063(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1064(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2227(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2228(.a(gate125inter0), .b(s_240), .O(gate125inter1));
  and2  gate2229(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2230(.a(s_240), .O(gate125inter3));
  inv1  gate2231(.a(s_241), .O(gate125inter4));
  nand2 gate2232(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2233(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2234(.a(G402), .O(gate125inter7));
  inv1  gate2235(.a(G403), .O(gate125inter8));
  nand2 gate2236(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2237(.a(s_241), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2238(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2239(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2240(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1653(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1654(.a(gate129inter0), .b(s_158), .O(gate129inter1));
  and2  gate1655(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1656(.a(s_158), .O(gate129inter3));
  inv1  gate1657(.a(s_159), .O(gate129inter4));
  nand2 gate1658(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1659(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1660(.a(G410), .O(gate129inter7));
  inv1  gate1661(.a(G411), .O(gate129inter8));
  nand2 gate1662(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1663(.a(s_159), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1664(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1665(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1666(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate2507(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2508(.a(gate133inter0), .b(s_280), .O(gate133inter1));
  and2  gate2509(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2510(.a(s_280), .O(gate133inter3));
  inv1  gate2511(.a(s_281), .O(gate133inter4));
  nand2 gate2512(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2513(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2514(.a(G418), .O(gate133inter7));
  inv1  gate2515(.a(G419), .O(gate133inter8));
  nand2 gate2516(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2517(.a(s_281), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2518(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2519(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2520(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1737(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1738(.a(gate134inter0), .b(s_170), .O(gate134inter1));
  and2  gate1739(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1740(.a(s_170), .O(gate134inter3));
  inv1  gate1741(.a(s_171), .O(gate134inter4));
  nand2 gate1742(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1743(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1744(.a(G420), .O(gate134inter7));
  inv1  gate1745(.a(G421), .O(gate134inter8));
  nand2 gate1746(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1747(.a(s_171), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1748(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1749(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1750(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1723(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1724(.a(gate136inter0), .b(s_168), .O(gate136inter1));
  and2  gate1725(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1726(.a(s_168), .O(gate136inter3));
  inv1  gate1727(.a(s_169), .O(gate136inter4));
  nand2 gate1728(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1729(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1730(.a(G424), .O(gate136inter7));
  inv1  gate1731(.a(G425), .O(gate136inter8));
  nand2 gate1732(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1733(.a(s_169), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1734(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1735(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1736(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1611(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1612(.a(gate138inter0), .b(s_152), .O(gate138inter1));
  and2  gate1613(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1614(.a(s_152), .O(gate138inter3));
  inv1  gate1615(.a(s_153), .O(gate138inter4));
  nand2 gate1616(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1617(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1618(.a(G432), .O(gate138inter7));
  inv1  gate1619(.a(G435), .O(gate138inter8));
  nand2 gate1620(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1621(.a(s_153), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1622(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1623(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1624(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate855(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate856(.a(gate139inter0), .b(s_44), .O(gate139inter1));
  and2  gate857(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate858(.a(s_44), .O(gate139inter3));
  inv1  gate859(.a(s_45), .O(gate139inter4));
  nand2 gate860(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate861(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate862(.a(G438), .O(gate139inter7));
  inv1  gate863(.a(G441), .O(gate139inter8));
  nand2 gate864(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate865(.a(s_45), .b(gate139inter3), .O(gate139inter10));
  nor2  gate866(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate867(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate868(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1527(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1528(.a(gate140inter0), .b(s_140), .O(gate140inter1));
  and2  gate1529(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1530(.a(s_140), .O(gate140inter3));
  inv1  gate1531(.a(s_141), .O(gate140inter4));
  nand2 gate1532(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1533(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1534(.a(G444), .O(gate140inter7));
  inv1  gate1535(.a(G447), .O(gate140inter8));
  nand2 gate1536(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1537(.a(s_141), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1538(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1539(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1540(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1205(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1206(.a(gate144inter0), .b(s_94), .O(gate144inter1));
  and2  gate1207(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1208(.a(s_94), .O(gate144inter3));
  inv1  gate1209(.a(s_95), .O(gate144inter4));
  nand2 gate1210(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1211(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1212(.a(G468), .O(gate144inter7));
  inv1  gate1213(.a(G471), .O(gate144inter8));
  nand2 gate1214(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1215(.a(s_95), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1216(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1217(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1218(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2003(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2004(.a(gate145inter0), .b(s_208), .O(gate145inter1));
  and2  gate2005(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2006(.a(s_208), .O(gate145inter3));
  inv1  gate2007(.a(s_209), .O(gate145inter4));
  nand2 gate2008(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2009(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2010(.a(G474), .O(gate145inter7));
  inv1  gate2011(.a(G477), .O(gate145inter8));
  nand2 gate2012(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2013(.a(s_209), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2014(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2015(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2016(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1163(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1164(.a(gate148inter0), .b(s_88), .O(gate148inter1));
  and2  gate1165(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1166(.a(s_88), .O(gate148inter3));
  inv1  gate1167(.a(s_89), .O(gate148inter4));
  nand2 gate1168(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1169(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1170(.a(G492), .O(gate148inter7));
  inv1  gate1171(.a(G495), .O(gate148inter8));
  nand2 gate1172(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1173(.a(s_89), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1174(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1175(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1176(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate995(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate996(.a(gate150inter0), .b(s_64), .O(gate150inter1));
  and2  gate997(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate998(.a(s_64), .O(gate150inter3));
  inv1  gate999(.a(s_65), .O(gate150inter4));
  nand2 gate1000(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1001(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1002(.a(G504), .O(gate150inter7));
  inv1  gate1003(.a(G507), .O(gate150inter8));
  nand2 gate1004(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1005(.a(s_65), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1006(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1007(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1008(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate785(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate786(.a(gate152inter0), .b(s_34), .O(gate152inter1));
  and2  gate787(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate788(.a(s_34), .O(gate152inter3));
  inv1  gate789(.a(s_35), .O(gate152inter4));
  nand2 gate790(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate791(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate792(.a(G516), .O(gate152inter7));
  inv1  gate793(.a(G519), .O(gate152inter8));
  nand2 gate794(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate795(.a(s_35), .b(gate152inter3), .O(gate152inter10));
  nor2  gate796(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate797(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate798(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate1597(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1598(.a(gate153inter0), .b(s_150), .O(gate153inter1));
  and2  gate1599(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1600(.a(s_150), .O(gate153inter3));
  inv1  gate1601(.a(s_151), .O(gate153inter4));
  nand2 gate1602(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1603(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1604(.a(G426), .O(gate153inter7));
  inv1  gate1605(.a(G522), .O(gate153inter8));
  nand2 gate1606(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1607(.a(s_151), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1608(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1609(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1610(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1359(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1360(.a(gate154inter0), .b(s_116), .O(gate154inter1));
  and2  gate1361(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1362(.a(s_116), .O(gate154inter3));
  inv1  gate1363(.a(s_117), .O(gate154inter4));
  nand2 gate1364(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1365(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1366(.a(G429), .O(gate154inter7));
  inv1  gate1367(.a(G522), .O(gate154inter8));
  nand2 gate1368(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1369(.a(s_117), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1370(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1371(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1372(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate2535(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2536(.a(gate156inter0), .b(s_284), .O(gate156inter1));
  and2  gate2537(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2538(.a(s_284), .O(gate156inter3));
  inv1  gate2539(.a(s_285), .O(gate156inter4));
  nand2 gate2540(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2541(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2542(.a(G435), .O(gate156inter7));
  inv1  gate2543(.a(G525), .O(gate156inter8));
  nand2 gate2544(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2545(.a(s_285), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2546(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2547(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2548(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2213(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2214(.a(gate157inter0), .b(s_238), .O(gate157inter1));
  and2  gate2215(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2216(.a(s_238), .O(gate157inter3));
  inv1  gate2217(.a(s_239), .O(gate157inter4));
  nand2 gate2218(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2219(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2220(.a(G438), .O(gate157inter7));
  inv1  gate2221(.a(G528), .O(gate157inter8));
  nand2 gate2222(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2223(.a(s_239), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2224(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2225(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2226(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1807(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1808(.a(gate160inter0), .b(s_180), .O(gate160inter1));
  and2  gate1809(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1810(.a(s_180), .O(gate160inter3));
  inv1  gate1811(.a(s_181), .O(gate160inter4));
  nand2 gate1812(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1813(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1814(.a(G447), .O(gate160inter7));
  inv1  gate1815(.a(G531), .O(gate160inter8));
  nand2 gate1816(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1817(.a(s_181), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1818(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1819(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1820(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1905(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1906(.a(gate162inter0), .b(s_194), .O(gate162inter1));
  and2  gate1907(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1908(.a(s_194), .O(gate162inter3));
  inv1  gate1909(.a(s_195), .O(gate162inter4));
  nand2 gate1910(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1911(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1912(.a(G453), .O(gate162inter7));
  inv1  gate1913(.a(G534), .O(gate162inter8));
  nand2 gate1914(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1915(.a(s_195), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1916(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1917(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1918(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2325(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2326(.a(gate163inter0), .b(s_254), .O(gate163inter1));
  and2  gate2327(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2328(.a(s_254), .O(gate163inter3));
  inv1  gate2329(.a(s_255), .O(gate163inter4));
  nand2 gate2330(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2331(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2332(.a(G456), .O(gate163inter7));
  inv1  gate2333(.a(G537), .O(gate163inter8));
  nand2 gate2334(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2335(.a(s_255), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2336(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2337(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2338(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate617(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate618(.a(gate164inter0), .b(s_10), .O(gate164inter1));
  and2  gate619(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate620(.a(s_10), .O(gate164inter3));
  inv1  gate621(.a(s_11), .O(gate164inter4));
  nand2 gate622(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate623(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate624(.a(G459), .O(gate164inter7));
  inv1  gate625(.a(G537), .O(gate164inter8));
  nand2 gate626(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate627(.a(s_11), .b(gate164inter3), .O(gate164inter10));
  nor2  gate628(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate629(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate630(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2073(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2074(.a(gate166inter0), .b(s_218), .O(gate166inter1));
  and2  gate2075(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2076(.a(s_218), .O(gate166inter3));
  inv1  gate2077(.a(s_219), .O(gate166inter4));
  nand2 gate2078(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2079(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2080(.a(G465), .O(gate166inter7));
  inv1  gate2081(.a(G540), .O(gate166inter8));
  nand2 gate2082(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2083(.a(s_219), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2084(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2085(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2086(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate2409(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate2410(.a(gate167inter0), .b(s_266), .O(gate167inter1));
  and2  gate2411(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate2412(.a(s_266), .O(gate167inter3));
  inv1  gate2413(.a(s_267), .O(gate167inter4));
  nand2 gate2414(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate2415(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate2416(.a(G468), .O(gate167inter7));
  inv1  gate2417(.a(G543), .O(gate167inter8));
  nand2 gate2418(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate2419(.a(s_267), .b(gate167inter3), .O(gate167inter10));
  nor2  gate2420(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate2421(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate2422(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate897(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate898(.a(gate173inter0), .b(s_50), .O(gate173inter1));
  and2  gate899(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate900(.a(s_50), .O(gate173inter3));
  inv1  gate901(.a(s_51), .O(gate173inter4));
  nand2 gate902(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate903(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate904(.a(G486), .O(gate173inter7));
  inv1  gate905(.a(G552), .O(gate173inter8));
  nand2 gate906(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate907(.a(s_51), .b(gate173inter3), .O(gate173inter10));
  nor2  gate908(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate909(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate910(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1583(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1584(.a(gate175inter0), .b(s_148), .O(gate175inter1));
  and2  gate1585(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1586(.a(s_148), .O(gate175inter3));
  inv1  gate1587(.a(s_149), .O(gate175inter4));
  nand2 gate1588(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1589(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1590(.a(G492), .O(gate175inter7));
  inv1  gate1591(.a(G555), .O(gate175inter8));
  nand2 gate1592(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1593(.a(s_149), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1594(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1595(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1596(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate2045(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2046(.a(gate176inter0), .b(s_214), .O(gate176inter1));
  and2  gate2047(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2048(.a(s_214), .O(gate176inter3));
  inv1  gate2049(.a(s_215), .O(gate176inter4));
  nand2 gate2050(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2051(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2052(.a(G495), .O(gate176inter7));
  inv1  gate2053(.a(G555), .O(gate176inter8));
  nand2 gate2054(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2055(.a(s_215), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2056(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2057(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2058(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate2619(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2620(.a(gate177inter0), .b(s_296), .O(gate177inter1));
  and2  gate2621(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2622(.a(s_296), .O(gate177inter3));
  inv1  gate2623(.a(s_297), .O(gate177inter4));
  nand2 gate2624(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2625(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2626(.a(G498), .O(gate177inter7));
  inv1  gate2627(.a(G558), .O(gate177inter8));
  nand2 gate2628(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2629(.a(s_297), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2630(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2631(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2632(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate2031(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2032(.a(gate178inter0), .b(s_212), .O(gate178inter1));
  and2  gate2033(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2034(.a(s_212), .O(gate178inter3));
  inv1  gate2035(.a(s_213), .O(gate178inter4));
  nand2 gate2036(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2037(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2038(.a(G501), .O(gate178inter7));
  inv1  gate2039(.a(G558), .O(gate178inter8));
  nand2 gate2040(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2041(.a(s_213), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2042(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2043(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2044(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate939(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate940(.a(gate184inter0), .b(s_56), .O(gate184inter1));
  and2  gate941(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate942(.a(s_56), .O(gate184inter3));
  inv1  gate943(.a(s_57), .O(gate184inter4));
  nand2 gate944(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate945(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate946(.a(G519), .O(gate184inter7));
  inv1  gate947(.a(G567), .O(gate184inter8));
  nand2 gate948(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate949(.a(s_57), .b(gate184inter3), .O(gate184inter10));
  nor2  gate950(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate951(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate952(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate2255(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2256(.a(gate186inter0), .b(s_244), .O(gate186inter1));
  and2  gate2257(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2258(.a(s_244), .O(gate186inter3));
  inv1  gate2259(.a(s_245), .O(gate186inter4));
  nand2 gate2260(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2261(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2262(.a(G572), .O(gate186inter7));
  inv1  gate2263(.a(G573), .O(gate186inter8));
  nand2 gate2264(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2265(.a(s_245), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2266(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2267(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2268(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1415(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1416(.a(gate189inter0), .b(s_124), .O(gate189inter1));
  and2  gate1417(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1418(.a(s_124), .O(gate189inter3));
  inv1  gate1419(.a(s_125), .O(gate189inter4));
  nand2 gate1420(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1421(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1422(.a(G578), .O(gate189inter7));
  inv1  gate1423(.a(G579), .O(gate189inter8));
  nand2 gate1424(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1425(.a(s_125), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1426(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1427(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1428(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1555(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1556(.a(gate191inter0), .b(s_144), .O(gate191inter1));
  and2  gate1557(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1558(.a(s_144), .O(gate191inter3));
  inv1  gate1559(.a(s_145), .O(gate191inter4));
  nand2 gate1560(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1561(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1562(.a(G582), .O(gate191inter7));
  inv1  gate1563(.a(G583), .O(gate191inter8));
  nand2 gate1564(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1565(.a(s_145), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1566(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1567(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1568(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1079(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1080(.a(gate194inter0), .b(s_76), .O(gate194inter1));
  and2  gate1081(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1082(.a(s_76), .O(gate194inter3));
  inv1  gate1083(.a(s_77), .O(gate194inter4));
  nand2 gate1084(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1085(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1086(.a(G588), .O(gate194inter7));
  inv1  gate1087(.a(G589), .O(gate194inter8));
  nand2 gate1088(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1089(.a(s_77), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1090(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1091(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1092(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1429(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1430(.a(gate195inter0), .b(s_126), .O(gate195inter1));
  and2  gate1431(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1432(.a(s_126), .O(gate195inter3));
  inv1  gate1433(.a(s_127), .O(gate195inter4));
  nand2 gate1434(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1435(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1436(.a(G590), .O(gate195inter7));
  inv1  gate1437(.a(G591), .O(gate195inter8));
  nand2 gate1438(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1439(.a(s_127), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1440(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1441(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1442(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate743(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate744(.a(gate197inter0), .b(s_28), .O(gate197inter1));
  and2  gate745(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate746(.a(s_28), .O(gate197inter3));
  inv1  gate747(.a(s_29), .O(gate197inter4));
  nand2 gate748(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate749(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate750(.a(G594), .O(gate197inter7));
  inv1  gate751(.a(G595), .O(gate197inter8));
  nand2 gate752(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate753(.a(s_29), .b(gate197inter3), .O(gate197inter10));
  nor2  gate754(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate755(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate756(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate883(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate884(.a(gate198inter0), .b(s_48), .O(gate198inter1));
  and2  gate885(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate886(.a(s_48), .O(gate198inter3));
  inv1  gate887(.a(s_49), .O(gate198inter4));
  nand2 gate888(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate889(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate890(.a(G596), .O(gate198inter7));
  inv1  gate891(.a(G597), .O(gate198inter8));
  nand2 gate892(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate893(.a(s_49), .b(gate198inter3), .O(gate198inter10));
  nor2  gate894(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate895(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate896(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1779(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1780(.a(gate199inter0), .b(s_176), .O(gate199inter1));
  and2  gate1781(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1782(.a(s_176), .O(gate199inter3));
  inv1  gate1783(.a(s_177), .O(gate199inter4));
  nand2 gate1784(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1785(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1786(.a(G598), .O(gate199inter7));
  inv1  gate1787(.a(G599), .O(gate199inter8));
  nand2 gate1788(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1789(.a(s_177), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1790(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1791(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1792(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1933(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1934(.a(gate200inter0), .b(s_198), .O(gate200inter1));
  and2  gate1935(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1936(.a(s_198), .O(gate200inter3));
  inv1  gate1937(.a(s_199), .O(gate200inter4));
  nand2 gate1938(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1939(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1940(.a(G600), .O(gate200inter7));
  inv1  gate1941(.a(G601), .O(gate200inter8));
  nand2 gate1942(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1943(.a(s_199), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1944(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1945(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1946(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate631(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate632(.a(gate203inter0), .b(s_12), .O(gate203inter1));
  and2  gate633(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate634(.a(s_12), .O(gate203inter3));
  inv1  gate635(.a(s_13), .O(gate203inter4));
  nand2 gate636(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate637(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate638(.a(G602), .O(gate203inter7));
  inv1  gate639(.a(G612), .O(gate203inter8));
  nand2 gate640(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate641(.a(s_13), .b(gate203inter3), .O(gate203inter10));
  nor2  gate642(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate643(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate644(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2087(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2088(.a(gate205inter0), .b(s_220), .O(gate205inter1));
  and2  gate2089(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2090(.a(s_220), .O(gate205inter3));
  inv1  gate2091(.a(s_221), .O(gate205inter4));
  nand2 gate2092(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2093(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2094(.a(G622), .O(gate205inter7));
  inv1  gate2095(.a(G627), .O(gate205inter8));
  nand2 gate2096(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2097(.a(s_221), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2098(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2099(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2100(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1149(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1150(.a(gate209inter0), .b(s_86), .O(gate209inter1));
  and2  gate1151(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1152(.a(s_86), .O(gate209inter3));
  inv1  gate1153(.a(s_87), .O(gate209inter4));
  nand2 gate1154(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1155(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1156(.a(G602), .O(gate209inter7));
  inv1  gate1157(.a(G666), .O(gate209inter8));
  nand2 gate1158(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1159(.a(s_87), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1160(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1161(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1162(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1443(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1444(.a(gate210inter0), .b(s_128), .O(gate210inter1));
  and2  gate1445(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1446(.a(s_128), .O(gate210inter3));
  inv1  gate1447(.a(s_129), .O(gate210inter4));
  nand2 gate1448(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1449(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1450(.a(G607), .O(gate210inter7));
  inv1  gate1451(.a(G666), .O(gate210inter8));
  nand2 gate1452(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1453(.a(s_129), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1454(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1455(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1456(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1765(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1766(.a(gate216inter0), .b(s_174), .O(gate216inter1));
  and2  gate1767(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1768(.a(s_174), .O(gate216inter3));
  inv1  gate1769(.a(s_175), .O(gate216inter4));
  nand2 gate1770(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1771(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1772(.a(G617), .O(gate216inter7));
  inv1  gate1773(.a(G675), .O(gate216inter8));
  nand2 gate1774(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1775(.a(s_175), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1776(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1777(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1778(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1107(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1108(.a(gate217inter0), .b(s_80), .O(gate217inter1));
  and2  gate1109(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1110(.a(s_80), .O(gate217inter3));
  inv1  gate1111(.a(s_81), .O(gate217inter4));
  nand2 gate1112(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1113(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1114(.a(G622), .O(gate217inter7));
  inv1  gate1115(.a(G678), .O(gate217inter8));
  nand2 gate1116(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1117(.a(s_81), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1118(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1119(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1120(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1457(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1458(.a(gate219inter0), .b(s_130), .O(gate219inter1));
  and2  gate1459(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1460(.a(s_130), .O(gate219inter3));
  inv1  gate1461(.a(s_131), .O(gate219inter4));
  nand2 gate1462(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1463(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1464(.a(G632), .O(gate219inter7));
  inv1  gate1465(.a(G681), .O(gate219inter8));
  nand2 gate1466(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1467(.a(s_131), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1468(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1469(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1470(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1387(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1388(.a(gate220inter0), .b(s_120), .O(gate220inter1));
  and2  gate1389(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1390(.a(s_120), .O(gate220inter3));
  inv1  gate1391(.a(s_121), .O(gate220inter4));
  nand2 gate1392(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1393(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1394(.a(G637), .O(gate220inter7));
  inv1  gate1395(.a(G681), .O(gate220inter8));
  nand2 gate1396(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1397(.a(s_121), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1398(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1399(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1400(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2311(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2312(.a(gate223inter0), .b(s_252), .O(gate223inter1));
  and2  gate2313(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2314(.a(s_252), .O(gate223inter3));
  inv1  gate2315(.a(s_253), .O(gate223inter4));
  nand2 gate2316(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2317(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2318(.a(G627), .O(gate223inter7));
  inv1  gate2319(.a(G687), .O(gate223inter8));
  nand2 gate2320(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2321(.a(s_253), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2322(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2323(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2324(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate967(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate968(.a(gate224inter0), .b(s_60), .O(gate224inter1));
  and2  gate969(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate970(.a(s_60), .O(gate224inter3));
  inv1  gate971(.a(s_61), .O(gate224inter4));
  nand2 gate972(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate973(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate974(.a(G637), .O(gate224inter7));
  inv1  gate975(.a(G687), .O(gate224inter8));
  nand2 gate976(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate977(.a(s_61), .b(gate224inter3), .O(gate224inter10));
  nor2  gate978(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate979(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate980(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1191(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1192(.a(gate226inter0), .b(s_92), .O(gate226inter1));
  and2  gate1193(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1194(.a(s_92), .O(gate226inter3));
  inv1  gate1195(.a(s_93), .O(gate226inter4));
  nand2 gate1196(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1197(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1198(.a(G692), .O(gate226inter7));
  inv1  gate1199(.a(G693), .O(gate226inter8));
  nand2 gate1200(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1201(.a(s_93), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1202(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1203(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1204(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2395(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2396(.a(gate231inter0), .b(s_264), .O(gate231inter1));
  and2  gate2397(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2398(.a(s_264), .O(gate231inter3));
  inv1  gate2399(.a(s_265), .O(gate231inter4));
  nand2 gate2400(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2401(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2402(.a(G702), .O(gate231inter7));
  inv1  gate2403(.a(G703), .O(gate231inter8));
  nand2 gate2404(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2405(.a(s_265), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2406(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2407(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2408(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate673(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate674(.a(gate232inter0), .b(s_18), .O(gate232inter1));
  and2  gate675(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate676(.a(s_18), .O(gate232inter3));
  inv1  gate677(.a(s_19), .O(gate232inter4));
  nand2 gate678(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate679(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate680(.a(G704), .O(gate232inter7));
  inv1  gate681(.a(G705), .O(gate232inter8));
  nand2 gate682(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate683(.a(s_19), .b(gate232inter3), .O(gate232inter10));
  nor2  gate684(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate685(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate686(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2381(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2382(.a(gate241inter0), .b(s_262), .O(gate241inter1));
  and2  gate2383(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2384(.a(s_262), .O(gate241inter3));
  inv1  gate2385(.a(s_263), .O(gate241inter4));
  nand2 gate2386(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2387(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2388(.a(G242), .O(gate241inter7));
  inv1  gate2389(.a(G730), .O(gate241inter8));
  nand2 gate2390(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2391(.a(s_263), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2392(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2393(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2394(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate2745(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2746(.a(gate244inter0), .b(s_314), .O(gate244inter1));
  and2  gate2747(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2748(.a(s_314), .O(gate244inter3));
  inv1  gate2749(.a(s_315), .O(gate244inter4));
  nand2 gate2750(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2751(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2752(.a(G721), .O(gate244inter7));
  inv1  gate2753(.a(G733), .O(gate244inter8));
  nand2 gate2754(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2755(.a(s_315), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2756(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2757(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2758(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate645(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate646(.a(gate246inter0), .b(s_14), .O(gate246inter1));
  and2  gate647(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate648(.a(s_14), .O(gate246inter3));
  inv1  gate649(.a(s_15), .O(gate246inter4));
  nand2 gate650(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate651(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate652(.a(G724), .O(gate246inter7));
  inv1  gate653(.a(G736), .O(gate246inter8));
  nand2 gate654(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate655(.a(s_15), .b(gate246inter3), .O(gate246inter10));
  nor2  gate656(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate657(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate658(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2647(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2648(.a(gate250inter0), .b(s_300), .O(gate250inter1));
  and2  gate2649(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2650(.a(s_300), .O(gate250inter3));
  inv1  gate2651(.a(s_301), .O(gate250inter4));
  nand2 gate2652(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2653(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2654(.a(G706), .O(gate250inter7));
  inv1  gate2655(.a(G742), .O(gate250inter8));
  nand2 gate2656(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2657(.a(s_301), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2658(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2659(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2660(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2465(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2466(.a(gate251inter0), .b(s_274), .O(gate251inter1));
  and2  gate2467(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2468(.a(s_274), .O(gate251inter3));
  inv1  gate2469(.a(s_275), .O(gate251inter4));
  nand2 gate2470(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2471(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2472(.a(G257), .O(gate251inter7));
  inv1  gate2473(.a(G745), .O(gate251inter8));
  nand2 gate2474(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2475(.a(s_275), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2476(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2477(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2478(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1317(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1318(.a(gate253inter0), .b(s_110), .O(gate253inter1));
  and2  gate1319(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1320(.a(s_110), .O(gate253inter3));
  inv1  gate1321(.a(s_111), .O(gate253inter4));
  nand2 gate1322(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1323(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1324(.a(G260), .O(gate253inter7));
  inv1  gate1325(.a(G748), .O(gate253inter8));
  nand2 gate1326(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1327(.a(s_111), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1328(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1329(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1330(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1023(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1024(.a(gate254inter0), .b(s_68), .O(gate254inter1));
  and2  gate1025(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1026(.a(s_68), .O(gate254inter3));
  inv1  gate1027(.a(s_69), .O(gate254inter4));
  nand2 gate1028(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1029(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1030(.a(G712), .O(gate254inter7));
  inv1  gate1031(.a(G748), .O(gate254inter8));
  nand2 gate1032(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1033(.a(s_69), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1034(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1035(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1036(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate2115(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2116(.a(gate255inter0), .b(s_224), .O(gate255inter1));
  and2  gate2117(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2118(.a(s_224), .O(gate255inter3));
  inv1  gate2119(.a(s_225), .O(gate255inter4));
  nand2 gate2120(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2121(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2122(.a(G263), .O(gate255inter7));
  inv1  gate2123(.a(G751), .O(gate255inter8));
  nand2 gate2124(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2125(.a(s_225), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2126(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2127(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2128(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1975(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1976(.a(gate256inter0), .b(s_204), .O(gate256inter1));
  and2  gate1977(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1978(.a(s_204), .O(gate256inter3));
  inv1  gate1979(.a(s_205), .O(gate256inter4));
  nand2 gate1980(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1981(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1982(.a(G715), .O(gate256inter7));
  inv1  gate1983(.a(G751), .O(gate256inter8));
  nand2 gate1984(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1985(.a(s_205), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1986(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1987(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1988(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate2521(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2522(.a(gate259inter0), .b(s_282), .O(gate259inter1));
  and2  gate2523(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2524(.a(s_282), .O(gate259inter3));
  inv1  gate2525(.a(s_283), .O(gate259inter4));
  nand2 gate2526(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2527(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2528(.a(G758), .O(gate259inter7));
  inv1  gate2529(.a(G759), .O(gate259inter8));
  nand2 gate2530(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2531(.a(s_283), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2532(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2533(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2534(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2773(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2774(.a(gate262inter0), .b(s_318), .O(gate262inter1));
  and2  gate2775(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2776(.a(s_318), .O(gate262inter3));
  inv1  gate2777(.a(s_319), .O(gate262inter4));
  nand2 gate2778(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2779(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2780(.a(G764), .O(gate262inter7));
  inv1  gate2781(.a(G765), .O(gate262inter8));
  nand2 gate2782(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2783(.a(s_319), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2784(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2785(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2786(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2661(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2662(.a(gate264inter0), .b(s_302), .O(gate264inter1));
  and2  gate2663(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2664(.a(s_302), .O(gate264inter3));
  inv1  gate2665(.a(s_303), .O(gate264inter4));
  nand2 gate2666(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2667(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2668(.a(G768), .O(gate264inter7));
  inv1  gate2669(.a(G769), .O(gate264inter8));
  nand2 gate2670(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2671(.a(s_303), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2672(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2673(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2674(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1667(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1668(.a(gate266inter0), .b(s_160), .O(gate266inter1));
  and2  gate1669(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1670(.a(s_160), .O(gate266inter3));
  inv1  gate1671(.a(s_161), .O(gate266inter4));
  nand2 gate1672(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1673(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1674(.a(G645), .O(gate266inter7));
  inv1  gate1675(.a(G773), .O(gate266inter8));
  nand2 gate1676(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1677(.a(s_161), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1678(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1679(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1680(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate827(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate828(.a(gate269inter0), .b(s_40), .O(gate269inter1));
  and2  gate829(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate830(.a(s_40), .O(gate269inter3));
  inv1  gate831(.a(s_41), .O(gate269inter4));
  nand2 gate832(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate833(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate834(.a(G654), .O(gate269inter7));
  inv1  gate835(.a(G782), .O(gate269inter8));
  nand2 gate836(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate837(.a(s_41), .b(gate269inter3), .O(gate269inter10));
  nor2  gate838(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate839(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate840(.a(gate269inter12), .b(gate269inter1), .O(G806));

  xor2  gate2241(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2242(.a(gate270inter0), .b(s_242), .O(gate270inter1));
  and2  gate2243(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2244(.a(s_242), .O(gate270inter3));
  inv1  gate2245(.a(s_243), .O(gate270inter4));
  nand2 gate2246(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2247(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2248(.a(G657), .O(gate270inter7));
  inv1  gate2249(.a(G785), .O(gate270inter8));
  nand2 gate2250(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2251(.a(s_243), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2252(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2253(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2254(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2423(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2424(.a(gate274inter0), .b(s_268), .O(gate274inter1));
  and2  gate2425(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2426(.a(s_268), .O(gate274inter3));
  inv1  gate2427(.a(s_269), .O(gate274inter4));
  nand2 gate2428(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2429(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2430(.a(G770), .O(gate274inter7));
  inv1  gate2431(.a(G794), .O(gate274inter8));
  nand2 gate2432(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2433(.a(s_269), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2434(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2435(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2436(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2185(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2186(.a(gate278inter0), .b(s_234), .O(gate278inter1));
  and2  gate2187(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2188(.a(s_234), .O(gate278inter3));
  inv1  gate2189(.a(s_235), .O(gate278inter4));
  nand2 gate2190(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2191(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2192(.a(G776), .O(gate278inter7));
  inv1  gate2193(.a(G800), .O(gate278inter8));
  nand2 gate2194(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2195(.a(s_235), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2196(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2197(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2198(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1821(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1822(.a(gate279inter0), .b(s_182), .O(gate279inter1));
  and2  gate1823(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1824(.a(s_182), .O(gate279inter3));
  inv1  gate1825(.a(s_183), .O(gate279inter4));
  nand2 gate1826(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1827(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1828(.a(G651), .O(gate279inter7));
  inv1  gate1829(.a(G803), .O(gate279inter8));
  nand2 gate1830(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1831(.a(s_183), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1832(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1833(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1834(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate981(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate982(.a(gate280inter0), .b(s_62), .O(gate280inter1));
  and2  gate983(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate984(.a(s_62), .O(gate280inter3));
  inv1  gate985(.a(s_63), .O(gate280inter4));
  nand2 gate986(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate987(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate988(.a(G779), .O(gate280inter7));
  inv1  gate989(.a(G803), .O(gate280inter8));
  nand2 gate990(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate991(.a(s_63), .b(gate280inter3), .O(gate280inter10));
  nor2  gate992(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate993(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate994(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1625(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1626(.a(gate281inter0), .b(s_154), .O(gate281inter1));
  and2  gate1627(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1628(.a(s_154), .O(gate281inter3));
  inv1  gate1629(.a(s_155), .O(gate281inter4));
  nand2 gate1630(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1631(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1632(.a(G654), .O(gate281inter7));
  inv1  gate1633(.a(G806), .O(gate281inter8));
  nand2 gate1634(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1635(.a(s_155), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1636(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1637(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1638(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1373(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1374(.a(gate286inter0), .b(s_118), .O(gate286inter1));
  and2  gate1375(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1376(.a(s_118), .O(gate286inter3));
  inv1  gate1377(.a(s_119), .O(gate286inter4));
  nand2 gate1378(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1379(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1380(.a(G788), .O(gate286inter7));
  inv1  gate1381(.a(G812), .O(gate286inter8));
  nand2 gate1382(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1383(.a(s_119), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1384(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1385(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1386(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate841(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate842(.a(gate287inter0), .b(s_42), .O(gate287inter1));
  and2  gate843(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate844(.a(s_42), .O(gate287inter3));
  inv1  gate845(.a(s_43), .O(gate287inter4));
  nand2 gate846(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate847(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate848(.a(G663), .O(gate287inter7));
  inv1  gate849(.a(G815), .O(gate287inter8));
  nand2 gate850(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate851(.a(s_43), .b(gate287inter3), .O(gate287inter10));
  nor2  gate852(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate853(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate854(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1849(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1850(.a(gate288inter0), .b(s_186), .O(gate288inter1));
  and2  gate1851(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1852(.a(s_186), .O(gate288inter3));
  inv1  gate1853(.a(s_187), .O(gate288inter4));
  nand2 gate1854(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1855(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1856(.a(G791), .O(gate288inter7));
  inv1  gate1857(.a(G815), .O(gate288inter8));
  nand2 gate1858(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1859(.a(s_187), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1860(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1861(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1862(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate869(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate870(.a(gate289inter0), .b(s_46), .O(gate289inter1));
  and2  gate871(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate872(.a(s_46), .O(gate289inter3));
  inv1  gate873(.a(s_47), .O(gate289inter4));
  nand2 gate874(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate875(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate876(.a(G818), .O(gate289inter7));
  inv1  gate877(.a(G819), .O(gate289inter8));
  nand2 gate878(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate879(.a(s_47), .b(gate289inter3), .O(gate289inter10));
  nor2  gate880(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate881(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate882(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2703(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2704(.a(gate389inter0), .b(s_308), .O(gate389inter1));
  and2  gate2705(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2706(.a(s_308), .O(gate389inter3));
  inv1  gate2707(.a(s_309), .O(gate389inter4));
  nand2 gate2708(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2709(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2710(.a(G3), .O(gate389inter7));
  inv1  gate2711(.a(G1042), .O(gate389inter8));
  nand2 gate2712(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2713(.a(s_309), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2714(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2715(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2716(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1681(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1682(.a(gate393inter0), .b(s_162), .O(gate393inter1));
  and2  gate1683(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1684(.a(s_162), .O(gate393inter3));
  inv1  gate1685(.a(s_163), .O(gate393inter4));
  nand2 gate1686(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1687(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1688(.a(G7), .O(gate393inter7));
  inv1  gate1689(.a(G1054), .O(gate393inter8));
  nand2 gate1690(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1691(.a(s_163), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1692(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1693(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1694(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2297(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2298(.a(gate395inter0), .b(s_250), .O(gate395inter1));
  and2  gate2299(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2300(.a(s_250), .O(gate395inter3));
  inv1  gate2301(.a(s_251), .O(gate395inter4));
  nand2 gate2302(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2303(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2304(.a(G9), .O(gate395inter7));
  inv1  gate2305(.a(G1060), .O(gate395inter8));
  nand2 gate2306(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2307(.a(s_251), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2308(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2309(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2310(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2451(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2452(.a(gate398inter0), .b(s_272), .O(gate398inter1));
  and2  gate2453(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2454(.a(s_272), .O(gate398inter3));
  inv1  gate2455(.a(s_273), .O(gate398inter4));
  nand2 gate2456(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2457(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2458(.a(G12), .O(gate398inter7));
  inv1  gate2459(.a(G1069), .O(gate398inter8));
  nand2 gate2460(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2461(.a(s_273), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2462(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2463(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2464(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2129(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2130(.a(gate402inter0), .b(s_226), .O(gate402inter1));
  and2  gate2131(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2132(.a(s_226), .O(gate402inter3));
  inv1  gate2133(.a(s_227), .O(gate402inter4));
  nand2 gate2134(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2135(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2136(.a(G16), .O(gate402inter7));
  inv1  gate2137(.a(G1081), .O(gate402inter8));
  nand2 gate2138(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2139(.a(s_227), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2140(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2141(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2142(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2143(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2144(.a(gate406inter0), .b(s_228), .O(gate406inter1));
  and2  gate2145(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2146(.a(s_228), .O(gate406inter3));
  inv1  gate2147(.a(s_229), .O(gate406inter4));
  nand2 gate2148(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2149(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2150(.a(G20), .O(gate406inter7));
  inv1  gate2151(.a(G1093), .O(gate406inter8));
  nand2 gate2152(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2153(.a(s_229), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2154(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2155(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2156(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate911(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate912(.a(gate408inter0), .b(s_52), .O(gate408inter1));
  and2  gate913(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate914(.a(s_52), .O(gate408inter3));
  inv1  gate915(.a(s_53), .O(gate408inter4));
  nand2 gate916(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate917(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate918(.a(G22), .O(gate408inter7));
  inv1  gate919(.a(G1099), .O(gate408inter8));
  nand2 gate920(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate921(.a(s_53), .b(gate408inter3), .O(gate408inter10));
  nor2  gate922(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate923(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate924(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate2101(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2102(.a(gate409inter0), .b(s_222), .O(gate409inter1));
  and2  gate2103(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2104(.a(s_222), .O(gate409inter3));
  inv1  gate2105(.a(s_223), .O(gate409inter4));
  nand2 gate2106(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2107(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2108(.a(G23), .O(gate409inter7));
  inv1  gate2109(.a(G1102), .O(gate409inter8));
  nand2 gate2110(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2111(.a(s_223), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2112(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2113(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2114(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate575(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate576(.a(gate411inter0), .b(s_4), .O(gate411inter1));
  and2  gate577(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate578(.a(s_4), .O(gate411inter3));
  inv1  gate579(.a(s_5), .O(gate411inter4));
  nand2 gate580(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate581(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate582(.a(G25), .O(gate411inter7));
  inv1  gate583(.a(G1108), .O(gate411inter8));
  nand2 gate584(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate585(.a(s_5), .b(gate411inter3), .O(gate411inter10));
  nor2  gate586(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate587(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate588(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate771(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate772(.a(gate418inter0), .b(s_32), .O(gate418inter1));
  and2  gate773(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate774(.a(s_32), .O(gate418inter3));
  inv1  gate775(.a(s_33), .O(gate418inter4));
  nand2 gate776(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate777(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate778(.a(G32), .O(gate418inter7));
  inv1  gate779(.a(G1129), .O(gate418inter8));
  nand2 gate780(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate781(.a(s_33), .b(gate418inter3), .O(gate418inter10));
  nor2  gate782(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate783(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate784(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1121(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1122(.a(gate419inter0), .b(s_82), .O(gate419inter1));
  and2  gate1123(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1124(.a(s_82), .O(gate419inter3));
  inv1  gate1125(.a(s_83), .O(gate419inter4));
  nand2 gate1126(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1127(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1128(.a(G1), .O(gate419inter7));
  inv1  gate1129(.a(G1132), .O(gate419inter8));
  nand2 gate1130(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1131(.a(s_83), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1132(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1133(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1134(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1863(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1864(.a(gate420inter0), .b(s_188), .O(gate420inter1));
  and2  gate1865(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1866(.a(s_188), .O(gate420inter3));
  inv1  gate1867(.a(s_189), .O(gate420inter4));
  nand2 gate1868(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1869(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1870(.a(G1036), .O(gate420inter7));
  inv1  gate1871(.a(G1132), .O(gate420inter8));
  nand2 gate1872(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1873(.a(s_189), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1874(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1875(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1876(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate2759(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2760(.a(gate423inter0), .b(s_316), .O(gate423inter1));
  and2  gate2761(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2762(.a(s_316), .O(gate423inter3));
  inv1  gate2763(.a(s_317), .O(gate423inter4));
  nand2 gate2764(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2765(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2766(.a(G3), .O(gate423inter7));
  inv1  gate2767(.a(G1138), .O(gate423inter8));
  nand2 gate2768(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2769(.a(s_317), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2770(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2771(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2772(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate953(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate954(.a(gate426inter0), .b(s_58), .O(gate426inter1));
  and2  gate955(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate956(.a(s_58), .O(gate426inter3));
  inv1  gate957(.a(s_59), .O(gate426inter4));
  nand2 gate958(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate959(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate960(.a(G1045), .O(gate426inter7));
  inv1  gate961(.a(G1141), .O(gate426inter8));
  nand2 gate962(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate963(.a(s_59), .b(gate426inter3), .O(gate426inter10));
  nor2  gate964(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate965(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate966(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate561(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate562(.a(gate428inter0), .b(s_2), .O(gate428inter1));
  and2  gate563(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate564(.a(s_2), .O(gate428inter3));
  inv1  gate565(.a(s_3), .O(gate428inter4));
  nand2 gate566(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate567(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate568(.a(G1048), .O(gate428inter7));
  inv1  gate569(.a(G1144), .O(gate428inter8));
  nand2 gate570(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate571(.a(s_3), .b(gate428inter3), .O(gate428inter10));
  nor2  gate572(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate573(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate574(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate2577(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2578(.a(gate429inter0), .b(s_290), .O(gate429inter1));
  and2  gate2579(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2580(.a(s_290), .O(gate429inter3));
  inv1  gate2581(.a(s_291), .O(gate429inter4));
  nand2 gate2582(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2583(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2584(.a(G6), .O(gate429inter7));
  inv1  gate2585(.a(G1147), .O(gate429inter8));
  nand2 gate2586(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2587(.a(s_291), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2588(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2589(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2590(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate687(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate688(.a(gate436inter0), .b(s_20), .O(gate436inter1));
  and2  gate689(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate690(.a(s_20), .O(gate436inter3));
  inv1  gate691(.a(s_21), .O(gate436inter4));
  nand2 gate692(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate693(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate694(.a(G1060), .O(gate436inter7));
  inv1  gate695(.a(G1156), .O(gate436inter8));
  nand2 gate696(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate697(.a(s_21), .b(gate436inter3), .O(gate436inter10));
  nor2  gate698(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate699(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate700(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate2437(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2438(.a(gate440inter0), .b(s_270), .O(gate440inter1));
  and2  gate2439(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2440(.a(s_270), .O(gate440inter3));
  inv1  gate2441(.a(s_271), .O(gate440inter4));
  nand2 gate2442(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2443(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2444(.a(G1066), .O(gate440inter7));
  inv1  gate2445(.a(G1162), .O(gate440inter8));
  nand2 gate2446(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2447(.a(s_271), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2448(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2449(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2450(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1947(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1948(.a(gate441inter0), .b(s_200), .O(gate441inter1));
  and2  gate1949(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1950(.a(s_200), .O(gate441inter3));
  inv1  gate1951(.a(s_201), .O(gate441inter4));
  nand2 gate1952(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1953(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1954(.a(G12), .O(gate441inter7));
  inv1  gate1955(.a(G1165), .O(gate441inter8));
  nand2 gate1956(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1957(.a(s_201), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1958(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1959(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1960(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1219(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1220(.a(gate442inter0), .b(s_96), .O(gate442inter1));
  and2  gate1221(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1222(.a(s_96), .O(gate442inter3));
  inv1  gate1223(.a(s_97), .O(gate442inter4));
  nand2 gate1224(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1225(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1226(.a(G1069), .O(gate442inter7));
  inv1  gate1227(.a(G1165), .O(gate442inter8));
  nand2 gate1228(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1229(.a(s_97), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1230(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1231(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1232(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1639(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1640(.a(gate443inter0), .b(s_156), .O(gate443inter1));
  and2  gate1641(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1642(.a(s_156), .O(gate443inter3));
  inv1  gate1643(.a(s_157), .O(gate443inter4));
  nand2 gate1644(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1645(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1646(.a(G13), .O(gate443inter7));
  inv1  gate1647(.a(G1168), .O(gate443inter8));
  nand2 gate1648(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1649(.a(s_157), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1650(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1651(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1652(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2059(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2060(.a(gate445inter0), .b(s_216), .O(gate445inter1));
  and2  gate2061(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2062(.a(s_216), .O(gate445inter3));
  inv1  gate2063(.a(s_217), .O(gate445inter4));
  nand2 gate2064(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2065(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2066(.a(G14), .O(gate445inter7));
  inv1  gate2067(.a(G1171), .O(gate445inter8));
  nand2 gate2068(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2069(.a(s_217), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2070(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2071(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2072(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate2171(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2172(.a(gate446inter0), .b(s_232), .O(gate446inter1));
  and2  gate2173(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2174(.a(s_232), .O(gate446inter3));
  inv1  gate2175(.a(s_233), .O(gate446inter4));
  nand2 gate2176(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2177(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2178(.a(G1075), .O(gate446inter7));
  inv1  gate2179(.a(G1171), .O(gate446inter8));
  nand2 gate2180(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2181(.a(s_233), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2182(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2183(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2184(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1485(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1486(.a(gate449inter0), .b(s_134), .O(gate449inter1));
  and2  gate1487(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1488(.a(s_134), .O(gate449inter3));
  inv1  gate1489(.a(s_135), .O(gate449inter4));
  nand2 gate1490(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1491(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1492(.a(G16), .O(gate449inter7));
  inv1  gate1493(.a(G1177), .O(gate449inter8));
  nand2 gate1494(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1495(.a(s_135), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1496(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1497(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1498(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1093(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1094(.a(gate452inter0), .b(s_78), .O(gate452inter1));
  and2  gate1095(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1096(.a(s_78), .O(gate452inter3));
  inv1  gate1097(.a(s_79), .O(gate452inter4));
  nand2 gate1098(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1099(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1100(.a(G1084), .O(gate452inter7));
  inv1  gate1101(.a(G1180), .O(gate452inter8));
  nand2 gate1102(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1103(.a(s_79), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1104(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1105(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1106(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2269(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2270(.a(gate455inter0), .b(s_246), .O(gate455inter1));
  and2  gate2271(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2272(.a(s_246), .O(gate455inter3));
  inv1  gate2273(.a(s_247), .O(gate455inter4));
  nand2 gate2274(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2275(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2276(.a(G19), .O(gate455inter7));
  inv1  gate2277(.a(G1186), .O(gate455inter8));
  nand2 gate2278(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2279(.a(s_247), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2280(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2281(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2282(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1835(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1836(.a(gate456inter0), .b(s_184), .O(gate456inter1));
  and2  gate1837(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1838(.a(s_184), .O(gate456inter3));
  inv1  gate1839(.a(s_185), .O(gate456inter4));
  nand2 gate1840(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1841(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1842(.a(G1090), .O(gate456inter7));
  inv1  gate1843(.a(G1186), .O(gate456inter8));
  nand2 gate1844(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1845(.a(s_185), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1846(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1847(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1848(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2815(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2816(.a(gate460inter0), .b(s_324), .O(gate460inter1));
  and2  gate2817(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2818(.a(s_324), .O(gate460inter3));
  inv1  gate2819(.a(s_325), .O(gate460inter4));
  nand2 gate2820(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2821(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2822(.a(G1096), .O(gate460inter7));
  inv1  gate2823(.a(G1192), .O(gate460inter8));
  nand2 gate2824(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2825(.a(s_325), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2826(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2827(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2828(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2017(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2018(.a(gate461inter0), .b(s_210), .O(gate461inter1));
  and2  gate2019(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2020(.a(s_210), .O(gate461inter3));
  inv1  gate2021(.a(s_211), .O(gate461inter4));
  nand2 gate2022(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2023(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2024(.a(G22), .O(gate461inter7));
  inv1  gate2025(.a(G1195), .O(gate461inter8));
  nand2 gate2026(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2027(.a(s_211), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2028(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2029(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2030(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1331(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1332(.a(gate463inter0), .b(s_112), .O(gate463inter1));
  and2  gate1333(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1334(.a(s_112), .O(gate463inter3));
  inv1  gate1335(.a(s_113), .O(gate463inter4));
  nand2 gate1336(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1337(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1338(.a(G23), .O(gate463inter7));
  inv1  gate1339(.a(G1198), .O(gate463inter8));
  nand2 gate1340(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1341(.a(s_113), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1342(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1343(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1344(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate799(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate800(.a(gate464inter0), .b(s_36), .O(gate464inter1));
  and2  gate801(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate802(.a(s_36), .O(gate464inter3));
  inv1  gate803(.a(s_37), .O(gate464inter4));
  nand2 gate804(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate805(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate806(.a(G1102), .O(gate464inter7));
  inv1  gate807(.a(G1198), .O(gate464inter8));
  nand2 gate808(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate809(.a(s_37), .b(gate464inter3), .O(gate464inter10));
  nor2  gate810(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate811(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate812(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1065(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1066(.a(gate465inter0), .b(s_74), .O(gate465inter1));
  and2  gate1067(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1068(.a(s_74), .O(gate465inter3));
  inv1  gate1069(.a(s_75), .O(gate465inter4));
  nand2 gate1070(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1071(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1072(.a(G24), .O(gate465inter7));
  inv1  gate1073(.a(G1201), .O(gate465inter8));
  nand2 gate1074(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1075(.a(s_75), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1076(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1077(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1078(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2605(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2606(.a(gate466inter0), .b(s_294), .O(gate466inter1));
  and2  gate2607(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2608(.a(s_294), .O(gate466inter3));
  inv1  gate2609(.a(s_295), .O(gate466inter4));
  nand2 gate2610(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2611(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2612(.a(G1105), .O(gate466inter7));
  inv1  gate2613(.a(G1201), .O(gate466inter8));
  nand2 gate2614(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2615(.a(s_295), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2616(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2617(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2618(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1009(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1010(.a(gate467inter0), .b(s_66), .O(gate467inter1));
  and2  gate1011(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1012(.a(s_66), .O(gate467inter3));
  inv1  gate1013(.a(s_67), .O(gate467inter4));
  nand2 gate1014(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1015(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1016(.a(G25), .O(gate467inter7));
  inv1  gate1017(.a(G1204), .O(gate467inter8));
  nand2 gate1018(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1019(.a(s_67), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1020(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1021(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1022(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1275(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1276(.a(gate472inter0), .b(s_104), .O(gate472inter1));
  and2  gate1277(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1278(.a(s_104), .O(gate472inter3));
  inv1  gate1279(.a(s_105), .O(gate472inter4));
  nand2 gate1280(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1281(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1282(.a(G1114), .O(gate472inter7));
  inv1  gate1283(.a(G1210), .O(gate472inter8));
  nand2 gate1284(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1285(.a(s_105), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1286(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1287(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1288(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1793(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1794(.a(gate474inter0), .b(s_178), .O(gate474inter1));
  and2  gate1795(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1796(.a(s_178), .O(gate474inter3));
  inv1  gate1797(.a(s_179), .O(gate474inter4));
  nand2 gate1798(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1799(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1800(.a(G1117), .O(gate474inter7));
  inv1  gate1801(.a(G1213), .O(gate474inter8));
  nand2 gate1802(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1803(.a(s_179), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1804(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1805(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1806(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2549(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2550(.a(gate482inter0), .b(s_286), .O(gate482inter1));
  and2  gate2551(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2552(.a(s_286), .O(gate482inter3));
  inv1  gate2553(.a(s_287), .O(gate482inter4));
  nand2 gate2554(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2555(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2556(.a(G1129), .O(gate482inter7));
  inv1  gate2557(.a(G1225), .O(gate482inter8));
  nand2 gate2558(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2559(.a(s_287), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2560(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2561(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2562(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1919(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1920(.a(gate483inter0), .b(s_196), .O(gate483inter1));
  and2  gate1921(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1922(.a(s_196), .O(gate483inter3));
  inv1  gate1923(.a(s_197), .O(gate483inter4));
  nand2 gate1924(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1925(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1926(.a(G1228), .O(gate483inter7));
  inv1  gate1927(.a(G1229), .O(gate483inter8));
  nand2 gate1928(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1929(.a(s_197), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1930(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1931(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1932(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1513(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1514(.a(gate485inter0), .b(s_138), .O(gate485inter1));
  and2  gate1515(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1516(.a(s_138), .O(gate485inter3));
  inv1  gate1517(.a(s_139), .O(gate485inter4));
  nand2 gate1518(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1519(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1520(.a(G1232), .O(gate485inter7));
  inv1  gate1521(.a(G1233), .O(gate485inter8));
  nand2 gate1522(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1523(.a(s_139), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1524(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1525(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1526(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate603(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate604(.a(gate486inter0), .b(s_8), .O(gate486inter1));
  and2  gate605(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate606(.a(s_8), .O(gate486inter3));
  inv1  gate607(.a(s_9), .O(gate486inter4));
  nand2 gate608(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate609(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate610(.a(G1234), .O(gate486inter7));
  inv1  gate611(.a(G1235), .O(gate486inter8));
  nand2 gate612(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate613(.a(s_9), .b(gate486inter3), .O(gate486inter10));
  nor2  gate614(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate615(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate616(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2339(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2340(.a(gate487inter0), .b(s_256), .O(gate487inter1));
  and2  gate2341(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2342(.a(s_256), .O(gate487inter3));
  inv1  gate2343(.a(s_257), .O(gate487inter4));
  nand2 gate2344(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2345(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2346(.a(G1236), .O(gate487inter7));
  inv1  gate2347(.a(G1237), .O(gate487inter8));
  nand2 gate2348(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2349(.a(s_257), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2350(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2351(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2352(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1541(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1542(.a(gate488inter0), .b(s_142), .O(gate488inter1));
  and2  gate1543(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1544(.a(s_142), .O(gate488inter3));
  inv1  gate1545(.a(s_143), .O(gate488inter4));
  nand2 gate1546(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1547(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1548(.a(G1238), .O(gate488inter7));
  inv1  gate1549(.a(G1239), .O(gate488inter8));
  nand2 gate1550(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1551(.a(s_143), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1552(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1553(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1554(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate2731(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2732(.a(gate494inter0), .b(s_312), .O(gate494inter1));
  and2  gate2733(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2734(.a(s_312), .O(gate494inter3));
  inv1  gate2735(.a(s_313), .O(gate494inter4));
  nand2 gate2736(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2737(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2738(.a(G1250), .O(gate494inter7));
  inv1  gate2739(.a(G1251), .O(gate494inter8));
  nand2 gate2740(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2741(.a(s_313), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2742(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2743(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2744(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2199(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2200(.a(gate495inter0), .b(s_236), .O(gate495inter1));
  and2  gate2201(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2202(.a(s_236), .O(gate495inter3));
  inv1  gate2203(.a(s_237), .O(gate495inter4));
  nand2 gate2204(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2205(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2206(.a(G1252), .O(gate495inter7));
  inv1  gate2207(.a(G1253), .O(gate495inter8));
  nand2 gate2208(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2209(.a(s_237), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2210(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2211(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2212(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1695(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1696(.a(gate502inter0), .b(s_164), .O(gate502inter1));
  and2  gate1697(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1698(.a(s_164), .O(gate502inter3));
  inv1  gate1699(.a(s_165), .O(gate502inter4));
  nand2 gate1700(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1701(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1702(.a(G1266), .O(gate502inter7));
  inv1  gate1703(.a(G1267), .O(gate502inter8));
  nand2 gate1704(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1705(.a(s_165), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1706(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1707(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1708(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2633(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2634(.a(gate503inter0), .b(s_298), .O(gate503inter1));
  and2  gate2635(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2636(.a(s_298), .O(gate503inter3));
  inv1  gate2637(.a(s_299), .O(gate503inter4));
  nand2 gate2638(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2639(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2640(.a(G1268), .O(gate503inter7));
  inv1  gate2641(.a(G1269), .O(gate503inter8));
  nand2 gate2642(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2643(.a(s_299), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2644(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2645(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2646(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate2843(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2844(.a(gate506inter0), .b(s_328), .O(gate506inter1));
  and2  gate2845(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2846(.a(s_328), .O(gate506inter3));
  inv1  gate2847(.a(s_329), .O(gate506inter4));
  nand2 gate2848(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2849(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2850(.a(G1274), .O(gate506inter7));
  inv1  gate2851(.a(G1275), .O(gate506inter8));
  nand2 gate2852(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2853(.a(s_329), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2854(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2855(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2856(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1135(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1136(.a(gate509inter0), .b(s_84), .O(gate509inter1));
  and2  gate1137(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1138(.a(s_84), .O(gate509inter3));
  inv1  gate1139(.a(s_85), .O(gate509inter4));
  nand2 gate1140(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1141(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1142(.a(G1280), .O(gate509inter7));
  inv1  gate1143(.a(G1281), .O(gate509inter8));
  nand2 gate1144(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1145(.a(s_85), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1146(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1147(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1148(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1961(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1962(.a(gate510inter0), .b(s_202), .O(gate510inter1));
  and2  gate1963(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1964(.a(s_202), .O(gate510inter3));
  inv1  gate1965(.a(s_203), .O(gate510inter4));
  nand2 gate1966(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1967(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1968(.a(G1282), .O(gate510inter7));
  inv1  gate1969(.a(G1283), .O(gate510inter8));
  nand2 gate1970(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1971(.a(s_203), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1972(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1973(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1974(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1247(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1248(.a(gate512inter0), .b(s_100), .O(gate512inter1));
  and2  gate1249(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1250(.a(s_100), .O(gate512inter3));
  inv1  gate1251(.a(s_101), .O(gate512inter4));
  nand2 gate1252(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1253(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1254(.a(G1286), .O(gate512inter7));
  inv1  gate1255(.a(G1287), .O(gate512inter8));
  nand2 gate1256(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1257(.a(s_101), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1258(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1259(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1260(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate715(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate716(.a(gate513inter0), .b(s_24), .O(gate513inter1));
  and2  gate717(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate718(.a(s_24), .O(gate513inter3));
  inv1  gate719(.a(s_25), .O(gate513inter4));
  nand2 gate720(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate721(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate722(.a(G1288), .O(gate513inter7));
  inv1  gate723(.a(G1289), .O(gate513inter8));
  nand2 gate724(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate725(.a(s_25), .b(gate513inter3), .O(gate513inter10));
  nor2  gate726(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate727(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate728(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1877(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1878(.a(gate514inter0), .b(s_190), .O(gate514inter1));
  and2  gate1879(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1880(.a(s_190), .O(gate514inter3));
  inv1  gate1881(.a(s_191), .O(gate514inter4));
  nand2 gate1882(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1883(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1884(.a(G1290), .O(gate514inter7));
  inv1  gate1885(.a(G1291), .O(gate514inter8));
  nand2 gate1886(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1887(.a(s_191), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1888(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1889(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1890(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule