module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1387(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1388(.a(gate12inter0), .b(s_120), .O(gate12inter1));
  and2  gate1389(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1390(.a(s_120), .O(gate12inter3));
  inv1  gate1391(.a(s_121), .O(gate12inter4));
  nand2 gate1392(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1393(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1394(.a(G7), .O(gate12inter7));
  inv1  gate1395(.a(G8), .O(gate12inter8));
  nand2 gate1396(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1397(.a(s_121), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1398(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1399(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1400(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1205(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1206(.a(gate13inter0), .b(s_94), .O(gate13inter1));
  and2  gate1207(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1208(.a(s_94), .O(gate13inter3));
  inv1  gate1209(.a(s_95), .O(gate13inter4));
  nand2 gate1210(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1211(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1212(.a(G9), .O(gate13inter7));
  inv1  gate1213(.a(G10), .O(gate13inter8));
  nand2 gate1214(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1215(.a(s_95), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1216(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1217(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1218(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1107(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1108(.a(gate14inter0), .b(s_80), .O(gate14inter1));
  and2  gate1109(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1110(.a(s_80), .O(gate14inter3));
  inv1  gate1111(.a(s_81), .O(gate14inter4));
  nand2 gate1112(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1113(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1114(.a(G11), .O(gate14inter7));
  inv1  gate1115(.a(G12), .O(gate14inter8));
  nand2 gate1116(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1117(.a(s_81), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1118(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1119(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1120(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate855(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate856(.a(gate23inter0), .b(s_44), .O(gate23inter1));
  and2  gate857(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate858(.a(s_44), .O(gate23inter3));
  inv1  gate859(.a(s_45), .O(gate23inter4));
  nand2 gate860(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate861(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate862(.a(G29), .O(gate23inter7));
  inv1  gate863(.a(G30), .O(gate23inter8));
  nand2 gate864(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate865(.a(s_45), .b(gate23inter3), .O(gate23inter10));
  nor2  gate866(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate867(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate868(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1345(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1346(.a(gate30inter0), .b(s_114), .O(gate30inter1));
  and2  gate1347(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1348(.a(s_114), .O(gate30inter3));
  inv1  gate1349(.a(s_115), .O(gate30inter4));
  nand2 gate1350(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1351(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1352(.a(G11), .O(gate30inter7));
  inv1  gate1353(.a(G15), .O(gate30inter8));
  nand2 gate1354(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1355(.a(s_115), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1356(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1357(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1358(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate1513(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1514(.a(gate31inter0), .b(s_138), .O(gate31inter1));
  and2  gate1515(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1516(.a(s_138), .O(gate31inter3));
  inv1  gate1517(.a(s_139), .O(gate31inter4));
  nand2 gate1518(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1519(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1520(.a(G4), .O(gate31inter7));
  inv1  gate1521(.a(G8), .O(gate31inter8));
  nand2 gate1522(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1523(.a(s_139), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1524(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1525(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1526(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1429(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1430(.a(gate45inter0), .b(s_126), .O(gate45inter1));
  and2  gate1431(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1432(.a(s_126), .O(gate45inter3));
  inv1  gate1433(.a(s_127), .O(gate45inter4));
  nand2 gate1434(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1435(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1436(.a(G5), .O(gate45inter7));
  inv1  gate1437(.a(G272), .O(gate45inter8));
  nand2 gate1438(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1439(.a(s_127), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1440(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1441(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1442(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1471(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1472(.a(gate46inter0), .b(s_132), .O(gate46inter1));
  and2  gate1473(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1474(.a(s_132), .O(gate46inter3));
  inv1  gate1475(.a(s_133), .O(gate46inter4));
  nand2 gate1476(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1477(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1478(.a(G6), .O(gate46inter7));
  inv1  gate1479(.a(G272), .O(gate46inter8));
  nand2 gate1480(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1481(.a(s_133), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1482(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1483(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1484(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1401(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1402(.a(gate49inter0), .b(s_122), .O(gate49inter1));
  and2  gate1403(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1404(.a(s_122), .O(gate49inter3));
  inv1  gate1405(.a(s_123), .O(gate49inter4));
  nand2 gate1406(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1407(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1408(.a(G9), .O(gate49inter7));
  inv1  gate1409(.a(G278), .O(gate49inter8));
  nand2 gate1410(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1411(.a(s_123), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1412(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1413(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1414(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate729(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate730(.a(gate51inter0), .b(s_26), .O(gate51inter1));
  and2  gate731(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate732(.a(s_26), .O(gate51inter3));
  inv1  gate733(.a(s_27), .O(gate51inter4));
  nand2 gate734(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate735(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate736(.a(G11), .O(gate51inter7));
  inv1  gate737(.a(G281), .O(gate51inter8));
  nand2 gate738(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate739(.a(s_27), .b(gate51inter3), .O(gate51inter10));
  nor2  gate740(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate741(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate742(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate701(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate702(.a(gate55inter0), .b(s_22), .O(gate55inter1));
  and2  gate703(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate704(.a(s_22), .O(gate55inter3));
  inv1  gate705(.a(s_23), .O(gate55inter4));
  nand2 gate706(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate707(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate708(.a(G15), .O(gate55inter7));
  inv1  gate709(.a(G287), .O(gate55inter8));
  nand2 gate710(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate711(.a(s_23), .b(gate55inter3), .O(gate55inter10));
  nor2  gate712(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate713(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate714(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1331(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1332(.a(gate56inter0), .b(s_112), .O(gate56inter1));
  and2  gate1333(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1334(.a(s_112), .O(gate56inter3));
  inv1  gate1335(.a(s_113), .O(gate56inter4));
  nand2 gate1336(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1337(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1338(.a(G16), .O(gate56inter7));
  inv1  gate1339(.a(G287), .O(gate56inter8));
  nand2 gate1340(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1341(.a(s_113), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1342(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1343(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1344(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1569(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1570(.a(gate60inter0), .b(s_146), .O(gate60inter1));
  and2  gate1571(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1572(.a(s_146), .O(gate60inter3));
  inv1  gate1573(.a(s_147), .O(gate60inter4));
  nand2 gate1574(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1575(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1576(.a(G20), .O(gate60inter7));
  inv1  gate1577(.a(G293), .O(gate60inter8));
  nand2 gate1578(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1579(.a(s_147), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1580(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1581(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1582(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate589(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate590(.a(gate63inter0), .b(s_6), .O(gate63inter1));
  and2  gate591(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate592(.a(s_6), .O(gate63inter3));
  inv1  gate593(.a(s_7), .O(gate63inter4));
  nand2 gate594(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate595(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate596(.a(G23), .O(gate63inter7));
  inv1  gate597(.a(G299), .O(gate63inter8));
  nand2 gate598(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate599(.a(s_7), .b(gate63inter3), .O(gate63inter10));
  nor2  gate600(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate601(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate602(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1135(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1136(.a(gate64inter0), .b(s_84), .O(gate64inter1));
  and2  gate1137(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1138(.a(s_84), .O(gate64inter3));
  inv1  gate1139(.a(s_85), .O(gate64inter4));
  nand2 gate1140(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1141(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1142(.a(G24), .O(gate64inter7));
  inv1  gate1143(.a(G299), .O(gate64inter8));
  nand2 gate1144(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1145(.a(s_85), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1146(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1147(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1148(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate743(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate744(.a(gate67inter0), .b(s_28), .O(gate67inter1));
  and2  gate745(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate746(.a(s_28), .O(gate67inter3));
  inv1  gate747(.a(s_29), .O(gate67inter4));
  nand2 gate748(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate749(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate750(.a(G27), .O(gate67inter7));
  inv1  gate751(.a(G305), .O(gate67inter8));
  nand2 gate752(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate753(.a(s_29), .b(gate67inter3), .O(gate67inter10));
  nor2  gate754(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate755(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate756(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1079(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1080(.a(gate70inter0), .b(s_76), .O(gate70inter1));
  and2  gate1081(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1082(.a(s_76), .O(gate70inter3));
  inv1  gate1083(.a(s_77), .O(gate70inter4));
  nand2 gate1084(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1085(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1086(.a(G30), .O(gate70inter7));
  inv1  gate1087(.a(G308), .O(gate70inter8));
  nand2 gate1088(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1089(.a(s_77), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1090(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1091(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1092(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1247(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1248(.a(gate73inter0), .b(s_100), .O(gate73inter1));
  and2  gate1249(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1250(.a(s_100), .O(gate73inter3));
  inv1  gate1251(.a(s_101), .O(gate73inter4));
  nand2 gate1252(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1253(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1254(.a(G1), .O(gate73inter7));
  inv1  gate1255(.a(G314), .O(gate73inter8));
  nand2 gate1256(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1257(.a(s_101), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1258(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1259(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1260(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1457(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1458(.a(gate86inter0), .b(s_130), .O(gate86inter1));
  and2  gate1459(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1460(.a(s_130), .O(gate86inter3));
  inv1  gate1461(.a(s_131), .O(gate86inter4));
  nand2 gate1462(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1463(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1464(.a(G8), .O(gate86inter7));
  inv1  gate1465(.a(G332), .O(gate86inter8));
  nand2 gate1466(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1467(.a(s_131), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1468(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1469(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1470(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1359(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1360(.a(gate87inter0), .b(s_116), .O(gate87inter1));
  and2  gate1361(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1362(.a(s_116), .O(gate87inter3));
  inv1  gate1363(.a(s_117), .O(gate87inter4));
  nand2 gate1364(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1365(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1366(.a(G12), .O(gate87inter7));
  inv1  gate1367(.a(G335), .O(gate87inter8));
  nand2 gate1368(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1369(.a(s_117), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1370(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1371(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1372(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate617(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate618(.a(gate88inter0), .b(s_10), .O(gate88inter1));
  and2  gate619(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate620(.a(s_10), .O(gate88inter3));
  inv1  gate621(.a(s_11), .O(gate88inter4));
  nand2 gate622(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate623(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate624(.a(G16), .O(gate88inter7));
  inv1  gate625(.a(G335), .O(gate88inter8));
  nand2 gate626(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate627(.a(s_11), .b(gate88inter3), .O(gate88inter10));
  nor2  gate628(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate629(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate630(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1555(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1556(.a(gate96inter0), .b(s_144), .O(gate96inter1));
  and2  gate1557(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1558(.a(s_144), .O(gate96inter3));
  inv1  gate1559(.a(s_145), .O(gate96inter4));
  nand2 gate1560(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1561(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1562(.a(G30), .O(gate96inter7));
  inv1  gate1563(.a(G347), .O(gate96inter8));
  nand2 gate1564(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1565(.a(s_145), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1566(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1567(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1568(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate967(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate968(.a(gate99inter0), .b(s_60), .O(gate99inter1));
  and2  gate969(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate970(.a(s_60), .O(gate99inter3));
  inv1  gate971(.a(s_61), .O(gate99inter4));
  nand2 gate972(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate973(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate974(.a(G27), .O(gate99inter7));
  inv1  gate975(.a(G353), .O(gate99inter8));
  nand2 gate976(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate977(.a(s_61), .b(gate99inter3), .O(gate99inter10));
  nor2  gate978(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate979(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate980(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate785(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate786(.a(gate100inter0), .b(s_34), .O(gate100inter1));
  and2  gate787(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate788(.a(s_34), .O(gate100inter3));
  inv1  gate789(.a(s_35), .O(gate100inter4));
  nand2 gate790(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate791(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate792(.a(G31), .O(gate100inter7));
  inv1  gate793(.a(G353), .O(gate100inter8));
  nand2 gate794(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate795(.a(s_35), .b(gate100inter3), .O(gate100inter10));
  nor2  gate796(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate797(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate798(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate883(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate884(.a(gate110inter0), .b(s_48), .O(gate110inter1));
  and2  gate885(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate886(.a(s_48), .O(gate110inter3));
  inv1  gate887(.a(s_49), .O(gate110inter4));
  nand2 gate888(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate889(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate890(.a(G372), .O(gate110inter7));
  inv1  gate891(.a(G373), .O(gate110inter8));
  nand2 gate892(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate893(.a(s_49), .b(gate110inter3), .O(gate110inter10));
  nor2  gate894(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate895(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate896(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate547(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate548(.a(gate113inter0), .b(s_0), .O(gate113inter1));
  and2  gate549(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate550(.a(s_0), .O(gate113inter3));
  inv1  gate551(.a(s_1), .O(gate113inter4));
  nand2 gate552(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate553(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate554(.a(G378), .O(gate113inter7));
  inv1  gate555(.a(G379), .O(gate113inter8));
  nand2 gate556(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate557(.a(s_1), .b(gate113inter3), .O(gate113inter10));
  nor2  gate558(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate559(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate560(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate715(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate716(.a(gate121inter0), .b(s_24), .O(gate121inter1));
  and2  gate717(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate718(.a(s_24), .O(gate121inter3));
  inv1  gate719(.a(s_25), .O(gate121inter4));
  nand2 gate720(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate721(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate722(.a(G394), .O(gate121inter7));
  inv1  gate723(.a(G395), .O(gate121inter8));
  nand2 gate724(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate725(.a(s_25), .b(gate121inter3), .O(gate121inter10));
  nor2  gate726(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate727(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate728(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1415(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1416(.a(gate137inter0), .b(s_124), .O(gate137inter1));
  and2  gate1417(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1418(.a(s_124), .O(gate137inter3));
  inv1  gate1419(.a(s_125), .O(gate137inter4));
  nand2 gate1420(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1421(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1422(.a(G426), .O(gate137inter7));
  inv1  gate1423(.a(G429), .O(gate137inter8));
  nand2 gate1424(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1425(.a(s_125), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1426(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1427(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1428(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate953(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate954(.a(gate141inter0), .b(s_58), .O(gate141inter1));
  and2  gate955(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate956(.a(s_58), .O(gate141inter3));
  inv1  gate957(.a(s_59), .O(gate141inter4));
  nand2 gate958(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate959(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate960(.a(G450), .O(gate141inter7));
  inv1  gate961(.a(G453), .O(gate141inter8));
  nand2 gate962(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate963(.a(s_59), .b(gate141inter3), .O(gate141inter10));
  nor2  gate964(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate965(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate966(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1191(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1192(.a(gate148inter0), .b(s_92), .O(gate148inter1));
  and2  gate1193(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1194(.a(s_92), .O(gate148inter3));
  inv1  gate1195(.a(s_93), .O(gate148inter4));
  nand2 gate1196(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1197(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1198(.a(G492), .O(gate148inter7));
  inv1  gate1199(.a(G495), .O(gate148inter8));
  nand2 gate1200(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1201(.a(s_93), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1202(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1203(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1204(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate659(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate660(.a(gate149inter0), .b(s_16), .O(gate149inter1));
  and2  gate661(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate662(.a(s_16), .O(gate149inter3));
  inv1  gate663(.a(s_17), .O(gate149inter4));
  nand2 gate664(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate665(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate666(.a(G498), .O(gate149inter7));
  inv1  gate667(.a(G501), .O(gate149inter8));
  nand2 gate668(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate669(.a(s_17), .b(gate149inter3), .O(gate149inter10));
  nor2  gate670(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate671(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate672(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate673(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate674(.a(gate161inter0), .b(s_18), .O(gate161inter1));
  and2  gate675(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate676(.a(s_18), .O(gate161inter3));
  inv1  gate677(.a(s_19), .O(gate161inter4));
  nand2 gate678(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate679(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate680(.a(G450), .O(gate161inter7));
  inv1  gate681(.a(G534), .O(gate161inter8));
  nand2 gate682(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate683(.a(s_19), .b(gate161inter3), .O(gate161inter10));
  nor2  gate684(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate685(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate686(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1373(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1374(.a(gate167inter0), .b(s_118), .O(gate167inter1));
  and2  gate1375(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1376(.a(s_118), .O(gate167inter3));
  inv1  gate1377(.a(s_119), .O(gate167inter4));
  nand2 gate1378(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1379(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1380(.a(G468), .O(gate167inter7));
  inv1  gate1381(.a(G543), .O(gate167inter8));
  nand2 gate1382(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1383(.a(s_119), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1384(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1385(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1386(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate813(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate814(.a(gate168inter0), .b(s_38), .O(gate168inter1));
  and2  gate815(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate816(.a(s_38), .O(gate168inter3));
  inv1  gate817(.a(s_39), .O(gate168inter4));
  nand2 gate818(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate819(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate820(.a(G471), .O(gate168inter7));
  inv1  gate821(.a(G543), .O(gate168inter8));
  nand2 gate822(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate823(.a(s_39), .b(gate168inter3), .O(gate168inter10));
  nor2  gate824(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate825(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate826(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1499(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1500(.a(gate169inter0), .b(s_136), .O(gate169inter1));
  and2  gate1501(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1502(.a(s_136), .O(gate169inter3));
  inv1  gate1503(.a(s_137), .O(gate169inter4));
  nand2 gate1504(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1505(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1506(.a(G474), .O(gate169inter7));
  inv1  gate1507(.a(G546), .O(gate169inter8));
  nand2 gate1508(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1509(.a(s_137), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1510(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1511(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1512(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate799(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate800(.a(gate173inter0), .b(s_36), .O(gate173inter1));
  and2  gate801(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate802(.a(s_36), .O(gate173inter3));
  inv1  gate803(.a(s_37), .O(gate173inter4));
  nand2 gate804(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate805(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate806(.a(G486), .O(gate173inter7));
  inv1  gate807(.a(G552), .O(gate173inter8));
  nand2 gate808(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate809(.a(s_37), .b(gate173inter3), .O(gate173inter10));
  nor2  gate810(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate811(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate812(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate981(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate982(.a(gate179inter0), .b(s_62), .O(gate179inter1));
  and2  gate983(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate984(.a(s_62), .O(gate179inter3));
  inv1  gate985(.a(s_63), .O(gate179inter4));
  nand2 gate986(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate987(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate988(.a(G504), .O(gate179inter7));
  inv1  gate989(.a(G561), .O(gate179inter8));
  nand2 gate990(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate991(.a(s_63), .b(gate179inter3), .O(gate179inter10));
  nor2  gate992(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate993(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate994(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1597(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1598(.a(gate189inter0), .b(s_150), .O(gate189inter1));
  and2  gate1599(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1600(.a(s_150), .O(gate189inter3));
  inv1  gate1601(.a(s_151), .O(gate189inter4));
  nand2 gate1602(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1603(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1604(.a(G578), .O(gate189inter7));
  inv1  gate1605(.a(G579), .O(gate189inter8));
  nand2 gate1606(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1607(.a(s_151), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1608(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1609(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1610(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate827(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate828(.a(gate196inter0), .b(s_40), .O(gate196inter1));
  and2  gate829(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate830(.a(s_40), .O(gate196inter3));
  inv1  gate831(.a(s_41), .O(gate196inter4));
  nand2 gate832(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate833(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate834(.a(G592), .O(gate196inter7));
  inv1  gate835(.a(G593), .O(gate196inter8));
  nand2 gate836(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate837(.a(s_41), .b(gate196inter3), .O(gate196inter10));
  nor2  gate838(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate839(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate840(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1485(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1486(.a(gate198inter0), .b(s_134), .O(gate198inter1));
  and2  gate1487(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1488(.a(s_134), .O(gate198inter3));
  inv1  gate1489(.a(s_135), .O(gate198inter4));
  nand2 gate1490(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1491(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1492(.a(G596), .O(gate198inter7));
  inv1  gate1493(.a(G597), .O(gate198inter8));
  nand2 gate1494(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1495(.a(s_135), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1496(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1497(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1498(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1163(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1164(.a(gate201inter0), .b(s_88), .O(gate201inter1));
  and2  gate1165(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1166(.a(s_88), .O(gate201inter3));
  inv1  gate1167(.a(s_89), .O(gate201inter4));
  nand2 gate1168(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1169(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1170(.a(G602), .O(gate201inter7));
  inv1  gate1171(.a(G607), .O(gate201inter8));
  nand2 gate1172(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1173(.a(s_89), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1174(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1175(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1176(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate575(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate576(.a(gate210inter0), .b(s_4), .O(gate210inter1));
  and2  gate577(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate578(.a(s_4), .O(gate210inter3));
  inv1  gate579(.a(s_5), .O(gate210inter4));
  nand2 gate580(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate581(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate582(.a(G607), .O(gate210inter7));
  inv1  gate583(.a(G666), .O(gate210inter8));
  nand2 gate584(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate585(.a(s_5), .b(gate210inter3), .O(gate210inter10));
  nor2  gate586(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate587(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate588(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate771(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate772(.a(gate211inter0), .b(s_32), .O(gate211inter1));
  and2  gate773(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate774(.a(s_32), .O(gate211inter3));
  inv1  gate775(.a(s_33), .O(gate211inter4));
  nand2 gate776(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate777(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate778(.a(G612), .O(gate211inter7));
  inv1  gate779(.a(G669), .O(gate211inter8));
  nand2 gate780(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate781(.a(s_33), .b(gate211inter3), .O(gate211inter10));
  nor2  gate782(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate783(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate784(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate925(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate926(.a(gate225inter0), .b(s_54), .O(gate225inter1));
  and2  gate927(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate928(.a(s_54), .O(gate225inter3));
  inv1  gate929(.a(s_55), .O(gate225inter4));
  nand2 gate930(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate931(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate932(.a(G690), .O(gate225inter7));
  inv1  gate933(.a(G691), .O(gate225inter8));
  nand2 gate934(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate935(.a(s_55), .b(gate225inter3), .O(gate225inter10));
  nor2  gate936(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate937(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate938(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1009(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1010(.a(gate234inter0), .b(s_66), .O(gate234inter1));
  and2  gate1011(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1012(.a(s_66), .O(gate234inter3));
  inv1  gate1013(.a(s_67), .O(gate234inter4));
  nand2 gate1014(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1015(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1016(.a(G245), .O(gate234inter7));
  inv1  gate1017(.a(G721), .O(gate234inter8));
  nand2 gate1018(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1019(.a(s_67), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1020(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1021(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1022(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1219(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1220(.a(gate241inter0), .b(s_96), .O(gate241inter1));
  and2  gate1221(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1222(.a(s_96), .O(gate241inter3));
  inv1  gate1223(.a(s_97), .O(gate241inter4));
  nand2 gate1224(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1225(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1226(.a(G242), .O(gate241inter7));
  inv1  gate1227(.a(G730), .O(gate241inter8));
  nand2 gate1228(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1229(.a(s_97), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1230(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1231(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1232(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1583(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1584(.a(gate247inter0), .b(s_148), .O(gate247inter1));
  and2  gate1585(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1586(.a(s_148), .O(gate247inter3));
  inv1  gate1587(.a(s_149), .O(gate247inter4));
  nand2 gate1588(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1589(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1590(.a(G251), .O(gate247inter7));
  inv1  gate1591(.a(G739), .O(gate247inter8));
  nand2 gate1592(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1593(.a(s_149), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1594(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1595(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1596(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1527(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1528(.a(gate261inter0), .b(s_140), .O(gate261inter1));
  and2  gate1529(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1530(.a(s_140), .O(gate261inter3));
  inv1  gate1531(.a(s_141), .O(gate261inter4));
  nand2 gate1532(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1533(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1534(.a(G762), .O(gate261inter7));
  inv1  gate1535(.a(G763), .O(gate261inter8));
  nand2 gate1536(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1537(.a(s_141), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1538(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1539(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1540(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate687(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate688(.a(gate277inter0), .b(s_20), .O(gate277inter1));
  and2  gate689(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate690(.a(s_20), .O(gate277inter3));
  inv1  gate691(.a(s_21), .O(gate277inter4));
  nand2 gate692(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate693(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate694(.a(G648), .O(gate277inter7));
  inv1  gate695(.a(G800), .O(gate277inter8));
  nand2 gate696(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate697(.a(s_21), .b(gate277inter3), .O(gate277inter10));
  nor2  gate698(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate699(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate700(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1541(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1542(.a(gate281inter0), .b(s_142), .O(gate281inter1));
  and2  gate1543(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1544(.a(s_142), .O(gate281inter3));
  inv1  gate1545(.a(s_143), .O(gate281inter4));
  nand2 gate1546(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1547(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1548(.a(G654), .O(gate281inter7));
  inv1  gate1549(.a(G806), .O(gate281inter8));
  nand2 gate1550(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1551(.a(s_143), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1552(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1553(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1554(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate995(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate996(.a(gate284inter0), .b(s_64), .O(gate284inter1));
  and2  gate997(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate998(.a(s_64), .O(gate284inter3));
  inv1  gate999(.a(s_65), .O(gate284inter4));
  nand2 gate1000(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1001(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1002(.a(G785), .O(gate284inter7));
  inv1  gate1003(.a(G809), .O(gate284inter8));
  nand2 gate1004(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1005(.a(s_65), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1006(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1007(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1008(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate757(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate758(.a(gate285inter0), .b(s_30), .O(gate285inter1));
  and2  gate759(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate760(.a(s_30), .O(gate285inter3));
  inv1  gate761(.a(s_31), .O(gate285inter4));
  nand2 gate762(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate763(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate764(.a(G660), .O(gate285inter7));
  inv1  gate765(.a(G812), .O(gate285inter8));
  nand2 gate766(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate767(.a(s_31), .b(gate285inter3), .O(gate285inter10));
  nor2  gate768(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate769(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate770(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1261(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1262(.a(gate289inter0), .b(s_102), .O(gate289inter1));
  and2  gate1263(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1264(.a(s_102), .O(gate289inter3));
  inv1  gate1265(.a(s_103), .O(gate289inter4));
  nand2 gate1266(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1267(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1268(.a(G818), .O(gate289inter7));
  inv1  gate1269(.a(G819), .O(gate289inter8));
  nand2 gate1270(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1271(.a(s_103), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1272(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1273(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1274(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1149(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1150(.a(gate293inter0), .b(s_86), .O(gate293inter1));
  and2  gate1151(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1152(.a(s_86), .O(gate293inter3));
  inv1  gate1153(.a(s_87), .O(gate293inter4));
  nand2 gate1154(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1155(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1156(.a(G828), .O(gate293inter7));
  inv1  gate1157(.a(G829), .O(gate293inter8));
  nand2 gate1158(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1159(.a(s_87), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1160(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1161(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1162(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate603(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate604(.a(gate294inter0), .b(s_8), .O(gate294inter1));
  and2  gate605(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate606(.a(s_8), .O(gate294inter3));
  inv1  gate607(.a(s_9), .O(gate294inter4));
  nand2 gate608(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate609(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate610(.a(G832), .O(gate294inter7));
  inv1  gate611(.a(G833), .O(gate294inter8));
  nand2 gate612(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate613(.a(s_9), .b(gate294inter3), .O(gate294inter10));
  nor2  gate614(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate615(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate616(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate939(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate940(.a(gate392inter0), .b(s_56), .O(gate392inter1));
  and2  gate941(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate942(.a(s_56), .O(gate392inter3));
  inv1  gate943(.a(s_57), .O(gate392inter4));
  nand2 gate944(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate945(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate946(.a(G6), .O(gate392inter7));
  inv1  gate947(.a(G1051), .O(gate392inter8));
  nand2 gate948(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate949(.a(s_57), .b(gate392inter3), .O(gate392inter10));
  nor2  gate950(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate951(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate952(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1303(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1304(.a(gate407inter0), .b(s_108), .O(gate407inter1));
  and2  gate1305(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1306(.a(s_108), .O(gate407inter3));
  inv1  gate1307(.a(s_109), .O(gate407inter4));
  nand2 gate1308(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1309(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1310(.a(G21), .O(gate407inter7));
  inv1  gate1311(.a(G1096), .O(gate407inter8));
  nand2 gate1312(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1313(.a(s_109), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1314(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1315(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1316(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1289(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1290(.a(gate411inter0), .b(s_106), .O(gate411inter1));
  and2  gate1291(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1292(.a(s_106), .O(gate411inter3));
  inv1  gate1293(.a(s_107), .O(gate411inter4));
  nand2 gate1294(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1295(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1296(.a(G25), .O(gate411inter7));
  inv1  gate1297(.a(G1108), .O(gate411inter8));
  nand2 gate1298(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1299(.a(s_107), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1300(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1301(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1302(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate561(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate562(.a(gate415inter0), .b(s_2), .O(gate415inter1));
  and2  gate563(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate564(.a(s_2), .O(gate415inter3));
  inv1  gate565(.a(s_3), .O(gate415inter4));
  nand2 gate566(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate567(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate568(.a(G29), .O(gate415inter7));
  inv1  gate569(.a(G1120), .O(gate415inter8));
  nand2 gate570(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate571(.a(s_3), .b(gate415inter3), .O(gate415inter10));
  nor2  gate572(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate573(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate574(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1121(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1122(.a(gate416inter0), .b(s_82), .O(gate416inter1));
  and2  gate1123(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1124(.a(s_82), .O(gate416inter3));
  inv1  gate1125(.a(s_83), .O(gate416inter4));
  nand2 gate1126(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1127(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1128(.a(G30), .O(gate416inter7));
  inv1  gate1129(.a(G1123), .O(gate416inter8));
  nand2 gate1130(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1131(.a(s_83), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1132(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1133(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1134(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1317(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1318(.a(gate421inter0), .b(s_110), .O(gate421inter1));
  and2  gate1319(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1320(.a(s_110), .O(gate421inter3));
  inv1  gate1321(.a(s_111), .O(gate421inter4));
  nand2 gate1322(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1323(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1324(.a(G2), .O(gate421inter7));
  inv1  gate1325(.a(G1135), .O(gate421inter8));
  nand2 gate1326(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1327(.a(s_111), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1328(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1329(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1330(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate897(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate898(.a(gate423inter0), .b(s_50), .O(gate423inter1));
  and2  gate899(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate900(.a(s_50), .O(gate423inter3));
  inv1  gate901(.a(s_51), .O(gate423inter4));
  nand2 gate902(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate903(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate904(.a(G3), .O(gate423inter7));
  inv1  gate905(.a(G1138), .O(gate423inter8));
  nand2 gate906(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate907(.a(s_51), .b(gate423inter3), .O(gate423inter10));
  nor2  gate908(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate909(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate910(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate841(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate842(.a(gate433inter0), .b(s_42), .O(gate433inter1));
  and2  gate843(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate844(.a(s_42), .O(gate433inter3));
  inv1  gate845(.a(s_43), .O(gate433inter4));
  nand2 gate846(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate847(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate848(.a(G8), .O(gate433inter7));
  inv1  gate849(.a(G1153), .O(gate433inter8));
  nand2 gate850(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate851(.a(s_43), .b(gate433inter3), .O(gate433inter10));
  nor2  gate852(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate853(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate854(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1233(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1234(.a(gate444inter0), .b(s_98), .O(gate444inter1));
  and2  gate1235(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1236(.a(s_98), .O(gate444inter3));
  inv1  gate1237(.a(s_99), .O(gate444inter4));
  nand2 gate1238(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1239(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1240(.a(G1072), .O(gate444inter7));
  inv1  gate1241(.a(G1168), .O(gate444inter8));
  nand2 gate1242(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1243(.a(s_99), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1244(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1245(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1246(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1177(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1178(.a(gate446inter0), .b(s_90), .O(gate446inter1));
  and2  gate1179(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1180(.a(s_90), .O(gate446inter3));
  inv1  gate1181(.a(s_91), .O(gate446inter4));
  nand2 gate1182(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1183(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1184(.a(G1075), .O(gate446inter7));
  inv1  gate1185(.a(G1171), .O(gate446inter8));
  nand2 gate1186(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1187(.a(s_91), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1188(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1189(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1190(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1065(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1066(.a(gate469inter0), .b(s_74), .O(gate469inter1));
  and2  gate1067(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1068(.a(s_74), .O(gate469inter3));
  inv1  gate1069(.a(s_75), .O(gate469inter4));
  nand2 gate1070(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1071(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1072(.a(G26), .O(gate469inter7));
  inv1  gate1073(.a(G1207), .O(gate469inter8));
  nand2 gate1074(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1075(.a(s_75), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1076(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1077(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1078(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1023(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1024(.a(gate472inter0), .b(s_68), .O(gate472inter1));
  and2  gate1025(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1026(.a(s_68), .O(gate472inter3));
  inv1  gate1027(.a(s_69), .O(gate472inter4));
  nand2 gate1028(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1029(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1030(.a(G1114), .O(gate472inter7));
  inv1  gate1031(.a(G1210), .O(gate472inter8));
  nand2 gate1032(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1033(.a(s_69), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1034(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1035(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1036(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1443(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1444(.a(gate473inter0), .b(s_128), .O(gate473inter1));
  and2  gate1445(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1446(.a(s_128), .O(gate473inter3));
  inv1  gate1447(.a(s_129), .O(gate473inter4));
  nand2 gate1448(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1449(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1450(.a(G28), .O(gate473inter7));
  inv1  gate1451(.a(G1213), .O(gate473inter8));
  nand2 gate1452(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1453(.a(s_129), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1454(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1455(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1456(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1093(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1094(.a(gate477inter0), .b(s_78), .O(gate477inter1));
  and2  gate1095(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1096(.a(s_78), .O(gate477inter3));
  inv1  gate1097(.a(s_79), .O(gate477inter4));
  nand2 gate1098(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1099(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1100(.a(G30), .O(gate477inter7));
  inv1  gate1101(.a(G1219), .O(gate477inter8));
  nand2 gate1102(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1103(.a(s_79), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1104(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1105(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1106(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate645(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate646(.a(gate480inter0), .b(s_14), .O(gate480inter1));
  and2  gate647(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate648(.a(s_14), .O(gate480inter3));
  inv1  gate649(.a(s_15), .O(gate480inter4));
  nand2 gate650(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate651(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate652(.a(G1126), .O(gate480inter7));
  inv1  gate653(.a(G1222), .O(gate480inter8));
  nand2 gate654(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate655(.a(s_15), .b(gate480inter3), .O(gate480inter10));
  nor2  gate656(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate657(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate658(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1275(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1276(.a(gate483inter0), .b(s_104), .O(gate483inter1));
  and2  gate1277(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1278(.a(s_104), .O(gate483inter3));
  inv1  gate1279(.a(s_105), .O(gate483inter4));
  nand2 gate1280(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1281(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1282(.a(G1228), .O(gate483inter7));
  inv1  gate1283(.a(G1229), .O(gate483inter8));
  nand2 gate1284(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1285(.a(s_105), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1286(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1287(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1288(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1051(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1052(.a(gate484inter0), .b(s_72), .O(gate484inter1));
  and2  gate1053(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1054(.a(s_72), .O(gate484inter3));
  inv1  gate1055(.a(s_73), .O(gate484inter4));
  nand2 gate1056(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1057(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1058(.a(G1230), .O(gate484inter7));
  inv1  gate1059(.a(G1231), .O(gate484inter8));
  nand2 gate1060(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1061(.a(s_73), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1062(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1063(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1064(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate869(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate870(.a(gate497inter0), .b(s_46), .O(gate497inter1));
  and2  gate871(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate872(.a(s_46), .O(gate497inter3));
  inv1  gate873(.a(s_47), .O(gate497inter4));
  nand2 gate874(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate875(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate876(.a(G1256), .O(gate497inter7));
  inv1  gate877(.a(G1257), .O(gate497inter8));
  nand2 gate878(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate879(.a(s_47), .b(gate497inter3), .O(gate497inter10));
  nor2  gate880(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate881(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate882(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate631(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate632(.a(gate502inter0), .b(s_12), .O(gate502inter1));
  and2  gate633(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate634(.a(s_12), .O(gate502inter3));
  inv1  gate635(.a(s_13), .O(gate502inter4));
  nand2 gate636(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate637(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate638(.a(G1266), .O(gate502inter7));
  inv1  gate639(.a(G1267), .O(gate502inter8));
  nand2 gate640(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate641(.a(s_13), .b(gate502inter3), .O(gate502inter10));
  nor2  gate642(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate643(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate644(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate911(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate912(.a(gate507inter0), .b(s_52), .O(gate507inter1));
  and2  gate913(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate914(.a(s_52), .O(gate507inter3));
  inv1  gate915(.a(s_53), .O(gate507inter4));
  nand2 gate916(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate917(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate918(.a(G1276), .O(gate507inter7));
  inv1  gate919(.a(G1277), .O(gate507inter8));
  nand2 gate920(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate921(.a(s_53), .b(gate507inter3), .O(gate507inter10));
  nor2  gate922(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate923(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate924(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1037(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1038(.a(gate510inter0), .b(s_70), .O(gate510inter1));
  and2  gate1039(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1040(.a(s_70), .O(gate510inter3));
  inv1  gate1041(.a(s_71), .O(gate510inter4));
  nand2 gate1042(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1043(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1044(.a(G1282), .O(gate510inter7));
  inv1  gate1045(.a(G1283), .O(gate510inter8));
  nand2 gate1046(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1047(.a(s_71), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1048(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1049(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1050(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule