module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1275(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1276(.a(gate11inter0), .b(s_104), .O(gate11inter1));
  and2  gate1277(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1278(.a(s_104), .O(gate11inter3));
  inv1  gate1279(.a(s_105), .O(gate11inter4));
  nand2 gate1280(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1281(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1282(.a(G5), .O(gate11inter7));
  inv1  gate1283(.a(G6), .O(gate11inter8));
  nand2 gate1284(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1285(.a(s_105), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1286(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1287(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1288(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate925(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate926(.a(gate12inter0), .b(s_54), .O(gate12inter1));
  and2  gate927(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate928(.a(s_54), .O(gate12inter3));
  inv1  gate929(.a(s_55), .O(gate12inter4));
  nand2 gate930(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate931(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate932(.a(G7), .O(gate12inter7));
  inv1  gate933(.a(G8), .O(gate12inter8));
  nand2 gate934(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate935(.a(s_55), .b(gate12inter3), .O(gate12inter10));
  nor2  gate936(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate937(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate938(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1989(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1990(.a(gate13inter0), .b(s_206), .O(gate13inter1));
  and2  gate1991(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1992(.a(s_206), .O(gate13inter3));
  inv1  gate1993(.a(s_207), .O(gate13inter4));
  nand2 gate1994(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1995(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1996(.a(G9), .O(gate13inter7));
  inv1  gate1997(.a(G10), .O(gate13inter8));
  nand2 gate1998(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1999(.a(s_207), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2000(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2001(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2002(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate547(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate548(.a(gate14inter0), .b(s_0), .O(gate14inter1));
  and2  gate549(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate550(.a(s_0), .O(gate14inter3));
  inv1  gate551(.a(s_1), .O(gate14inter4));
  nand2 gate552(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate553(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate554(.a(G11), .O(gate14inter7));
  inv1  gate555(.a(G12), .O(gate14inter8));
  nand2 gate556(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate557(.a(s_1), .b(gate14inter3), .O(gate14inter10));
  nor2  gate558(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate559(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate560(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1345(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1346(.a(gate18inter0), .b(s_114), .O(gate18inter1));
  and2  gate1347(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1348(.a(s_114), .O(gate18inter3));
  inv1  gate1349(.a(s_115), .O(gate18inter4));
  nand2 gate1350(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1351(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1352(.a(G19), .O(gate18inter7));
  inv1  gate1353(.a(G20), .O(gate18inter8));
  nand2 gate1354(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1355(.a(s_115), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1356(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1357(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1358(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1975(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1976(.a(gate29inter0), .b(s_204), .O(gate29inter1));
  and2  gate1977(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1978(.a(s_204), .O(gate29inter3));
  inv1  gate1979(.a(s_205), .O(gate29inter4));
  nand2 gate1980(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1981(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1982(.a(G3), .O(gate29inter7));
  inv1  gate1983(.a(G7), .O(gate29inter8));
  nand2 gate1984(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1985(.a(s_205), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1986(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1987(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1988(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1597(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1598(.a(gate32inter0), .b(s_150), .O(gate32inter1));
  and2  gate1599(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1600(.a(s_150), .O(gate32inter3));
  inv1  gate1601(.a(s_151), .O(gate32inter4));
  nand2 gate1602(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1603(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1604(.a(G12), .O(gate32inter7));
  inv1  gate1605(.a(G16), .O(gate32inter8));
  nand2 gate1606(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1607(.a(s_151), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1608(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1609(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1610(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1639(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1640(.a(gate33inter0), .b(s_156), .O(gate33inter1));
  and2  gate1641(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1642(.a(s_156), .O(gate33inter3));
  inv1  gate1643(.a(s_157), .O(gate33inter4));
  nand2 gate1644(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1645(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1646(.a(G17), .O(gate33inter7));
  inv1  gate1647(.a(G21), .O(gate33inter8));
  nand2 gate1648(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1649(.a(s_157), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1650(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1651(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1652(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1303(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1304(.a(gate34inter0), .b(s_108), .O(gate34inter1));
  and2  gate1305(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1306(.a(s_108), .O(gate34inter3));
  inv1  gate1307(.a(s_109), .O(gate34inter4));
  nand2 gate1308(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1309(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1310(.a(G25), .O(gate34inter7));
  inv1  gate1311(.a(G29), .O(gate34inter8));
  nand2 gate1312(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1313(.a(s_109), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1314(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1315(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1316(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1807(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1808(.a(gate43inter0), .b(s_180), .O(gate43inter1));
  and2  gate1809(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1810(.a(s_180), .O(gate43inter3));
  inv1  gate1811(.a(s_181), .O(gate43inter4));
  nand2 gate1812(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1813(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1814(.a(G3), .O(gate43inter7));
  inv1  gate1815(.a(G269), .O(gate43inter8));
  nand2 gate1816(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1817(.a(s_181), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1818(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1819(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1820(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1009(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1010(.a(gate44inter0), .b(s_66), .O(gate44inter1));
  and2  gate1011(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1012(.a(s_66), .O(gate44inter3));
  inv1  gate1013(.a(s_67), .O(gate44inter4));
  nand2 gate1014(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1015(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1016(.a(G4), .O(gate44inter7));
  inv1  gate1017(.a(G269), .O(gate44inter8));
  nand2 gate1018(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1019(.a(s_67), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1020(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1021(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1022(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1121(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1122(.a(gate45inter0), .b(s_82), .O(gate45inter1));
  and2  gate1123(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1124(.a(s_82), .O(gate45inter3));
  inv1  gate1125(.a(s_83), .O(gate45inter4));
  nand2 gate1126(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1127(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1128(.a(G5), .O(gate45inter7));
  inv1  gate1129(.a(G272), .O(gate45inter8));
  nand2 gate1130(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1131(.a(s_83), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1132(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1133(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1134(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate939(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate940(.a(gate47inter0), .b(s_56), .O(gate47inter1));
  and2  gate941(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate942(.a(s_56), .O(gate47inter3));
  inv1  gate943(.a(s_57), .O(gate47inter4));
  nand2 gate944(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate945(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate946(.a(G7), .O(gate47inter7));
  inv1  gate947(.a(G275), .O(gate47inter8));
  nand2 gate948(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate949(.a(s_57), .b(gate47inter3), .O(gate47inter10));
  nor2  gate950(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate951(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate952(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate995(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate996(.a(gate50inter0), .b(s_64), .O(gate50inter1));
  and2  gate997(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate998(.a(s_64), .O(gate50inter3));
  inv1  gate999(.a(s_65), .O(gate50inter4));
  nand2 gate1000(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1001(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1002(.a(G10), .O(gate50inter7));
  inv1  gate1003(.a(G278), .O(gate50inter8));
  nand2 gate1004(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1005(.a(s_65), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1006(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1007(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1008(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate785(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate786(.a(gate59inter0), .b(s_34), .O(gate59inter1));
  and2  gate787(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate788(.a(s_34), .O(gate59inter3));
  inv1  gate789(.a(s_35), .O(gate59inter4));
  nand2 gate790(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate791(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate792(.a(G19), .O(gate59inter7));
  inv1  gate793(.a(G293), .O(gate59inter8));
  nand2 gate794(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate795(.a(s_35), .b(gate59inter3), .O(gate59inter10));
  nor2  gate796(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate797(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate798(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate1485(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1486(.a(gate60inter0), .b(s_134), .O(gate60inter1));
  and2  gate1487(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1488(.a(s_134), .O(gate60inter3));
  inv1  gate1489(.a(s_135), .O(gate60inter4));
  nand2 gate1490(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1491(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1492(.a(G20), .O(gate60inter7));
  inv1  gate1493(.a(G293), .O(gate60inter8));
  nand2 gate1494(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1495(.a(s_135), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1496(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1497(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1498(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate687(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate688(.a(gate66inter0), .b(s_20), .O(gate66inter1));
  and2  gate689(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate690(.a(s_20), .O(gate66inter3));
  inv1  gate691(.a(s_21), .O(gate66inter4));
  nand2 gate692(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate693(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate694(.a(G26), .O(gate66inter7));
  inv1  gate695(.a(G302), .O(gate66inter8));
  nand2 gate696(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate697(.a(s_21), .b(gate66inter3), .O(gate66inter10));
  nor2  gate698(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate699(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate700(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1149(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1150(.a(gate77inter0), .b(s_86), .O(gate77inter1));
  and2  gate1151(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1152(.a(s_86), .O(gate77inter3));
  inv1  gate1153(.a(s_87), .O(gate77inter4));
  nand2 gate1154(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1155(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1156(.a(G2), .O(gate77inter7));
  inv1  gate1157(.a(G320), .O(gate77inter8));
  nand2 gate1158(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1159(.a(s_87), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1160(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1161(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1162(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2087(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2088(.a(gate80inter0), .b(s_220), .O(gate80inter1));
  and2  gate2089(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2090(.a(s_220), .O(gate80inter3));
  inv1  gate2091(.a(s_221), .O(gate80inter4));
  nand2 gate2092(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2093(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2094(.a(G14), .O(gate80inter7));
  inv1  gate2095(.a(G323), .O(gate80inter8));
  nand2 gate2096(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2097(.a(s_221), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2098(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2099(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2100(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1387(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1388(.a(gate82inter0), .b(s_120), .O(gate82inter1));
  and2  gate1389(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1390(.a(s_120), .O(gate82inter3));
  inv1  gate1391(.a(s_121), .O(gate82inter4));
  nand2 gate1392(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1393(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1394(.a(G7), .O(gate82inter7));
  inv1  gate1395(.a(G326), .O(gate82inter8));
  nand2 gate1396(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1397(.a(s_121), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1398(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1399(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1400(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1331(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1332(.a(gate84inter0), .b(s_112), .O(gate84inter1));
  and2  gate1333(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1334(.a(s_112), .O(gate84inter3));
  inv1  gate1335(.a(s_113), .O(gate84inter4));
  nand2 gate1336(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1337(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1338(.a(G15), .O(gate84inter7));
  inv1  gate1339(.a(G329), .O(gate84inter8));
  nand2 gate1340(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1341(.a(s_113), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1342(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1343(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1344(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1541(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1542(.a(gate88inter0), .b(s_142), .O(gate88inter1));
  and2  gate1543(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1544(.a(s_142), .O(gate88inter3));
  inv1  gate1545(.a(s_143), .O(gate88inter4));
  nand2 gate1546(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1547(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1548(.a(G16), .O(gate88inter7));
  inv1  gate1549(.a(G335), .O(gate88inter8));
  nand2 gate1550(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1551(.a(s_143), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1552(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1553(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1554(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate589(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate590(.a(gate90inter0), .b(s_6), .O(gate90inter1));
  and2  gate591(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate592(.a(s_6), .O(gate90inter3));
  inv1  gate593(.a(s_7), .O(gate90inter4));
  nand2 gate594(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate595(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate596(.a(G21), .O(gate90inter7));
  inv1  gate597(.a(G338), .O(gate90inter8));
  nand2 gate598(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate599(.a(s_7), .b(gate90inter3), .O(gate90inter10));
  nor2  gate600(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate601(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate602(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate1527(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1528(.a(gate91inter0), .b(s_140), .O(gate91inter1));
  and2  gate1529(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1530(.a(s_140), .O(gate91inter3));
  inv1  gate1531(.a(s_141), .O(gate91inter4));
  nand2 gate1532(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1533(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1534(.a(G25), .O(gate91inter7));
  inv1  gate1535(.a(G341), .O(gate91inter8));
  nand2 gate1536(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1537(.a(s_141), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1538(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1539(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1540(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate715(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate716(.a(gate96inter0), .b(s_24), .O(gate96inter1));
  and2  gate717(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate718(.a(s_24), .O(gate96inter3));
  inv1  gate719(.a(s_25), .O(gate96inter4));
  nand2 gate720(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate721(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate722(.a(G30), .O(gate96inter7));
  inv1  gate723(.a(G347), .O(gate96inter8));
  nand2 gate724(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate725(.a(s_25), .b(gate96inter3), .O(gate96inter10));
  nor2  gate726(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate727(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate728(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate911(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate912(.a(gate97inter0), .b(s_52), .O(gate97inter1));
  and2  gate913(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate914(.a(s_52), .O(gate97inter3));
  inv1  gate915(.a(s_53), .O(gate97inter4));
  nand2 gate916(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate917(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate918(.a(G19), .O(gate97inter7));
  inv1  gate919(.a(G350), .O(gate97inter8));
  nand2 gate920(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate921(.a(s_53), .b(gate97inter3), .O(gate97inter10));
  nor2  gate922(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate923(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate924(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1513(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1514(.a(gate106inter0), .b(s_138), .O(gate106inter1));
  and2  gate1515(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1516(.a(s_138), .O(gate106inter3));
  inv1  gate1517(.a(s_139), .O(gate106inter4));
  nand2 gate1518(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1519(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1520(.a(G364), .O(gate106inter7));
  inv1  gate1521(.a(G365), .O(gate106inter8));
  nand2 gate1522(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1523(.a(s_139), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1524(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1525(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1526(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate701(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate702(.a(gate109inter0), .b(s_22), .O(gate109inter1));
  and2  gate703(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate704(.a(s_22), .O(gate109inter3));
  inv1  gate705(.a(s_23), .O(gate109inter4));
  nand2 gate706(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate707(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate708(.a(G370), .O(gate109inter7));
  inv1  gate709(.a(G371), .O(gate109inter8));
  nand2 gate710(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate711(.a(s_23), .b(gate109inter3), .O(gate109inter10));
  nor2  gate712(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate713(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate714(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate2045(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate2046(.a(gate113inter0), .b(s_214), .O(gate113inter1));
  and2  gate2047(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate2048(.a(s_214), .O(gate113inter3));
  inv1  gate2049(.a(s_215), .O(gate113inter4));
  nand2 gate2050(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate2051(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate2052(.a(G378), .O(gate113inter7));
  inv1  gate2053(.a(G379), .O(gate113inter8));
  nand2 gate2054(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate2055(.a(s_215), .b(gate113inter3), .O(gate113inter10));
  nor2  gate2056(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate2057(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate2058(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate897(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate898(.a(gate116inter0), .b(s_50), .O(gate116inter1));
  and2  gate899(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate900(.a(s_50), .O(gate116inter3));
  inv1  gate901(.a(s_51), .O(gate116inter4));
  nand2 gate902(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate903(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate904(.a(G384), .O(gate116inter7));
  inv1  gate905(.a(G385), .O(gate116inter8));
  nand2 gate906(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate907(.a(s_51), .b(gate116inter3), .O(gate116inter10));
  nor2  gate908(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate909(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate910(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1051(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1052(.a(gate118inter0), .b(s_72), .O(gate118inter1));
  and2  gate1053(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1054(.a(s_72), .O(gate118inter3));
  inv1  gate1055(.a(s_73), .O(gate118inter4));
  nand2 gate1056(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1057(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1058(.a(G388), .O(gate118inter7));
  inv1  gate1059(.a(G389), .O(gate118inter8));
  nand2 gate1060(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1061(.a(s_73), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1062(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1063(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1064(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1835(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1836(.a(gate130inter0), .b(s_184), .O(gate130inter1));
  and2  gate1837(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1838(.a(s_184), .O(gate130inter3));
  inv1  gate1839(.a(s_185), .O(gate130inter4));
  nand2 gate1840(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1841(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1842(.a(G412), .O(gate130inter7));
  inv1  gate1843(.a(G413), .O(gate130inter8));
  nand2 gate1844(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1845(.a(s_185), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1846(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1847(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1848(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2003(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2004(.a(gate140inter0), .b(s_208), .O(gate140inter1));
  and2  gate2005(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2006(.a(s_208), .O(gate140inter3));
  inv1  gate2007(.a(s_209), .O(gate140inter4));
  nand2 gate2008(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2009(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2010(.a(G444), .O(gate140inter7));
  inv1  gate2011(.a(G447), .O(gate140inter8));
  nand2 gate2012(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2013(.a(s_209), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2014(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2015(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2016(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1219(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1220(.a(gate144inter0), .b(s_96), .O(gate144inter1));
  and2  gate1221(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1222(.a(s_96), .O(gate144inter3));
  inv1  gate1223(.a(s_97), .O(gate144inter4));
  nand2 gate1224(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1225(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1226(.a(G468), .O(gate144inter7));
  inv1  gate1227(.a(G471), .O(gate144inter8));
  nand2 gate1228(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1229(.a(s_97), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1230(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1231(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1232(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate771(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate772(.a(gate145inter0), .b(s_32), .O(gate145inter1));
  and2  gate773(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate774(.a(s_32), .O(gate145inter3));
  inv1  gate775(.a(s_33), .O(gate145inter4));
  nand2 gate776(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate777(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate778(.a(G474), .O(gate145inter7));
  inv1  gate779(.a(G477), .O(gate145inter8));
  nand2 gate780(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate781(.a(s_33), .b(gate145inter3), .O(gate145inter10));
  nor2  gate782(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate783(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate784(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2031(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2032(.a(gate152inter0), .b(s_212), .O(gate152inter1));
  and2  gate2033(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2034(.a(s_212), .O(gate152inter3));
  inv1  gate2035(.a(s_213), .O(gate152inter4));
  nand2 gate2036(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2037(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2038(.a(G516), .O(gate152inter7));
  inv1  gate2039(.a(G519), .O(gate152inter8));
  nand2 gate2040(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2041(.a(s_213), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2042(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2043(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2044(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1191(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1192(.a(gate155inter0), .b(s_92), .O(gate155inter1));
  and2  gate1193(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1194(.a(s_92), .O(gate155inter3));
  inv1  gate1195(.a(s_93), .O(gate155inter4));
  nand2 gate1196(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1197(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1198(.a(G432), .O(gate155inter7));
  inv1  gate1199(.a(G525), .O(gate155inter8));
  nand2 gate1200(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1201(.a(s_93), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1202(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1203(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1204(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1205(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1206(.a(gate158inter0), .b(s_94), .O(gate158inter1));
  and2  gate1207(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1208(.a(s_94), .O(gate158inter3));
  inv1  gate1209(.a(s_95), .O(gate158inter4));
  nand2 gate1210(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1211(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1212(.a(G441), .O(gate158inter7));
  inv1  gate1213(.a(G528), .O(gate158inter8));
  nand2 gate1214(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1215(.a(s_95), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1216(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1217(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1218(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1667(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1668(.a(gate163inter0), .b(s_160), .O(gate163inter1));
  and2  gate1669(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1670(.a(s_160), .O(gate163inter3));
  inv1  gate1671(.a(s_161), .O(gate163inter4));
  nand2 gate1672(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1673(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1674(.a(G456), .O(gate163inter7));
  inv1  gate1675(.a(G537), .O(gate163inter8));
  nand2 gate1676(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1677(.a(s_161), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1678(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1679(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1680(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate869(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate870(.a(gate164inter0), .b(s_46), .O(gate164inter1));
  and2  gate871(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate872(.a(s_46), .O(gate164inter3));
  inv1  gate873(.a(s_47), .O(gate164inter4));
  nand2 gate874(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate875(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate876(.a(G459), .O(gate164inter7));
  inv1  gate877(.a(G537), .O(gate164inter8));
  nand2 gate878(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate879(.a(s_47), .b(gate164inter3), .O(gate164inter10));
  nor2  gate880(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate881(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate882(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1317(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1318(.a(gate179inter0), .b(s_110), .O(gate179inter1));
  and2  gate1319(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1320(.a(s_110), .O(gate179inter3));
  inv1  gate1321(.a(s_111), .O(gate179inter4));
  nand2 gate1322(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1323(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1324(.a(G504), .O(gate179inter7));
  inv1  gate1325(.a(G561), .O(gate179inter8));
  nand2 gate1326(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1327(.a(s_111), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1328(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1329(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1330(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate2017(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate2018(.a(gate181inter0), .b(s_210), .O(gate181inter1));
  and2  gate2019(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate2020(.a(s_210), .O(gate181inter3));
  inv1  gate2021(.a(s_211), .O(gate181inter4));
  nand2 gate2022(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate2023(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate2024(.a(G510), .O(gate181inter7));
  inv1  gate2025(.a(G564), .O(gate181inter8));
  nand2 gate2026(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate2027(.a(s_211), .b(gate181inter3), .O(gate181inter10));
  nor2  gate2028(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate2029(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate2030(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1261(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1262(.a(gate183inter0), .b(s_102), .O(gate183inter1));
  and2  gate1263(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1264(.a(s_102), .O(gate183inter3));
  inv1  gate1265(.a(s_103), .O(gate183inter4));
  nand2 gate1266(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1267(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1268(.a(G516), .O(gate183inter7));
  inv1  gate1269(.a(G567), .O(gate183inter8));
  nand2 gate1270(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1271(.a(s_103), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1272(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1273(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1274(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1821(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1822(.a(gate184inter0), .b(s_182), .O(gate184inter1));
  and2  gate1823(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1824(.a(s_182), .O(gate184inter3));
  inv1  gate1825(.a(s_183), .O(gate184inter4));
  nand2 gate1826(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1827(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1828(.a(G519), .O(gate184inter7));
  inv1  gate1829(.a(G567), .O(gate184inter8));
  nand2 gate1830(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1831(.a(s_183), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1832(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1833(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1834(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate855(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate856(.a(gate185inter0), .b(s_44), .O(gate185inter1));
  and2  gate857(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate858(.a(s_44), .O(gate185inter3));
  inv1  gate859(.a(s_45), .O(gate185inter4));
  nand2 gate860(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate861(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate862(.a(G570), .O(gate185inter7));
  inv1  gate863(.a(G571), .O(gate185inter8));
  nand2 gate864(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate865(.a(s_45), .b(gate185inter3), .O(gate185inter10));
  nor2  gate866(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate867(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate868(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1933(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1934(.a(gate189inter0), .b(s_198), .O(gate189inter1));
  and2  gate1935(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1936(.a(s_198), .O(gate189inter3));
  inv1  gate1937(.a(s_199), .O(gate189inter4));
  nand2 gate1938(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1939(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1940(.a(G578), .O(gate189inter7));
  inv1  gate1941(.a(G579), .O(gate189inter8));
  nand2 gate1942(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1943(.a(s_199), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1944(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1945(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1946(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1359(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1360(.a(gate190inter0), .b(s_116), .O(gate190inter1));
  and2  gate1361(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1362(.a(s_116), .O(gate190inter3));
  inv1  gate1363(.a(s_117), .O(gate190inter4));
  nand2 gate1364(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1365(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1366(.a(G580), .O(gate190inter7));
  inv1  gate1367(.a(G581), .O(gate190inter8));
  nand2 gate1368(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1369(.a(s_117), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1370(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1371(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1372(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1709(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1710(.a(gate196inter0), .b(s_166), .O(gate196inter1));
  and2  gate1711(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1712(.a(s_166), .O(gate196inter3));
  inv1  gate1713(.a(s_167), .O(gate196inter4));
  nand2 gate1714(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1715(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1716(.a(G592), .O(gate196inter7));
  inv1  gate1717(.a(G593), .O(gate196inter8));
  nand2 gate1718(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1719(.a(s_167), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1720(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1721(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1722(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1079(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1080(.a(gate197inter0), .b(s_76), .O(gate197inter1));
  and2  gate1081(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1082(.a(s_76), .O(gate197inter3));
  inv1  gate1083(.a(s_77), .O(gate197inter4));
  nand2 gate1084(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1085(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1086(.a(G594), .O(gate197inter7));
  inv1  gate1087(.a(G595), .O(gate197inter8));
  nand2 gate1088(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1089(.a(s_77), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1090(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1091(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1092(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1625(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1626(.a(gate200inter0), .b(s_154), .O(gate200inter1));
  and2  gate1627(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1628(.a(s_154), .O(gate200inter3));
  inv1  gate1629(.a(s_155), .O(gate200inter4));
  nand2 gate1630(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1631(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1632(.a(G600), .O(gate200inter7));
  inv1  gate1633(.a(G601), .O(gate200inter8));
  nand2 gate1634(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1635(.a(s_155), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1636(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1637(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1638(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1849(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1850(.a(gate201inter0), .b(s_186), .O(gate201inter1));
  and2  gate1851(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1852(.a(s_186), .O(gate201inter3));
  inv1  gate1853(.a(s_187), .O(gate201inter4));
  nand2 gate1854(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1855(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1856(.a(G602), .O(gate201inter7));
  inv1  gate1857(.a(G607), .O(gate201inter8));
  nand2 gate1858(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1859(.a(s_187), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1860(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1861(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1862(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate673(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate674(.a(gate203inter0), .b(s_18), .O(gate203inter1));
  and2  gate675(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate676(.a(s_18), .O(gate203inter3));
  inv1  gate677(.a(s_19), .O(gate203inter4));
  nand2 gate678(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate679(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate680(.a(G602), .O(gate203inter7));
  inv1  gate681(.a(G612), .O(gate203inter8));
  nand2 gate682(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate683(.a(s_19), .b(gate203inter3), .O(gate203inter10));
  nor2  gate684(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate685(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate686(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1471(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1472(.a(gate204inter0), .b(s_132), .O(gate204inter1));
  and2  gate1473(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1474(.a(s_132), .O(gate204inter3));
  inv1  gate1475(.a(s_133), .O(gate204inter4));
  nand2 gate1476(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1477(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1478(.a(G607), .O(gate204inter7));
  inv1  gate1479(.a(G617), .O(gate204inter8));
  nand2 gate1480(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1481(.a(s_133), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1482(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1483(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1484(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1023(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1024(.a(gate207inter0), .b(s_68), .O(gate207inter1));
  and2  gate1025(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1026(.a(s_68), .O(gate207inter3));
  inv1  gate1027(.a(s_69), .O(gate207inter4));
  nand2 gate1028(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1029(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1030(.a(G622), .O(gate207inter7));
  inv1  gate1031(.a(G632), .O(gate207inter8));
  nand2 gate1032(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1033(.a(s_69), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1034(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1035(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1036(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1401(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1402(.a(gate213inter0), .b(s_122), .O(gate213inter1));
  and2  gate1403(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1404(.a(s_122), .O(gate213inter3));
  inv1  gate1405(.a(s_123), .O(gate213inter4));
  nand2 gate1406(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1407(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1408(.a(G602), .O(gate213inter7));
  inv1  gate1409(.a(G672), .O(gate213inter8));
  nand2 gate1410(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1411(.a(s_123), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1412(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1413(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1414(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1037(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1038(.a(gate214inter0), .b(s_70), .O(gate214inter1));
  and2  gate1039(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1040(.a(s_70), .O(gate214inter3));
  inv1  gate1041(.a(s_71), .O(gate214inter4));
  nand2 gate1042(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1043(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1044(.a(G612), .O(gate214inter7));
  inv1  gate1045(.a(G672), .O(gate214inter8));
  nand2 gate1046(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1047(.a(s_71), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1048(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1049(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1050(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate799(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate800(.a(gate222inter0), .b(s_36), .O(gate222inter1));
  and2  gate801(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate802(.a(s_36), .O(gate222inter3));
  inv1  gate803(.a(s_37), .O(gate222inter4));
  nand2 gate804(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate805(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate806(.a(G632), .O(gate222inter7));
  inv1  gate807(.a(G684), .O(gate222inter8));
  nand2 gate808(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate809(.a(s_37), .b(gate222inter3), .O(gate222inter10));
  nor2  gate810(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate811(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate812(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1457(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1458(.a(gate224inter0), .b(s_130), .O(gate224inter1));
  and2  gate1459(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1460(.a(s_130), .O(gate224inter3));
  inv1  gate1461(.a(s_131), .O(gate224inter4));
  nand2 gate1462(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1463(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1464(.a(G637), .O(gate224inter7));
  inv1  gate1465(.a(G687), .O(gate224inter8));
  nand2 gate1466(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1467(.a(s_131), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1468(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1469(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1470(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1695(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1696(.a(gate226inter0), .b(s_164), .O(gate226inter1));
  and2  gate1697(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1698(.a(s_164), .O(gate226inter3));
  inv1  gate1699(.a(s_165), .O(gate226inter4));
  nand2 gate1700(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1701(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1702(.a(G692), .O(gate226inter7));
  inv1  gate1703(.a(G693), .O(gate226inter8));
  nand2 gate1704(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1705(.a(s_165), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1706(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1707(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1708(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1233(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1234(.a(gate238inter0), .b(s_98), .O(gate238inter1));
  and2  gate1235(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1236(.a(s_98), .O(gate238inter3));
  inv1  gate1237(.a(s_99), .O(gate238inter4));
  nand2 gate1238(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1239(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1240(.a(G257), .O(gate238inter7));
  inv1  gate1241(.a(G709), .O(gate238inter8));
  nand2 gate1242(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1243(.a(s_99), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1244(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1245(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1246(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate953(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate954(.a(gate242inter0), .b(s_58), .O(gate242inter1));
  and2  gate955(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate956(.a(s_58), .O(gate242inter3));
  inv1  gate957(.a(s_59), .O(gate242inter4));
  nand2 gate958(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate959(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate960(.a(G718), .O(gate242inter7));
  inv1  gate961(.a(G730), .O(gate242inter8));
  nand2 gate962(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate963(.a(s_59), .b(gate242inter3), .O(gate242inter10));
  nor2  gate964(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate965(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate966(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate743(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate744(.a(gate244inter0), .b(s_28), .O(gate244inter1));
  and2  gate745(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate746(.a(s_28), .O(gate244inter3));
  inv1  gate747(.a(s_29), .O(gate244inter4));
  nand2 gate748(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate749(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate750(.a(G721), .O(gate244inter7));
  inv1  gate751(.a(G733), .O(gate244inter8));
  nand2 gate752(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate753(.a(s_29), .b(gate244inter3), .O(gate244inter10));
  nor2  gate754(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate755(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate756(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1653(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1654(.a(gate249inter0), .b(s_158), .O(gate249inter1));
  and2  gate1655(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1656(.a(s_158), .O(gate249inter3));
  inv1  gate1657(.a(s_159), .O(gate249inter4));
  nand2 gate1658(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1659(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1660(.a(G254), .O(gate249inter7));
  inv1  gate1661(.a(G742), .O(gate249inter8));
  nand2 gate1662(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1663(.a(s_159), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1664(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1665(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1666(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate603(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate604(.a(gate253inter0), .b(s_8), .O(gate253inter1));
  and2  gate605(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate606(.a(s_8), .O(gate253inter3));
  inv1  gate607(.a(s_9), .O(gate253inter4));
  nand2 gate608(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate609(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate610(.a(G260), .O(gate253inter7));
  inv1  gate611(.a(G748), .O(gate253inter8));
  nand2 gate612(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate613(.a(s_9), .b(gate253inter3), .O(gate253inter10));
  nor2  gate614(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate615(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate616(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate617(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate618(.a(gate254inter0), .b(s_10), .O(gate254inter1));
  and2  gate619(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate620(.a(s_10), .O(gate254inter3));
  inv1  gate621(.a(s_11), .O(gate254inter4));
  nand2 gate622(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate623(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate624(.a(G712), .O(gate254inter7));
  inv1  gate625(.a(G748), .O(gate254inter8));
  nand2 gate626(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate627(.a(s_11), .b(gate254inter3), .O(gate254inter10));
  nor2  gate628(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate629(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate630(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1093(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1094(.a(gate262inter0), .b(s_78), .O(gate262inter1));
  and2  gate1095(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1096(.a(s_78), .O(gate262inter3));
  inv1  gate1097(.a(s_79), .O(gate262inter4));
  nand2 gate1098(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1099(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1100(.a(G764), .O(gate262inter7));
  inv1  gate1101(.a(G765), .O(gate262inter8));
  nand2 gate1102(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1103(.a(s_79), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1104(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1105(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1106(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate659(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate660(.a(gate268inter0), .b(s_16), .O(gate268inter1));
  and2  gate661(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate662(.a(s_16), .O(gate268inter3));
  inv1  gate663(.a(s_17), .O(gate268inter4));
  nand2 gate664(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate665(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate666(.a(G651), .O(gate268inter7));
  inv1  gate667(.a(G779), .O(gate268inter8));
  nand2 gate668(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate669(.a(s_17), .b(gate268inter3), .O(gate268inter10));
  nor2  gate670(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate671(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate672(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate827(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate828(.a(gate272inter0), .b(s_40), .O(gate272inter1));
  and2  gate829(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate830(.a(s_40), .O(gate272inter3));
  inv1  gate831(.a(s_41), .O(gate272inter4));
  nand2 gate832(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate833(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate834(.a(G663), .O(gate272inter7));
  inv1  gate835(.a(G791), .O(gate272inter8));
  nand2 gate836(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate837(.a(s_41), .b(gate272inter3), .O(gate272inter10));
  nor2  gate838(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate839(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate840(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1863(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1864(.a(gate273inter0), .b(s_188), .O(gate273inter1));
  and2  gate1865(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1866(.a(s_188), .O(gate273inter3));
  inv1  gate1867(.a(s_189), .O(gate273inter4));
  nand2 gate1868(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1869(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1870(.a(G642), .O(gate273inter7));
  inv1  gate1871(.a(G794), .O(gate273inter8));
  nand2 gate1872(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1873(.a(s_189), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1874(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1875(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1876(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1443(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1444(.a(gate275inter0), .b(s_128), .O(gate275inter1));
  and2  gate1445(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1446(.a(s_128), .O(gate275inter3));
  inv1  gate1447(.a(s_129), .O(gate275inter4));
  nand2 gate1448(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1449(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1450(.a(G645), .O(gate275inter7));
  inv1  gate1451(.a(G797), .O(gate275inter8));
  nand2 gate1452(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1453(.a(s_129), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1454(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1455(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1456(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1163(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1164(.a(gate285inter0), .b(s_88), .O(gate285inter1));
  and2  gate1165(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1166(.a(s_88), .O(gate285inter3));
  inv1  gate1167(.a(s_89), .O(gate285inter4));
  nand2 gate1168(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1169(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1170(.a(G660), .O(gate285inter7));
  inv1  gate1171(.a(G812), .O(gate285inter8));
  nand2 gate1172(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1173(.a(s_89), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1174(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1175(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1176(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1891(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1892(.a(gate287inter0), .b(s_192), .O(gate287inter1));
  and2  gate1893(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1894(.a(s_192), .O(gate287inter3));
  inv1  gate1895(.a(s_193), .O(gate287inter4));
  nand2 gate1896(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1897(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1898(.a(G663), .O(gate287inter7));
  inv1  gate1899(.a(G815), .O(gate287inter8));
  nand2 gate1900(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1901(.a(s_193), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1902(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1903(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1904(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate981(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate982(.a(gate288inter0), .b(s_62), .O(gate288inter1));
  and2  gate983(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate984(.a(s_62), .O(gate288inter3));
  inv1  gate985(.a(s_63), .O(gate288inter4));
  nand2 gate986(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate987(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate988(.a(G791), .O(gate288inter7));
  inv1  gate989(.a(G815), .O(gate288inter8));
  nand2 gate990(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate991(.a(s_63), .b(gate288inter3), .O(gate288inter10));
  nor2  gate992(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate993(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate994(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate645(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate646(.a(gate289inter0), .b(s_14), .O(gate289inter1));
  and2  gate647(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate648(.a(s_14), .O(gate289inter3));
  inv1  gate649(.a(s_15), .O(gate289inter4));
  nand2 gate650(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate651(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate652(.a(G818), .O(gate289inter7));
  inv1  gate653(.a(G819), .O(gate289inter8));
  nand2 gate654(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate655(.a(s_15), .b(gate289inter3), .O(gate289inter10));
  nor2  gate656(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate657(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate658(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate575(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate576(.a(gate387inter0), .b(s_4), .O(gate387inter1));
  and2  gate577(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate578(.a(s_4), .O(gate387inter3));
  inv1  gate579(.a(s_5), .O(gate387inter4));
  nand2 gate580(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate581(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate582(.a(G1), .O(gate387inter7));
  inv1  gate583(.a(G1036), .O(gate387inter8));
  nand2 gate584(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate585(.a(s_5), .b(gate387inter3), .O(gate387inter10));
  nor2  gate586(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate587(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate588(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1373(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1374(.a(gate388inter0), .b(s_118), .O(gate388inter1));
  and2  gate1375(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1376(.a(s_118), .O(gate388inter3));
  inv1  gate1377(.a(s_119), .O(gate388inter4));
  nand2 gate1378(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1379(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1380(.a(G2), .O(gate388inter7));
  inv1  gate1381(.a(G1039), .O(gate388inter8));
  nand2 gate1382(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1383(.a(s_119), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1384(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1385(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1386(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1429(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1430(.a(gate389inter0), .b(s_126), .O(gate389inter1));
  and2  gate1431(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1432(.a(s_126), .O(gate389inter3));
  inv1  gate1433(.a(s_127), .O(gate389inter4));
  nand2 gate1434(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1435(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1436(.a(G3), .O(gate389inter7));
  inv1  gate1437(.a(G1042), .O(gate389inter8));
  nand2 gate1438(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1439(.a(s_127), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1440(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1441(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1442(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate841(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate842(.a(gate392inter0), .b(s_42), .O(gate392inter1));
  and2  gate843(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate844(.a(s_42), .O(gate392inter3));
  inv1  gate845(.a(s_43), .O(gate392inter4));
  nand2 gate846(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate847(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate848(.a(G6), .O(gate392inter7));
  inv1  gate849(.a(G1051), .O(gate392inter8));
  nand2 gate850(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate851(.a(s_43), .b(gate392inter3), .O(gate392inter10));
  nor2  gate852(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate853(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate854(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1107(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1108(.a(gate393inter0), .b(s_80), .O(gate393inter1));
  and2  gate1109(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1110(.a(s_80), .O(gate393inter3));
  inv1  gate1111(.a(s_81), .O(gate393inter4));
  nand2 gate1112(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1113(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1114(.a(G7), .O(gate393inter7));
  inv1  gate1115(.a(G1054), .O(gate393inter8));
  nand2 gate1116(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1117(.a(s_81), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1118(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1119(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1120(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1723(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1724(.a(gate395inter0), .b(s_168), .O(gate395inter1));
  and2  gate1725(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1726(.a(s_168), .O(gate395inter3));
  inv1  gate1727(.a(s_169), .O(gate395inter4));
  nand2 gate1728(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1729(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1730(.a(G9), .O(gate395inter7));
  inv1  gate1731(.a(G1060), .O(gate395inter8));
  nand2 gate1732(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1733(.a(s_169), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1734(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1735(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1736(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate1065(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1066(.a(gate396inter0), .b(s_74), .O(gate396inter1));
  and2  gate1067(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1068(.a(s_74), .O(gate396inter3));
  inv1  gate1069(.a(s_75), .O(gate396inter4));
  nand2 gate1070(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1071(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1072(.a(G10), .O(gate396inter7));
  inv1  gate1073(.a(G1063), .O(gate396inter8));
  nand2 gate1074(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1075(.a(s_75), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1076(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1077(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1078(.a(gate396inter12), .b(gate396inter1), .O(G1159));

  xor2  gate729(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate730(.a(gate397inter0), .b(s_26), .O(gate397inter1));
  and2  gate731(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate732(.a(s_26), .O(gate397inter3));
  inv1  gate733(.a(s_27), .O(gate397inter4));
  nand2 gate734(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate735(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate736(.a(G11), .O(gate397inter7));
  inv1  gate737(.a(G1066), .O(gate397inter8));
  nand2 gate738(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate739(.a(s_27), .b(gate397inter3), .O(gate397inter10));
  nor2  gate740(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate741(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate742(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1779(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1780(.a(gate398inter0), .b(s_176), .O(gate398inter1));
  and2  gate1781(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1782(.a(s_176), .O(gate398inter3));
  inv1  gate1783(.a(s_177), .O(gate398inter4));
  nand2 gate1784(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1785(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1786(.a(G12), .O(gate398inter7));
  inv1  gate1787(.a(G1069), .O(gate398inter8));
  nand2 gate1788(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1789(.a(s_177), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1790(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1791(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1792(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1961(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1962(.a(gate408inter0), .b(s_202), .O(gate408inter1));
  and2  gate1963(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1964(.a(s_202), .O(gate408inter3));
  inv1  gate1965(.a(s_203), .O(gate408inter4));
  nand2 gate1966(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1967(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1968(.a(G22), .O(gate408inter7));
  inv1  gate1969(.a(G1099), .O(gate408inter8));
  nand2 gate1970(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1971(.a(s_203), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1972(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1973(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1974(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1247(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1248(.a(gate409inter0), .b(s_100), .O(gate409inter1));
  and2  gate1249(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1250(.a(s_100), .O(gate409inter3));
  inv1  gate1251(.a(s_101), .O(gate409inter4));
  nand2 gate1252(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1253(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1254(.a(G23), .O(gate409inter7));
  inv1  gate1255(.a(G1102), .O(gate409inter8));
  nand2 gate1256(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1257(.a(s_101), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1258(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1259(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1260(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate883(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate884(.a(gate411inter0), .b(s_48), .O(gate411inter1));
  and2  gate885(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate886(.a(s_48), .O(gate411inter3));
  inv1  gate887(.a(s_49), .O(gate411inter4));
  nand2 gate888(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate889(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate890(.a(G25), .O(gate411inter7));
  inv1  gate891(.a(G1108), .O(gate411inter8));
  nand2 gate892(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate893(.a(s_49), .b(gate411inter3), .O(gate411inter10));
  nor2  gate894(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate895(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate896(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1877(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1878(.a(gate414inter0), .b(s_190), .O(gate414inter1));
  and2  gate1879(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1880(.a(s_190), .O(gate414inter3));
  inv1  gate1881(.a(s_191), .O(gate414inter4));
  nand2 gate1882(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1883(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1884(.a(G28), .O(gate414inter7));
  inv1  gate1885(.a(G1117), .O(gate414inter8));
  nand2 gate1886(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1887(.a(s_191), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1888(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1889(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1890(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate561(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate562(.a(gate415inter0), .b(s_2), .O(gate415inter1));
  and2  gate563(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate564(.a(s_2), .O(gate415inter3));
  inv1  gate565(.a(s_3), .O(gate415inter4));
  nand2 gate566(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate567(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate568(.a(G29), .O(gate415inter7));
  inv1  gate569(.a(G1120), .O(gate415inter8));
  nand2 gate570(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate571(.a(s_3), .b(gate415inter3), .O(gate415inter10));
  nor2  gate572(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate573(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate574(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1177(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1178(.a(gate417inter0), .b(s_90), .O(gate417inter1));
  and2  gate1179(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1180(.a(s_90), .O(gate417inter3));
  inv1  gate1181(.a(s_91), .O(gate417inter4));
  nand2 gate1182(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1183(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1184(.a(G31), .O(gate417inter7));
  inv1  gate1185(.a(G1126), .O(gate417inter8));
  nand2 gate1186(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1187(.a(s_91), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1188(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1189(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1190(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate967(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate968(.a(gate433inter0), .b(s_60), .O(gate433inter1));
  and2  gate969(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate970(.a(s_60), .O(gate433inter3));
  inv1  gate971(.a(s_61), .O(gate433inter4));
  nand2 gate972(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate973(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate974(.a(G8), .O(gate433inter7));
  inv1  gate975(.a(G1153), .O(gate433inter8));
  nand2 gate976(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate977(.a(s_61), .b(gate433inter3), .O(gate433inter10));
  nor2  gate978(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate979(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate980(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1681(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1682(.a(gate434inter0), .b(s_162), .O(gate434inter1));
  and2  gate1683(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1684(.a(s_162), .O(gate434inter3));
  inv1  gate1685(.a(s_163), .O(gate434inter4));
  nand2 gate1686(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1687(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1688(.a(G1057), .O(gate434inter7));
  inv1  gate1689(.a(G1153), .O(gate434inter8));
  nand2 gate1690(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1691(.a(s_163), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1692(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1693(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1694(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1751(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1752(.a(gate440inter0), .b(s_172), .O(gate440inter1));
  and2  gate1753(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1754(.a(s_172), .O(gate440inter3));
  inv1  gate1755(.a(s_173), .O(gate440inter4));
  nand2 gate1756(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1757(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1758(.a(G1066), .O(gate440inter7));
  inv1  gate1759(.a(G1162), .O(gate440inter8));
  nand2 gate1760(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1761(.a(s_173), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1762(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1763(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1764(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate757(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate758(.a(gate444inter0), .b(s_30), .O(gate444inter1));
  and2  gate759(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate760(.a(s_30), .O(gate444inter3));
  inv1  gate761(.a(s_31), .O(gate444inter4));
  nand2 gate762(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate763(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate764(.a(G1072), .O(gate444inter7));
  inv1  gate765(.a(G1168), .O(gate444inter8));
  nand2 gate766(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate767(.a(s_31), .b(gate444inter3), .O(gate444inter10));
  nor2  gate768(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate769(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate770(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate631(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate632(.a(gate451inter0), .b(s_12), .O(gate451inter1));
  and2  gate633(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate634(.a(s_12), .O(gate451inter3));
  inv1  gate635(.a(s_13), .O(gate451inter4));
  nand2 gate636(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate637(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate638(.a(G17), .O(gate451inter7));
  inv1  gate639(.a(G1180), .O(gate451inter8));
  nand2 gate640(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate641(.a(s_13), .b(gate451inter3), .O(gate451inter10));
  nor2  gate642(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate643(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate644(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1611(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1612(.a(gate452inter0), .b(s_152), .O(gate452inter1));
  and2  gate1613(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1614(.a(s_152), .O(gate452inter3));
  inv1  gate1615(.a(s_153), .O(gate452inter4));
  nand2 gate1616(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1617(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1618(.a(G1084), .O(gate452inter7));
  inv1  gate1619(.a(G1180), .O(gate452inter8));
  nand2 gate1620(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1621(.a(s_153), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1622(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1623(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1624(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate1737(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1738(.a(gate453inter0), .b(s_170), .O(gate453inter1));
  and2  gate1739(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1740(.a(s_170), .O(gate453inter3));
  inv1  gate1741(.a(s_171), .O(gate453inter4));
  nand2 gate1742(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1743(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1744(.a(G18), .O(gate453inter7));
  inv1  gate1745(.a(G1183), .O(gate453inter8));
  nand2 gate1746(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1747(.a(s_171), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1748(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1749(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1750(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1765(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1766(.a(gate454inter0), .b(s_174), .O(gate454inter1));
  and2  gate1767(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1768(.a(s_174), .O(gate454inter3));
  inv1  gate1769(.a(s_175), .O(gate454inter4));
  nand2 gate1770(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1771(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1772(.a(G1087), .O(gate454inter7));
  inv1  gate1773(.a(G1183), .O(gate454inter8));
  nand2 gate1774(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1775(.a(s_175), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1776(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1777(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1778(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1569(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1570(.a(gate455inter0), .b(s_146), .O(gate455inter1));
  and2  gate1571(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1572(.a(s_146), .O(gate455inter3));
  inv1  gate1573(.a(s_147), .O(gate455inter4));
  nand2 gate1574(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1575(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1576(.a(G19), .O(gate455inter7));
  inv1  gate1577(.a(G1186), .O(gate455inter8));
  nand2 gate1578(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1579(.a(s_147), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1580(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1581(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1582(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1135(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1136(.a(gate456inter0), .b(s_84), .O(gate456inter1));
  and2  gate1137(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1138(.a(s_84), .O(gate456inter3));
  inv1  gate1139(.a(s_85), .O(gate456inter4));
  nand2 gate1140(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1141(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1142(.a(G1090), .O(gate456inter7));
  inv1  gate1143(.a(G1186), .O(gate456inter8));
  nand2 gate1144(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1145(.a(s_85), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1146(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1147(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1148(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate2059(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2060(.a(gate462inter0), .b(s_216), .O(gate462inter1));
  and2  gate2061(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2062(.a(s_216), .O(gate462inter3));
  inv1  gate2063(.a(s_217), .O(gate462inter4));
  nand2 gate2064(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2065(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2066(.a(G1099), .O(gate462inter7));
  inv1  gate2067(.a(G1195), .O(gate462inter8));
  nand2 gate2068(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2069(.a(s_217), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2070(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2071(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2072(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate813(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate814(.a(gate469inter0), .b(s_38), .O(gate469inter1));
  and2  gate815(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate816(.a(s_38), .O(gate469inter3));
  inv1  gate817(.a(s_39), .O(gate469inter4));
  nand2 gate818(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate819(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate820(.a(G26), .O(gate469inter7));
  inv1  gate821(.a(G1207), .O(gate469inter8));
  nand2 gate822(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate823(.a(s_39), .b(gate469inter3), .O(gate469inter10));
  nor2  gate824(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate825(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate826(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1583(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1584(.a(gate471inter0), .b(s_148), .O(gate471inter1));
  and2  gate1585(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1586(.a(s_148), .O(gate471inter3));
  inv1  gate1587(.a(s_149), .O(gate471inter4));
  nand2 gate1588(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1589(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1590(.a(G27), .O(gate471inter7));
  inv1  gate1591(.a(G1210), .O(gate471inter8));
  nand2 gate1592(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1593(.a(s_149), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1594(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1595(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1596(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1555(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1556(.a(gate482inter0), .b(s_144), .O(gate482inter1));
  and2  gate1557(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1558(.a(s_144), .O(gate482inter3));
  inv1  gate1559(.a(s_145), .O(gate482inter4));
  nand2 gate1560(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1561(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1562(.a(G1129), .O(gate482inter7));
  inv1  gate1563(.a(G1225), .O(gate482inter8));
  nand2 gate1564(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1565(.a(s_145), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1566(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1567(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1568(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1905(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1906(.a(gate485inter0), .b(s_194), .O(gate485inter1));
  and2  gate1907(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1908(.a(s_194), .O(gate485inter3));
  inv1  gate1909(.a(s_195), .O(gate485inter4));
  nand2 gate1910(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1911(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1912(.a(G1232), .O(gate485inter7));
  inv1  gate1913(.a(G1233), .O(gate485inter8));
  nand2 gate1914(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1915(.a(s_195), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1916(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1917(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1918(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1415(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1416(.a(gate497inter0), .b(s_124), .O(gate497inter1));
  and2  gate1417(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1418(.a(s_124), .O(gate497inter3));
  inv1  gate1419(.a(s_125), .O(gate497inter4));
  nand2 gate1420(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1421(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1422(.a(G1256), .O(gate497inter7));
  inv1  gate1423(.a(G1257), .O(gate497inter8));
  nand2 gate1424(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1425(.a(s_125), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1426(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1427(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1428(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1793(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1794(.a(gate500inter0), .b(s_178), .O(gate500inter1));
  and2  gate1795(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1796(.a(s_178), .O(gate500inter3));
  inv1  gate1797(.a(s_179), .O(gate500inter4));
  nand2 gate1798(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1799(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1800(.a(G1262), .O(gate500inter7));
  inv1  gate1801(.a(G1263), .O(gate500inter8));
  nand2 gate1802(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1803(.a(s_179), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1804(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1805(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1806(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1919(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1920(.a(gate505inter0), .b(s_196), .O(gate505inter1));
  and2  gate1921(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1922(.a(s_196), .O(gate505inter3));
  inv1  gate1923(.a(s_197), .O(gate505inter4));
  nand2 gate1924(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1925(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1926(.a(G1272), .O(gate505inter7));
  inv1  gate1927(.a(G1273), .O(gate505inter8));
  nand2 gate1928(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1929(.a(s_197), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1930(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1931(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1932(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1289(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1290(.a(gate507inter0), .b(s_106), .O(gate507inter1));
  and2  gate1291(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1292(.a(s_106), .O(gate507inter3));
  inv1  gate1293(.a(s_107), .O(gate507inter4));
  nand2 gate1294(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1295(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1296(.a(G1276), .O(gate507inter7));
  inv1  gate1297(.a(G1277), .O(gate507inter8));
  nand2 gate1298(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1299(.a(s_107), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1300(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1301(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1302(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1499(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1500(.a(gate510inter0), .b(s_136), .O(gate510inter1));
  and2  gate1501(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1502(.a(s_136), .O(gate510inter3));
  inv1  gate1503(.a(s_137), .O(gate510inter4));
  nand2 gate1504(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1505(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1506(.a(G1282), .O(gate510inter7));
  inv1  gate1507(.a(G1283), .O(gate510inter8));
  nand2 gate1508(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1509(.a(s_137), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1510(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1511(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1512(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate2073(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2074(.a(gate512inter0), .b(s_218), .O(gate512inter1));
  and2  gate2075(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2076(.a(s_218), .O(gate512inter3));
  inv1  gate2077(.a(s_219), .O(gate512inter4));
  nand2 gate2078(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2079(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2080(.a(G1286), .O(gate512inter7));
  inv1  gate2081(.a(G1287), .O(gate512inter8));
  nand2 gate2082(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2083(.a(s_219), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2084(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2085(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2086(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1947(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1948(.a(gate514inter0), .b(s_200), .O(gate514inter1));
  and2  gate1949(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1950(.a(s_200), .O(gate514inter3));
  inv1  gate1951(.a(s_201), .O(gate514inter4));
  nand2 gate1952(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1953(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1954(.a(G1290), .O(gate514inter7));
  inv1  gate1955(.a(G1291), .O(gate514inter8));
  nand2 gate1956(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1957(.a(s_201), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1958(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1959(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1960(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule