module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;
wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877, gate298inter0, gate298inter1, gate298inter2, gate298inter3, gate298inter4, gate298inter5, gate298inter6, gate298inter7, gate298inter8, gate298inter9, gate298inter10, gate298inter11, gate298inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate299inter0, gate299inter1, gate299inter2, gate299inter3, gate299inter4, gate299inter5, gate299inter6, gate299inter7, gate299inter8, gate299inter9, gate299inter10, gate299inter11, gate299inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate305inter0, gate305inter1, gate305inter2, gate305inter3, gate305inter4, gate305inter5, gate305inter6, gate305inter7, gate305inter8, gate305inter9, gate305inter10, gate305inter11, gate305inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate316inter0, gate316inter1, gate316inter2, gate316inter3, gate316inter4, gate316inter5, gate316inter6, gate316inter7, gate316inter8, gate316inter9, gate316inter10, gate316inter11, gate316inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate335inter0, gate335inter1, gate335inter2, gate335inter3, gate335inter4, gate335inter5, gate335inter6, gate335inter7, gate335inter8, gate335inter9, gate335inter10, gate335inter11, gate335inter12, gate363inter0, gate363inter1, gate363inter2, gate363inter3, gate363inter4, gate363inter5, gate363inter6, gate363inter7, gate363inter8, gate363inter9, gate363inter10, gate363inter11, gate363inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate333inter0, gate333inter1, gate333inter2, gate333inter3, gate333inter4, gate333inter5, gate333inter6, gate333inter7, gate333inter8, gate333inter9, gate333inter10, gate333inter11, gate333inter12, gate322inter0, gate322inter1, gate322inter2, gate322inter3, gate322inter4, gate322inter5, gate322inter6, gate322inter7, gate322inter8, gate322inter9, gate322inter10, gate322inter11, gate322inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate312inter0, gate312inter1, gate312inter2, gate312inter3, gate312inter4, gate312inter5, gate312inter6, gate312inter7, gate312inter8, gate312inter9, gate312inter10, gate312inter11, gate312inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate313inter0, gate313inter1, gate313inter2, gate313inter3, gate313inter4, gate313inter5, gate313inter6, gate313inter7, gate313inter8, gate313inter9, gate313inter10, gate313inter11, gate313inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate362inter0, gate362inter1, gate362inter2, gate362inter3, gate362inter4, gate362inter5, gate362inter6, gate362inter7, gate362inter8, gate362inter9, gate362inter10, gate362inter11, gate362inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12;


nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );

  xor2  gate524(.a(N96), .b(N91), .O(gate20inter0));
  nand2 gate525(.a(gate20inter0), .b(s_20), .O(gate20inter1));
  and2  gate526(.a(N96), .b(N91), .O(gate20inter2));
  inv1  gate527(.a(s_20), .O(gate20inter3));
  inv1  gate528(.a(s_21), .O(gate20inter4));
  nand2 gate529(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate530(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate531(.a(N91), .O(gate20inter7));
  inv1  gate532(.a(N96), .O(gate20inter8));
  nand2 gate533(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate534(.a(s_21), .b(gate20inter3), .O(gate20inter10));
  nor2  gate535(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate536(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate537(.a(gate20inter12), .b(gate20inter1), .O(N301));
or2 gate21( .a(N91), .b(N96), .O(N302) );
nand2 gate22( .a(N101), .b(N106), .O(N303) );
or2 gate23( .a(N101), .b(N106), .O(N304) );

  xor2  gate496(.a(N116), .b(N111), .O(gate24inter0));
  nand2 gate497(.a(gate24inter0), .b(s_16), .O(gate24inter1));
  and2  gate498(.a(N116), .b(N111), .O(gate24inter2));
  inv1  gate499(.a(s_16), .O(gate24inter3));
  inv1  gate500(.a(s_17), .O(gate24inter4));
  nand2 gate501(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate502(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate503(.a(N111), .O(gate24inter7));
  inv1  gate504(.a(N116), .O(gate24inter8));
  nand2 gate505(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate506(.a(s_17), .b(gate24inter3), .O(gate24inter10));
  nor2  gate507(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate508(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate509(.a(gate24inter12), .b(gate24inter1), .O(N305));
or2 gate25( .a(N111), .b(N116), .O(N306) );

  xor2  gate888(.a(N126), .b(N121), .O(gate26inter0));
  nand2 gate889(.a(gate26inter0), .b(s_72), .O(gate26inter1));
  and2  gate890(.a(N126), .b(N121), .O(gate26inter2));
  inv1  gate891(.a(s_72), .O(gate26inter3));
  inv1  gate892(.a(s_73), .O(gate26inter4));
  nand2 gate893(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate894(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate895(.a(N121), .O(gate26inter7));
  inv1  gate896(.a(N126), .O(gate26inter8));
  nand2 gate897(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate898(.a(s_73), .b(gate26inter3), .O(gate26inter10));
  nor2  gate899(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate900(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate901(.a(gate26inter12), .b(gate26inter1), .O(N307));
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );
nand2 gate33( .a(N59), .b(N156), .O(N319) );
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17), .b(N42), .O(N323) );
nand2 gate36( .a(N159), .b(N165), .O(N324) );
or2 gate37( .a(N159), .b(N165), .O(N325) );

  xor2  gate790(.a(N177), .b(N171), .O(gate38inter0));
  nand2 gate791(.a(gate38inter0), .b(s_58), .O(gate38inter1));
  and2  gate792(.a(N177), .b(N171), .O(gate38inter2));
  inv1  gate793(.a(s_58), .O(gate38inter3));
  inv1  gate794(.a(s_59), .O(gate38inter4));
  nand2 gate795(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate796(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate797(.a(N171), .O(gate38inter7));
  inv1  gate798(.a(N177), .O(gate38inter8));
  nand2 gate799(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate800(.a(s_59), .b(gate38inter3), .O(gate38inter10));
  nor2  gate801(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate802(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate803(.a(gate38inter12), .b(gate38inter1), .O(N326));
or2 gate39( .a(N171), .b(N177), .O(N327) );

  xor2  gate916(.a(N189), .b(N183), .O(gate40inter0));
  nand2 gate917(.a(gate40inter0), .b(s_76), .O(gate40inter1));
  and2  gate918(.a(N189), .b(N183), .O(gate40inter2));
  inv1  gate919(.a(s_76), .O(gate40inter3));
  inv1  gate920(.a(s_77), .O(gate40inter4));
  nand2 gate921(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate922(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate923(.a(N183), .O(gate40inter7));
  inv1  gate924(.a(N189), .O(gate40inter8));
  nand2 gate925(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate926(.a(s_77), .b(gate40inter3), .O(gate40inter10));
  nor2  gate927(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate928(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate929(.a(gate40inter12), .b(gate40inter1), .O(N328));
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
and2 gate49( .a(N255), .b(N259), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );

  xor2  gate1070(.a(N284), .b(N280), .O(gate60inter0));
  nand2 gate1071(.a(gate60inter0), .b(s_98), .O(gate60inter1));
  and2  gate1072(.a(N284), .b(N280), .O(gate60inter2));
  inv1  gate1073(.a(s_98), .O(gate60inter3));
  inv1  gate1074(.a(s_99), .O(gate60inter4));
  nand2 gate1075(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1076(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1077(.a(N280), .O(gate60inter7));
  inv1  gate1078(.a(N284), .O(gate60inter8));
  nand2 gate1079(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1080(.a(s_99), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1081(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1082(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1083(.a(gate60inter12), .b(gate60inter1), .O(N348));
or2 gate61( .a(N280), .b(N285), .O(N349) );
or2 gate62( .a(N280), .b(N286), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );

  xor2  gate776(.a(N298), .b(N89), .O(gate67inter0));
  nand2 gate777(.a(gate67inter0), .b(s_56), .O(gate67inter1));
  and2  gate778(.a(N298), .b(N89), .O(gate67inter2));
  inv1  gate779(.a(s_56), .O(gate67inter3));
  inv1  gate780(.a(s_57), .O(gate67inter4));
  nand2 gate781(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate782(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate783(.a(N89), .O(gate67inter7));
  inv1  gate784(.a(N298), .O(gate67inter8));
  nand2 gate785(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate786(.a(s_57), .b(gate67inter3), .O(gate67inter10));
  nor2  gate787(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate788(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate789(.a(gate67inter12), .b(gate67inter1), .O(N355));
and2 gate68( .a(N90), .b(N298), .O(N356) );

  xor2  gate1014(.a(N302), .b(N301), .O(gate69inter0));
  nand2 gate1015(.a(gate69inter0), .b(s_90), .O(gate69inter1));
  and2  gate1016(.a(N302), .b(N301), .O(gate69inter2));
  inv1  gate1017(.a(s_90), .O(gate69inter3));
  inv1  gate1018(.a(s_91), .O(gate69inter4));
  nand2 gate1019(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1020(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1021(.a(N301), .O(gate69inter7));
  inv1  gate1022(.a(N302), .O(gate69inter8));
  nand2 gate1023(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1024(.a(s_91), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1025(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1026(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1027(.a(gate69inter12), .b(gate69inter1), .O(N357));

  xor2  gate874(.a(N304), .b(N303), .O(gate70inter0));
  nand2 gate875(.a(gate70inter0), .b(s_70), .O(gate70inter1));
  and2  gate876(.a(N304), .b(N303), .O(gate70inter2));
  inv1  gate877(.a(s_70), .O(gate70inter3));
  inv1  gate878(.a(s_71), .O(gate70inter4));
  nand2 gate879(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate880(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate881(.a(N303), .O(gate70inter7));
  inv1  gate882(.a(N304), .O(gate70inter8));
  nand2 gate883(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate884(.a(s_71), .b(gate70inter3), .O(gate70inter10));
  nor2  gate885(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate886(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate887(.a(gate70inter12), .b(gate70inter1), .O(N360));

  xor2  gate944(.a(N306), .b(N305), .O(gate71inter0));
  nand2 gate945(.a(gate71inter0), .b(s_80), .O(gate71inter1));
  and2  gate946(.a(N306), .b(N305), .O(gate71inter2));
  inv1  gate947(.a(s_80), .O(gate71inter3));
  inv1  gate948(.a(s_81), .O(gate71inter4));
  nand2 gate949(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate950(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate951(.a(N305), .O(gate71inter7));
  inv1  gate952(.a(N306), .O(gate71inter8));
  nand2 gate953(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate954(.a(s_81), .b(gate71inter3), .O(gate71inter10));
  nor2  gate955(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate956(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate957(.a(gate71inter12), .b(gate71inter1), .O(N363));

  xor2  gate818(.a(N308), .b(N307), .O(gate72inter0));
  nand2 gate819(.a(gate72inter0), .b(s_62), .O(gate72inter1));
  and2  gate820(.a(N308), .b(N307), .O(gate72inter2));
  inv1  gate821(.a(s_62), .O(gate72inter3));
  inv1  gate822(.a(s_63), .O(gate72inter4));
  nand2 gate823(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate824(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate825(.a(N307), .O(gate72inter7));
  inv1  gate826(.a(N308), .O(gate72inter8));
  nand2 gate827(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate828(.a(s_63), .b(gate72inter3), .O(gate72inter10));
  nor2  gate829(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate830(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate831(.a(gate72inter12), .b(gate72inter1), .O(N366));
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );
nand2 gate76( .a(N326), .b(N327), .O(N379) );
nand2 gate77( .a(N328), .b(N329), .O(N382) );

  xor2  gate398(.a(N331), .b(N330), .O(gate78inter0));
  nand2 gate399(.a(gate78inter0), .b(s_2), .O(gate78inter1));
  and2  gate400(.a(N331), .b(N330), .O(gate78inter2));
  inv1  gate401(.a(s_2), .O(gate78inter3));
  inv1  gate402(.a(s_3), .O(gate78inter4));
  nand2 gate403(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate404(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate405(.a(N330), .O(gate78inter7));
  inv1  gate406(.a(N331), .O(gate78inter8));
  nand2 gate407(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate408(.a(s_3), .b(gate78inter3), .O(gate78inter10));
  nor2  gate409(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate410(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate411(.a(gate78inter12), .b(gate78inter1), .O(N385));
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );

  xor2  gate860(.a(N352), .b(N347), .O(gate96inter0));
  nand2 gate861(.a(gate96inter0), .b(s_68), .O(gate96inter1));
  and2  gate862(.a(N352), .b(N347), .O(gate96inter2));
  inv1  gate863(.a(s_68), .O(gate96inter3));
  inv1  gate864(.a(s_69), .O(gate96inter4));
  nand2 gate865(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate866(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate867(.a(N347), .O(gate96inter7));
  inv1  gate868(.a(N352), .O(gate96inter8));
  nand2 gate869(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate870(.a(s_69), .b(gate96inter3), .O(gate96inter10));
  nor2  gate871(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate872(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate873(.a(gate96inter12), .b(gate96inter1), .O(N410));
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );

  xor2  gate426(.a(N425), .b(N406), .O(gate126inter0));
  nand2 gate427(.a(gate126inter0), .b(s_6), .O(gate126inter1));
  and2  gate428(.a(N425), .b(N406), .O(gate126inter2));
  inv1  gate429(.a(s_6), .O(gate126inter3));
  inv1  gate430(.a(s_7), .O(gate126inter4));
  nand2 gate431(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate432(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate433(.a(N406), .O(gate126inter7));
  inv1  gate434(.a(N425), .O(gate126inter8));
  nand2 gate435(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate436(.a(s_7), .b(gate126inter3), .O(gate126inter10));
  nor2  gate437(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate438(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate439(.a(gate126inter12), .b(gate126inter1), .O(N460));

  xor2  gate692(.a(N426), .b(N409), .O(gate127inter0));
  nand2 gate693(.a(gate127inter0), .b(s_44), .O(gate127inter1));
  and2  gate694(.a(N426), .b(N409), .O(gate127inter2));
  inv1  gate695(.a(s_44), .O(gate127inter3));
  inv1  gate696(.a(s_45), .O(gate127inter4));
  nand2 gate697(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate698(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate699(.a(N409), .O(gate127inter7));
  inv1  gate700(.a(N426), .O(gate127inter8));
  nand2 gate701(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate702(.a(s_45), .b(gate127inter3), .O(gate127inter10));
  nor2  gate703(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate704(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate705(.a(gate127inter12), .b(gate127inter1), .O(N463));
nand2 gate128( .a(N442), .b(N410), .O(N466) );
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );

  xor2  gate846(.a(N1), .b(N443), .O(gate137inter0));
  nand2 gate847(.a(gate137inter0), .b(s_66), .O(gate137inter1));
  and2  gate848(.a(N1), .b(N443), .O(gate137inter2));
  inv1  gate849(.a(s_66), .O(gate137inter3));
  inv1  gate850(.a(s_67), .O(gate137inter4));
  nand2 gate851(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate852(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate853(.a(N443), .O(gate137inter7));
  inv1  gate854(.a(N1), .O(gate137inter8));
  nand2 gate855(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate856(.a(s_67), .b(gate137inter3), .O(gate137inter10));
  nor2  gate857(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate858(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate859(.a(gate137inter12), .b(gate137inter1), .O(N483));
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );

  xor2  gate538(.a(N444), .b(N413), .O(gate142inter0));
  nand2 gate539(.a(gate142inter0), .b(s_22), .O(gate142inter1));
  and2  gate540(.a(N444), .b(N413), .O(gate142inter2));
  inv1  gate541(.a(s_22), .O(gate142inter3));
  inv1  gate542(.a(s_23), .O(gate142inter4));
  nand2 gate543(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate544(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate545(.a(N413), .O(gate142inter7));
  inv1  gate546(.a(N444), .O(gate142inter8));
  nand2 gate547(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate548(.a(s_23), .b(gate142inter3), .O(gate142inter10));
  nor2  gate549(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate550(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate551(.a(gate142inter12), .b(gate142inter1), .O(N492));

  xor2  gate804(.a(N445), .b(N416), .O(gate143inter0));
  nand2 gate805(.a(gate143inter0), .b(s_60), .O(gate143inter1));
  and2  gate806(.a(N445), .b(N416), .O(gate143inter2));
  inv1  gate807(.a(s_60), .O(gate143inter3));
  inv1  gate808(.a(s_61), .O(gate143inter4));
  nand2 gate809(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate810(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate811(.a(N416), .O(gate143inter7));
  inv1  gate812(.a(N445), .O(gate143inter8));
  nand2 gate813(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate814(.a(s_61), .b(gate143inter3), .O(gate143inter10));
  nor2  gate815(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate816(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate817(.a(gate143inter12), .b(gate143inter1), .O(N495));
nand2 gate144( .a(N130), .b(N460), .O(N498) );
or2 gate145( .a(N130), .b(N460), .O(N499) );

  xor2  gate552(.a(N135), .b(N463), .O(gate146inter0));
  nand2 gate553(.a(gate146inter0), .b(s_24), .O(gate146inter1));
  and2  gate554(.a(N135), .b(N463), .O(gate146inter2));
  inv1  gate555(.a(s_24), .O(gate146inter3));
  inv1  gate556(.a(s_25), .O(gate146inter4));
  nand2 gate557(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate558(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate559(.a(N463), .O(gate146inter7));
  inv1  gate560(.a(N135), .O(gate146inter8));
  nand2 gate561(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate562(.a(s_25), .b(gate146inter3), .O(gate146inter10));
  nor2  gate563(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate564(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate565(.a(gate146inter12), .b(gate146inter1), .O(N500));
or2 gate147( .a(N463), .b(N135), .O(N501) );
and2 gate148( .a(N91), .b(N466), .O(N502) );
nor2 gate149( .a(N475), .b(N476), .O(N503) );
and2 gate150( .a(N96), .b(N466), .O(N504) );
nor2 gate151( .a(N477), .b(N478), .O(N505) );
and2 gate152( .a(N101), .b(N466), .O(N506) );
nor2 gate153( .a(N479), .b(N480), .O(N507) );
and2 gate154( .a(N106), .b(N466), .O(N508) );
nor2 gate155( .a(N481), .b(N482), .O(N509) );
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );

  xor2  gate1084(.a(N492), .b(N130), .O(gate164inter0));
  nand2 gate1085(.a(gate164inter0), .b(s_100), .O(gate164inter1));
  and2  gate1086(.a(N492), .b(N130), .O(gate164inter2));
  inv1  gate1087(.a(s_100), .O(gate164inter3));
  inv1  gate1088(.a(s_101), .O(gate164inter4));
  nand2 gate1089(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1090(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1091(.a(N130), .O(gate164inter7));
  inv1  gate1092(.a(N492), .O(gate164inter8));
  nand2 gate1093(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1094(.a(s_101), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1095(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1096(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1097(.a(gate164inter12), .b(gate164inter1), .O(N518));
or2 gate165( .a(N130), .b(N492), .O(N519) );

  xor2  gate566(.a(N207), .b(N495), .O(gate166inter0));
  nand2 gate567(.a(gate166inter0), .b(s_26), .O(gate166inter1));
  and2  gate568(.a(N207), .b(N495), .O(gate166inter2));
  inv1  gate569(.a(s_26), .O(gate166inter3));
  inv1  gate570(.a(s_27), .O(gate166inter4));
  nand2 gate571(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate572(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate573(.a(N495), .O(gate166inter7));
  inv1  gate574(.a(N207), .O(gate166inter8));
  nand2 gate575(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate576(.a(s_27), .b(gate166inter3), .O(gate166inter10));
  nor2  gate577(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate578(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate579(.a(gate166inter12), .b(gate166inter1), .O(N520));
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
and2 gate170( .a(N451), .b(N171), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );
nand2 gate173( .a(N451), .b(N189), .O(N527) );

  xor2  gate1000(.a(N195), .b(N451), .O(gate174inter0));
  nand2 gate1001(.a(gate174inter0), .b(s_88), .O(gate174inter1));
  and2  gate1002(.a(N195), .b(N451), .O(gate174inter2));
  inv1  gate1003(.a(s_88), .O(gate174inter3));
  inv1  gate1004(.a(s_89), .O(gate174inter4));
  nand2 gate1005(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1006(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1007(.a(N451), .O(gate174inter7));
  inv1  gate1008(.a(N195), .O(gate174inter8));
  nand2 gate1009(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1010(.a(s_89), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1011(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1012(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1013(.a(gate174inter12), .b(gate174inter1), .O(N528));
nand2 gate175( .a(N451), .b(N201), .O(N529) );
nand2 gate176( .a(N498), .b(N499), .O(N530) );
nand2 gate177( .a(N500), .b(N501), .O(N533) );
nor2 gate178( .a(N309), .b(N502), .O(N536) );

  xor2  gate734(.a(N504), .b(N316), .O(gate179inter0));
  nand2 gate735(.a(gate179inter0), .b(s_50), .O(gate179inter1));
  and2  gate736(.a(N504), .b(N316), .O(gate179inter2));
  inv1  gate737(.a(s_50), .O(gate179inter3));
  inv1  gate738(.a(s_51), .O(gate179inter4));
  nand2 gate739(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate740(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate741(.a(N316), .O(gate179inter7));
  inv1  gate742(.a(N504), .O(gate179inter8));
  nand2 gate743(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate744(.a(s_51), .b(gate179inter3), .O(gate179inter10));
  nor2  gate745(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate746(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate747(.a(gate179inter12), .b(gate179inter1), .O(N537));
nor2 gate180( .a(N317), .b(N506), .O(N538) );

  xor2  gate1056(.a(N508), .b(N318), .O(gate181inter0));
  nand2 gate1057(.a(gate181inter0), .b(s_96), .O(gate181inter1));
  and2  gate1058(.a(N508), .b(N318), .O(gate181inter2));
  inv1  gate1059(.a(s_96), .O(gate181inter3));
  inv1  gate1060(.a(s_97), .O(gate181inter4));
  nand2 gate1061(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1062(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1063(.a(N318), .O(gate181inter7));
  inv1  gate1064(.a(N508), .O(gate181inter8));
  nand2 gate1065(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1066(.a(s_97), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1067(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1068(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1069(.a(gate181inter12), .b(gate181inter1), .O(N539));
nor2 gate182( .a(N510), .b(N511), .O(N540) );
nor2 gate183( .a(N512), .b(N513), .O(N541) );
nor2 gate184( .a(N514), .b(N515), .O(N542) );

  xor2  gate986(.a(N517), .b(N516), .O(gate185inter0));
  nand2 gate987(.a(gate185inter0), .b(s_86), .O(gate185inter1));
  and2  gate988(.a(N517), .b(N516), .O(gate185inter2));
  inv1  gate989(.a(s_86), .O(gate185inter3));
  inv1  gate990(.a(s_87), .O(gate185inter4));
  nand2 gate991(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate992(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate993(.a(N516), .O(gate185inter7));
  inv1  gate994(.a(N517), .O(gate185inter8));
  nand2 gate995(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate996(.a(s_87), .b(gate185inter3), .O(gate185inter10));
  nor2  gate997(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate998(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate999(.a(gate185inter12), .b(gate185inter1), .O(N543));

  xor2  gate1154(.a(N519), .b(N518), .O(gate186inter0));
  nand2 gate1155(.a(gate186inter0), .b(s_110), .O(gate186inter1));
  and2  gate1156(.a(N519), .b(N518), .O(gate186inter2));
  inv1  gate1157(.a(s_110), .O(gate186inter3));
  inv1  gate1158(.a(s_111), .O(gate186inter4));
  nand2 gate1159(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1160(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1161(.a(N518), .O(gate186inter7));
  inv1  gate1162(.a(N519), .O(gate186inter8));
  nand2 gate1163(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1164(.a(s_111), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1165(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1166(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1167(.a(gate186inter12), .b(gate186inter1), .O(N544));
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );

  xor2  gate1112(.a(N503), .b(N536), .O(gate191inter0));
  nand2 gate1113(.a(gate191inter0), .b(s_104), .O(gate191inter1));
  and2  gate1114(.a(N503), .b(N536), .O(gate191inter2));
  inv1  gate1115(.a(s_104), .O(gate191inter3));
  inv1  gate1116(.a(s_105), .O(gate191inter4));
  nand2 gate1117(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1118(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1119(.a(N536), .O(gate191inter7));
  inv1  gate1120(.a(N503), .O(gate191inter8));
  nand2 gate1121(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1122(.a(s_105), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1123(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1124(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1125(.a(gate191inter12), .b(gate191inter1), .O(N553));

  xor2  gate636(.a(N505), .b(N537), .O(gate192inter0));
  nand2 gate637(.a(gate192inter0), .b(s_36), .O(gate192inter1));
  and2  gate638(.a(N505), .b(N537), .O(gate192inter2));
  inv1  gate639(.a(s_36), .O(gate192inter3));
  inv1  gate640(.a(s_37), .O(gate192inter4));
  nand2 gate641(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate642(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate643(.a(N537), .O(gate192inter7));
  inv1  gate644(.a(N505), .O(gate192inter8));
  nand2 gate645(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate646(.a(s_37), .b(gate192inter3), .O(gate192inter10));
  nor2  gate647(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate648(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate649(.a(gate192inter12), .b(gate192inter1), .O(N557));
nand2 gate193( .a(N538), .b(N507), .O(N561) );
nand2 gate194( .a(N539), .b(N509), .O(N565) );
nand2 gate195( .a(N488), .b(N540), .O(N569) );

  xor2  gate1042(.a(N541), .b(N489), .O(gate196inter0));
  nand2 gate1043(.a(gate196inter0), .b(s_94), .O(gate196inter1));
  and2  gate1044(.a(N541), .b(N489), .O(gate196inter2));
  inv1  gate1045(.a(s_94), .O(gate196inter3));
  inv1  gate1046(.a(s_95), .O(gate196inter4));
  nand2 gate1047(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1048(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1049(.a(N489), .O(gate196inter7));
  inv1  gate1050(.a(N541), .O(gate196inter8));
  nand2 gate1051(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1052(.a(s_95), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1053(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1054(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1055(.a(gate196inter12), .b(gate196inter1), .O(N573));
nand2 gate197( .a(N490), .b(N542), .O(N577) );

  xor2  gate468(.a(N543), .b(N491), .O(gate198inter0));
  nand2 gate469(.a(gate198inter0), .b(s_12), .O(gate198inter1));
  and2  gate470(.a(N543), .b(N491), .O(gate198inter2));
  inv1  gate471(.a(s_12), .O(gate198inter3));
  inv1  gate472(.a(s_13), .O(gate198inter4));
  nand2 gate473(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate474(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate475(.a(N491), .O(gate198inter7));
  inv1  gate476(.a(N543), .O(gate198inter8));
  nand2 gate477(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate478(.a(s_13), .b(gate198inter3), .O(gate198inter10));
  nor2  gate479(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate480(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate481(.a(gate198inter12), .b(gate198inter1), .O(N581));
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );

  xor2  gate706(.a(N159), .b(N553), .O(gate204inter0));
  nand2 gate707(.a(gate204inter0), .b(s_46), .O(gate204inter1));
  and2  gate708(.a(N159), .b(N553), .O(gate204inter2));
  inv1  gate709(.a(s_46), .O(gate204inter3));
  inv1  gate710(.a(s_47), .O(gate204inter4));
  nand2 gate711(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate712(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate713(.a(N553), .O(gate204inter7));
  inv1  gate714(.a(N159), .O(gate204inter8));
  nand2 gate715(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate716(.a(s_47), .b(gate204inter3), .O(gate204inter10));
  nor2  gate717(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate718(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate719(.a(gate204inter12), .b(gate204inter1), .O(N590));
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );
nand2 gate207( .a(N557), .b(N165), .O(N597) );
or2 gate208( .a(N557), .b(N165), .O(N600) );
and2 gate209( .a(N246), .b(N557), .O(N605) );

  xor2  gate748(.a(N171), .b(N561), .O(gate210inter0));
  nand2 gate749(.a(gate210inter0), .b(s_52), .O(gate210inter1));
  and2  gate750(.a(N171), .b(N561), .O(gate210inter2));
  inv1  gate751(.a(s_52), .O(gate210inter3));
  inv1  gate752(.a(s_53), .O(gate210inter4));
  nand2 gate753(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate754(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate755(.a(N561), .O(gate210inter7));
  inv1  gate756(.a(N171), .O(gate210inter8));
  nand2 gate757(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate758(.a(s_53), .b(gate210inter3), .O(gate210inter10));
  nor2  gate759(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate760(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate761(.a(gate210inter12), .b(gate210inter1), .O(N606));
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );
nand2 gate213( .a(N565), .b(N177), .O(N616) );
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );

  xor2  gate1098(.a(N183), .b(N569), .O(gate216inter0));
  nand2 gate1099(.a(gate216inter0), .b(s_102), .O(gate216inter1));
  and2  gate1100(.a(N183), .b(N569), .O(gate216inter2));
  inv1  gate1101(.a(s_102), .O(gate216inter3));
  inv1  gate1102(.a(s_103), .O(gate216inter4));
  nand2 gate1103(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1104(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1105(.a(N569), .O(gate216inter7));
  inv1  gate1106(.a(N183), .O(gate216inter8));
  nand2 gate1107(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1108(.a(s_103), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1109(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1110(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1111(.a(gate216inter12), .b(gate216inter1), .O(N625));
or2 gate217( .a(N569), .b(N183), .O(N628) );
and2 gate218( .a(N246), .b(N569), .O(N631) );

  xor2  gate958(.a(N189), .b(N573), .O(gate219inter0));
  nand2 gate959(.a(gate219inter0), .b(s_82), .O(gate219inter1));
  and2  gate960(.a(N189), .b(N573), .O(gate219inter2));
  inv1  gate961(.a(s_82), .O(gate219inter3));
  inv1  gate962(.a(s_83), .O(gate219inter4));
  nand2 gate963(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate964(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate965(.a(N573), .O(gate219inter7));
  inv1  gate966(.a(N189), .O(gate219inter8));
  nand2 gate967(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate968(.a(s_83), .b(gate219inter3), .O(gate219inter10));
  nor2  gate969(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate970(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate971(.a(gate219inter12), .b(gate219inter1), .O(N632));
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );

  xor2  gate510(.a(N195), .b(N577), .O(gate222inter0));
  nand2 gate511(.a(gate222inter0), .b(s_18), .O(gate222inter1));
  and2  gate512(.a(N195), .b(N577), .O(gate222inter2));
  inv1  gate513(.a(s_18), .O(gate222inter3));
  inv1  gate514(.a(s_19), .O(gate222inter4));
  nand2 gate515(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate516(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate517(.a(N577), .O(gate222inter7));
  inv1  gate518(.a(N195), .O(gate222inter8));
  nand2 gate519(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate520(.a(s_19), .b(gate222inter3), .O(gate222inter10));
  nor2  gate521(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate522(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate523(.a(gate222inter12), .b(gate222inter1), .O(N641));
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );
nand2 gate225( .a(N581), .b(N201), .O(N651) );
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );
nor2 gate228( .a(N552), .b(N588), .O(N660) );

  xor2  gate454(.a(N589), .b(N587), .O(gate229inter0));
  nand2 gate455(.a(gate229inter0), .b(s_10), .O(gate229inter1));
  and2  gate456(.a(N589), .b(N587), .O(gate229inter2));
  inv1  gate457(.a(s_10), .O(gate229inter3));
  inv1  gate458(.a(s_11), .O(gate229inter4));
  nand2 gate459(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate460(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate461(.a(N587), .O(gate229inter7));
  inv1  gate462(.a(N589), .O(gate229inter8));
  nand2 gate463(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate464(.a(s_11), .b(gate229inter3), .O(gate229inter10));
  nor2  gate465(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate466(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate467(.a(gate229inter12), .b(gate229inter1), .O(N661));
inv1 gate230( .a(N590), .O(N662) );
and2 gate231( .a(N593), .b(N590), .O(N665) );
nor2 gate232( .a(N596), .b(N522), .O(N669) );
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );

  xor2  gate1126(.a(N523), .b(N605), .O(gate235inter0));
  nand2 gate1127(.a(gate235inter0), .b(s_106), .O(gate235inter1));
  and2  gate1128(.a(N523), .b(N605), .O(gate235inter2));
  inv1  gate1129(.a(s_106), .O(gate235inter3));
  inv1  gate1130(.a(s_107), .O(gate235inter4));
  nand2 gate1131(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1132(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1133(.a(N605), .O(gate235inter7));
  inv1  gate1134(.a(N523), .O(gate235inter8));
  nand2 gate1135(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1136(.a(s_107), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1137(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1138(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1139(.a(gate235inter12), .b(gate235inter1), .O(N677));
inv1 gate236( .a(N606), .O(N678) );
and2 gate237( .a(N609), .b(N606), .O(N682) );
nor2 gate238( .a(N615), .b(N524), .O(N686) );
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );

  xor2  gate650(.a(N525), .b(N624), .O(gate241inter0));
  nand2 gate651(.a(gate241inter0), .b(s_38), .O(gate241inter1));
  and2  gate652(.a(N525), .b(N624), .O(gate241inter2));
  inv1  gate653(.a(s_38), .O(gate241inter3));
  inv1  gate654(.a(s_39), .O(gate241inter4));
  nand2 gate655(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate656(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate657(.a(N624), .O(gate241inter7));
  inv1  gate658(.a(N525), .O(gate241inter8));
  nand2 gate659(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate660(.a(s_39), .b(gate241inter3), .O(gate241inter10));
  nor2  gate661(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate662(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate663(.a(gate241inter12), .b(gate241inter1), .O(N696));
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );
nor2 gate244( .a(N631), .b(N526), .O(N704) );
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );
nor2 gate247( .a(N337), .b(N640), .O(N712) );
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );
nor2 gate250( .a(N339), .b(N650), .O(N721) );
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );
nor2 gate253( .a(N341), .b(N659), .O(N731) );

  xor2  gate1028(.a(N261), .b(N654), .O(gate254inter0));
  nand2 gate1029(.a(gate254inter0), .b(s_92), .O(gate254inter1));
  and2  gate1030(.a(N261), .b(N654), .O(gate254inter2));
  inv1  gate1031(.a(s_92), .O(gate254inter3));
  inv1  gate1032(.a(s_93), .O(gate254inter4));
  nand2 gate1033(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1034(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1035(.a(N654), .O(gate254inter7));
  inv1  gate1036(.a(N261), .O(gate254inter8));
  nand2 gate1037(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1038(.a(s_93), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1039(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1040(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1041(.a(gate254inter12), .b(gate254inter1), .O(N732));
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
and2 gate273( .a(N228), .b(N708), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );

  xor2  gate930(.a(N261), .b(N727), .O(gate279inter0));
  nand2 gate931(.a(gate279inter0), .b(s_78), .O(gate279inter1));
  and2  gate932(.a(N261), .b(N727), .O(gate279inter2));
  inv1  gate933(.a(s_78), .O(gate279inter3));
  inv1  gate934(.a(s_79), .O(gate279inter4));
  nand2 gate935(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate936(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate937(.a(N727), .O(gate279inter7));
  inv1  gate938(.a(N261), .O(gate279inter8));
  nand2 gate939(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate940(.a(s_79), .b(gate279inter3), .O(gate279inter10));
  nor2  gate941(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate942(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate943(.a(gate279inter12), .b(gate279inter1), .O(N757));
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );
nand2 gate284( .a(N635), .b(N713), .O(N762) );
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );

  xor2  gate972(.a(N737), .b(N736), .O(gate291inter0));
  nand2 gate973(.a(gate291inter0), .b(s_84), .O(gate291inter1));
  and2  gate974(.a(N737), .b(N736), .O(gate291inter2));
  inv1  gate975(.a(s_84), .O(gate291inter3));
  inv1  gate976(.a(s_85), .O(gate291inter4));
  nand2 gate977(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate978(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate979(.a(N736), .O(gate291inter7));
  inv1  gate980(.a(N737), .O(gate291inter8));
  nand2 gate981(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate982(.a(s_85), .b(gate291inter3), .O(gate291inter10));
  nor2  gate983(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate984(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate985(.a(gate291inter12), .b(gate291inter1), .O(N769));
nor2 gate292( .a(N739), .b(N740), .O(N770) );

  xor2  gate622(.a(N743), .b(N742), .O(gate293inter0));
  nand2 gate623(.a(gate293inter0), .b(s_34), .O(gate293inter1));
  and2  gate624(.a(N743), .b(N742), .O(gate293inter2));
  inv1  gate625(.a(s_34), .O(gate293inter3));
  inv1  gate626(.a(s_35), .O(gate293inter4));
  nand2 gate627(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate628(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate629(.a(N742), .O(gate293inter7));
  inv1  gate630(.a(N743), .O(gate293inter8));
  nand2 gate631(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate632(.a(s_35), .b(gate293inter3), .O(gate293inter10));
  nor2  gate633(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate634(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate635(.a(gate293inter12), .b(gate293inter1), .O(N771));

  xor2  gate720(.a(N746), .b(N745), .O(gate294inter0));
  nand2 gate721(.a(gate294inter0), .b(s_48), .O(gate294inter1));
  and2  gate722(.a(N746), .b(N745), .O(gate294inter2));
  inv1  gate723(.a(s_48), .O(gate294inter3));
  inv1  gate724(.a(s_49), .O(gate294inter4));
  nand2 gate725(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate726(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate727(.a(N745), .O(gate294inter7));
  inv1  gate728(.a(N746), .O(gate294inter8));
  nand2 gate729(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate730(.a(s_49), .b(gate294inter3), .O(gate294inter10));
  nor2  gate731(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate732(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate733(.a(gate294inter12), .b(gate294inter1), .O(N772));
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );
nor2 gate296( .a(N748), .b(N749), .O(N777) );
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );

  xor2  gate384(.a(N752), .b(N751), .O(gate298inter0));
  nand2 gate385(.a(gate298inter0), .b(s_0), .O(gate298inter1));
  and2  gate386(.a(N752), .b(N751), .O(gate298inter2));
  inv1  gate387(.a(s_0), .O(gate298inter3));
  inv1  gate388(.a(s_1), .O(gate298inter4));
  nand2 gate389(.a(gate298inter4), .b(gate298inter3), .O(gate298inter5));
  nor2  gate390(.a(gate298inter5), .b(gate298inter2), .O(gate298inter6));
  inv1  gate391(.a(N751), .O(gate298inter7));
  inv1  gate392(.a(N752), .O(gate298inter8));
  nand2 gate393(.a(gate298inter8), .b(gate298inter7), .O(gate298inter9));
  nand2 gate394(.a(s_1), .b(gate298inter3), .O(gate298inter10));
  nor2  gate395(.a(gate298inter10), .b(gate298inter9), .O(gate298inter11));
  nor2  gate396(.a(gate298inter11), .b(gate298inter6), .O(gate298inter12));
  nand2 gate397(.a(gate298inter12), .b(gate298inter1), .O(N781));

  xor2  gate412(.a(N732), .b(N756), .O(gate299inter0));
  nand2 gate413(.a(gate299inter0), .b(s_4), .O(gate299inter1));
  and2  gate414(.a(N732), .b(N756), .O(gate299inter2));
  inv1  gate415(.a(s_4), .O(gate299inter3));
  inv1  gate416(.a(s_5), .O(gate299inter4));
  nand2 gate417(.a(gate299inter4), .b(gate299inter3), .O(gate299inter5));
  nor2  gate418(.a(gate299inter5), .b(gate299inter2), .O(gate299inter6));
  inv1  gate419(.a(N756), .O(gate299inter7));
  inv1  gate420(.a(N732), .O(gate299inter8));
  nand2 gate421(.a(gate299inter8), .b(gate299inter7), .O(gate299inter9));
  nand2 gate422(.a(s_5), .b(gate299inter3), .O(gate299inter10));
  nor2  gate423(.a(gate299inter10), .b(gate299inter9), .O(gate299inter11));
  nor2  gate424(.a(gate299inter11), .b(gate299inter6), .O(gate299inter12));
  nand2 gate425(.a(gate299inter12), .b(gate299inter1), .O(N782));

  xor2  gate902(.a(N755), .b(N754), .O(gate300inter0));
  nand2 gate903(.a(gate300inter0), .b(s_74), .O(gate300inter1));
  and2  gate904(.a(N755), .b(N754), .O(gate300inter2));
  inv1  gate905(.a(s_74), .O(gate300inter3));
  inv1  gate906(.a(s_75), .O(gate300inter4));
  nand2 gate907(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate908(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate909(.a(N754), .O(gate300inter7));
  inv1  gate910(.a(N755), .O(gate300inter8));
  nand2 gate911(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate912(.a(s_75), .b(gate300inter3), .O(gate300inter10));
  nor2  gate913(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate914(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate915(.a(gate300inter12), .b(gate300inter1), .O(N785));
nor2 gate301( .a(N757), .b(N758), .O(N786) );
nor2 gate302( .a(N759), .b(N760), .O(N787) );
nor2 gate303( .a(N700), .b(N773), .O(N788) );
and2 gate304( .a(N700), .b(N773), .O(N789) );

  xor2  gate440(.a(N778), .b(N708), .O(gate305inter0));
  nand2 gate441(.a(gate305inter0), .b(s_8), .O(gate305inter1));
  and2  gate442(.a(N778), .b(N708), .O(gate305inter2));
  inv1  gate443(.a(s_8), .O(gate305inter3));
  inv1  gate444(.a(s_9), .O(gate305inter4));
  nand2 gate445(.a(gate305inter4), .b(gate305inter3), .O(gate305inter5));
  nor2  gate446(.a(gate305inter5), .b(gate305inter2), .O(gate305inter6));
  inv1  gate447(.a(N708), .O(gate305inter7));
  inv1  gate448(.a(N778), .O(gate305inter8));
  nand2 gate449(.a(gate305inter8), .b(gate305inter7), .O(gate305inter9));
  nand2 gate450(.a(s_9), .b(gate305inter3), .O(gate305inter10));
  nor2  gate451(.a(gate305inter10), .b(gate305inter9), .O(gate305inter11));
  nor2  gate452(.a(gate305inter11), .b(gate305inter6), .O(gate305inter12));
  nand2 gate453(.a(gate305inter12), .b(gate305inter1), .O(N790));
and2 gate306( .a(N708), .b(N778), .O(N791) );
nor2 gate307( .a(N717), .b(N782), .O(N792) );
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );
nand2 gate310( .a(N628), .b(N773), .O(N795) );
nand2 gate311( .a(N795), .b(N747), .O(N796) );

  xor2  gate762(.a(N789), .b(N788), .O(gate312inter0));
  nand2 gate763(.a(gate312inter0), .b(s_54), .O(gate312inter1));
  and2  gate764(.a(N789), .b(N788), .O(gate312inter2));
  inv1  gate765(.a(s_54), .O(gate312inter3));
  inv1  gate766(.a(s_55), .O(gate312inter4));
  nand2 gate767(.a(gate312inter4), .b(gate312inter3), .O(gate312inter5));
  nor2  gate768(.a(gate312inter5), .b(gate312inter2), .O(gate312inter6));
  inv1  gate769(.a(N788), .O(gate312inter7));
  inv1  gate770(.a(N789), .O(gate312inter8));
  nand2 gate771(.a(gate312inter8), .b(gate312inter7), .O(gate312inter9));
  nand2 gate772(.a(s_55), .b(gate312inter3), .O(gate312inter10));
  nor2  gate773(.a(gate312inter10), .b(gate312inter9), .O(gate312inter11));
  nor2  gate774(.a(gate312inter11), .b(gate312inter6), .O(gate312inter12));
  nand2 gate775(.a(gate312inter12), .b(gate312inter1), .O(N802));

  xor2  gate832(.a(N791), .b(N790), .O(gate313inter0));
  nand2 gate833(.a(gate313inter0), .b(s_64), .O(gate313inter1));
  and2  gate834(.a(N791), .b(N790), .O(gate313inter2));
  inv1  gate835(.a(s_64), .O(gate313inter3));
  inv1  gate836(.a(s_65), .O(gate313inter4));
  nand2 gate837(.a(gate313inter4), .b(gate313inter3), .O(gate313inter5));
  nor2  gate838(.a(gate313inter5), .b(gate313inter2), .O(gate313inter6));
  inv1  gate839(.a(N790), .O(gate313inter7));
  inv1  gate840(.a(N791), .O(gate313inter8));
  nand2 gate841(.a(gate313inter8), .b(gate313inter7), .O(gate313inter9));
  nand2 gate842(.a(s_65), .b(gate313inter3), .O(gate313inter10));
  nor2  gate843(.a(gate313inter10), .b(gate313inter9), .O(gate313inter11));
  nor2  gate844(.a(gate313inter11), .b(gate313inter6), .O(gate313inter12));
  nand2 gate845(.a(gate313inter12), .b(gate313inter1), .O(N803));

  xor2  gate580(.a(N793), .b(N792), .O(gate314inter0));
  nand2 gate581(.a(gate314inter0), .b(s_28), .O(gate314inter1));
  and2  gate582(.a(N793), .b(N792), .O(gate314inter2));
  inv1  gate583(.a(s_28), .O(gate314inter3));
  inv1  gate584(.a(s_29), .O(gate314inter4));
  nand2 gate585(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate586(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate587(.a(N792), .O(gate314inter7));
  inv1  gate588(.a(N793), .O(gate314inter8));
  nand2 gate589(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate590(.a(s_29), .b(gate314inter3), .O(gate314inter10));
  nor2  gate591(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate592(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate593(.a(gate314inter12), .b(gate314inter1), .O(N804));
nor2 gate315( .a(N340), .b(N794), .O(N805) );

  xor2  gate482(.a(N796), .b(N692), .O(gate316inter0));
  nand2 gate483(.a(gate316inter0), .b(s_14), .O(gate316inter1));
  and2  gate484(.a(N796), .b(N692), .O(gate316inter2));
  inv1  gate485(.a(s_14), .O(gate316inter3));
  inv1  gate486(.a(s_15), .O(gate316inter4));
  nand2 gate487(.a(gate316inter4), .b(gate316inter3), .O(gate316inter5));
  nor2  gate488(.a(gate316inter5), .b(gate316inter2), .O(gate316inter6));
  inv1  gate489(.a(N692), .O(gate316inter7));
  inv1  gate490(.a(N796), .O(gate316inter8));
  nand2 gate491(.a(gate316inter8), .b(gate316inter7), .O(gate316inter9));
  nand2 gate492(.a(s_15), .b(gate316inter3), .O(gate316inter10));
  nor2  gate493(.a(gate316inter10), .b(gate316inter9), .O(gate316inter11));
  nor2  gate494(.a(gate316inter11), .b(gate316inter6), .O(gate316inter12));
  nand2 gate495(.a(gate316inter12), .b(gate316inter1), .O(N806));
and2 gate317( .a(N692), .b(N796), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );

  xor2  gate678(.a(N796), .b(N619), .O(gate322inter0));
  nand2 gate679(.a(gate322inter0), .b(s_42), .O(gate322inter1));
  and2  gate680(.a(N796), .b(N619), .O(gate322inter2));
  inv1  gate681(.a(s_42), .O(gate322inter3));
  inv1  gate682(.a(s_43), .O(gate322inter4));
  nand2 gate683(.a(gate322inter4), .b(gate322inter3), .O(gate322inter5));
  nor2  gate684(.a(gate322inter5), .b(gate322inter2), .O(gate322inter6));
  inv1  gate685(.a(N619), .O(gate322inter7));
  inv1  gate686(.a(N796), .O(gate322inter8));
  nand2 gate687(.a(gate322inter8), .b(gate322inter7), .O(gate322inter9));
  nand2 gate688(.a(s_43), .b(gate322inter3), .O(gate322inter10));
  nor2  gate689(.a(gate322inter10), .b(gate322inter9), .O(gate322inter11));
  nor2  gate690(.a(gate322inter11), .b(gate322inter6), .O(gate322inter12));
  nand2 gate691(.a(gate322inter12), .b(gate322inter1), .O(N812));
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );
nand2 gate327( .a(N744), .b(N812), .O(N822) );
nor2 gate328( .a(N806), .b(N807), .O(N825) );
nor2 gate329( .a(N335), .b(N808), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );

  xor2  gate664(.a(N815), .b(N665), .O(gate333inter0));
  nand2 gate665(.a(gate333inter0), .b(s_40), .O(gate333inter1));
  and2  gate666(.a(N815), .b(N665), .O(gate333inter2));
  inv1  gate667(.a(s_40), .O(gate333inter3));
  inv1  gate668(.a(s_41), .O(gate333inter4));
  nand2 gate669(.a(gate333inter4), .b(gate333inter3), .O(gate333inter5));
  nor2  gate670(.a(gate333inter5), .b(gate333inter2), .O(gate333inter6));
  inv1  gate671(.a(N665), .O(gate333inter7));
  inv1  gate672(.a(N815), .O(gate333inter8));
  nand2 gate673(.a(gate333inter8), .b(gate333inter7), .O(gate333inter9));
  nand2 gate674(.a(s_41), .b(gate333inter3), .O(gate333inter10));
  nor2  gate675(.a(gate333inter10), .b(gate333inter9), .O(gate333inter11));
  nor2  gate676(.a(gate333inter11), .b(gate333inter6), .O(gate333inter12));
  nand2 gate677(.a(gate333inter12), .b(gate333inter1), .O(N830));
and2 gate334( .a(N665), .b(N815), .O(N831) );

  xor2  gate594(.a(N819), .b(N673), .O(gate335inter0));
  nand2 gate595(.a(gate335inter0), .b(s_30), .O(gate335inter1));
  and2  gate596(.a(N819), .b(N673), .O(gate335inter2));
  inv1  gate597(.a(s_30), .O(gate335inter3));
  inv1  gate598(.a(s_31), .O(gate335inter4));
  nand2 gate599(.a(gate335inter4), .b(gate335inter3), .O(gate335inter5));
  nor2  gate600(.a(gate335inter5), .b(gate335inter2), .O(gate335inter6));
  inv1  gate601(.a(N673), .O(gate335inter7));
  inv1  gate602(.a(N819), .O(gate335inter8));
  nand2 gate603(.a(gate335inter8), .b(gate335inter7), .O(gate335inter9));
  nand2 gate604(.a(s_31), .b(gate335inter3), .O(gate335inter10));
  nor2  gate605(.a(gate335inter10), .b(gate335inter9), .O(gate335inter11));
  nor2  gate606(.a(gate335inter11), .b(gate335inter6), .O(gate335inter12));
  nand2 gate607(.a(gate335inter12), .b(gate335inter1), .O(N832));
and2 gate336( .a(N673), .b(N819), .O(N833) );
nor2 gate337( .a(N682), .b(N822), .O(N834) );
and2 gate338( .a(N682), .b(N822), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
nand2 gate344( .a(N815), .b(N593), .O(N841) );
nor2 gate345( .a(N830), .b(N831), .O(N842) );
nor2 gate346( .a(N832), .b(N833), .O(N843) );
nor2 gate347( .a(N834), .b(N835), .O(N844) );
nor2 gate348( .a(N334), .b(N836), .O(N845) );
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
and2 gate354( .a(N219), .b(N842), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );

  xor2  gate1140(.a(N851), .b(N417), .O(gate362inter0));
  nand2 gate1141(.a(gate362inter0), .b(s_108), .O(gate362inter1));
  and2  gate1142(.a(N851), .b(N417), .O(gate362inter2));
  inv1  gate1143(.a(s_108), .O(gate362inter3));
  inv1  gate1144(.a(s_109), .O(gate362inter4));
  nand2 gate1145(.a(gate362inter4), .b(gate362inter3), .O(gate362inter5));
  nor2  gate1146(.a(gate362inter5), .b(gate362inter2), .O(gate362inter6));
  inv1  gate1147(.a(N417), .O(gate362inter7));
  inv1  gate1148(.a(N851), .O(gate362inter8));
  nand2 gate1149(.a(gate362inter8), .b(gate362inter7), .O(gate362inter9));
  nand2 gate1150(.a(s_109), .b(gate362inter3), .O(gate362inter10));
  nor2  gate1151(.a(gate362inter10), .b(gate362inter9), .O(gate362inter11));
  nor2  gate1152(.a(gate362inter11), .b(gate362inter6), .O(gate362inter12));
  nand2 gate1153(.a(gate362inter12), .b(gate362inter1), .O(N859));

  xor2  gate608(.a(N852), .b(N332), .O(gate363inter0));
  nand2 gate609(.a(gate363inter0), .b(s_32), .O(gate363inter1));
  and2  gate610(.a(N852), .b(N332), .O(gate363inter2));
  inv1  gate611(.a(s_32), .O(gate363inter3));
  inv1  gate612(.a(s_33), .O(gate363inter4));
  nand2 gate613(.a(gate363inter4), .b(gate363inter3), .O(gate363inter5));
  nor2  gate614(.a(gate363inter5), .b(gate363inter2), .O(gate363inter6));
  inv1  gate615(.a(N332), .O(gate363inter7));
  inv1  gate616(.a(N852), .O(gate363inter8));
  nand2 gate617(.a(gate363inter8), .b(gate363inter7), .O(gate363inter9));
  nand2 gate618(.a(s_33), .b(gate363inter3), .O(gate363inter10));
  nor2  gate619(.a(gate363inter10), .b(gate363inter9), .O(gate363inter11));
  nor2  gate620(.a(gate363inter11), .b(gate363inter6), .O(gate363inter12));
  nand2 gate621(.a(gate363inter12), .b(gate363inter1), .O(N860));
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

endmodule