module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381, s_382, s_383, s_384, s_385, s_386, s_387, s_388, s_389, s_390, s_391, s_392, s_393, s_394, s_395, s_396, s_397, s_398, s_399, s_400, s_401;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2297(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2298(.a(gate11inter0), .b(s_250), .O(gate11inter1));
  and2  gate2299(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2300(.a(s_250), .O(gate11inter3));
  inv1  gate2301(.a(s_251), .O(gate11inter4));
  nand2 gate2302(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2303(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2304(.a(G5), .O(gate11inter7));
  inv1  gate2305(.a(G6), .O(gate11inter8));
  nand2 gate2306(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2307(.a(s_251), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2308(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2309(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2310(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1709(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1710(.a(gate12inter0), .b(s_166), .O(gate12inter1));
  and2  gate1711(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1712(.a(s_166), .O(gate12inter3));
  inv1  gate1713(.a(s_167), .O(gate12inter4));
  nand2 gate1714(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1715(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1716(.a(G7), .O(gate12inter7));
  inv1  gate1717(.a(G8), .O(gate12inter8));
  nand2 gate1718(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1719(.a(s_167), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1720(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1721(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1722(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2157(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2158(.a(gate14inter0), .b(s_230), .O(gate14inter1));
  and2  gate2159(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2160(.a(s_230), .O(gate14inter3));
  inv1  gate2161(.a(s_231), .O(gate14inter4));
  nand2 gate2162(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2163(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2164(.a(G11), .O(gate14inter7));
  inv1  gate2165(.a(G12), .O(gate14inter8));
  nand2 gate2166(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2167(.a(s_231), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2168(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2169(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2170(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1415(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1416(.a(gate16inter0), .b(s_124), .O(gate16inter1));
  and2  gate1417(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1418(.a(s_124), .O(gate16inter3));
  inv1  gate1419(.a(s_125), .O(gate16inter4));
  nand2 gate1420(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1421(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1422(.a(G15), .O(gate16inter7));
  inv1  gate1423(.a(G16), .O(gate16inter8));
  nand2 gate1424(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1425(.a(s_125), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1426(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1427(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1428(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate2311(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2312(.a(gate18inter0), .b(s_252), .O(gate18inter1));
  and2  gate2313(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2314(.a(s_252), .O(gate18inter3));
  inv1  gate2315(.a(s_253), .O(gate18inter4));
  nand2 gate2316(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2317(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2318(.a(G19), .O(gate18inter7));
  inv1  gate2319(.a(G20), .O(gate18inter8));
  nand2 gate2320(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2321(.a(s_253), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2322(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2323(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2324(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1373(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1374(.a(gate19inter0), .b(s_118), .O(gate19inter1));
  and2  gate1375(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1376(.a(s_118), .O(gate19inter3));
  inv1  gate1377(.a(s_119), .O(gate19inter4));
  nand2 gate1378(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1379(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1380(.a(G21), .O(gate19inter7));
  inv1  gate1381(.a(G22), .O(gate19inter8));
  nand2 gate1382(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1383(.a(s_119), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1384(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1385(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1386(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1653(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1654(.a(gate20inter0), .b(s_158), .O(gate20inter1));
  and2  gate1655(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1656(.a(s_158), .O(gate20inter3));
  inv1  gate1657(.a(s_159), .O(gate20inter4));
  nand2 gate1658(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1659(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1660(.a(G23), .O(gate20inter7));
  inv1  gate1661(.a(G24), .O(gate20inter8));
  nand2 gate1662(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1663(.a(s_159), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1664(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1665(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1666(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1919(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1920(.a(gate21inter0), .b(s_196), .O(gate21inter1));
  and2  gate1921(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1922(.a(s_196), .O(gate21inter3));
  inv1  gate1923(.a(s_197), .O(gate21inter4));
  nand2 gate1924(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1925(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1926(.a(G25), .O(gate21inter7));
  inv1  gate1927(.a(G26), .O(gate21inter8));
  nand2 gate1928(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1929(.a(s_197), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1930(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1931(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1932(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate715(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate716(.a(gate28inter0), .b(s_24), .O(gate28inter1));
  and2  gate717(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate718(.a(s_24), .O(gate28inter3));
  inv1  gate719(.a(s_25), .O(gate28inter4));
  nand2 gate720(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate721(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate722(.a(G10), .O(gate28inter7));
  inv1  gate723(.a(G14), .O(gate28inter8));
  nand2 gate724(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate725(.a(s_25), .b(gate28inter3), .O(gate28inter10));
  nor2  gate726(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate727(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate728(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate799(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate800(.a(gate29inter0), .b(s_36), .O(gate29inter1));
  and2  gate801(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate802(.a(s_36), .O(gate29inter3));
  inv1  gate803(.a(s_37), .O(gate29inter4));
  nand2 gate804(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate805(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate806(.a(G3), .O(gate29inter7));
  inv1  gate807(.a(G7), .O(gate29inter8));
  nand2 gate808(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate809(.a(s_37), .b(gate29inter3), .O(gate29inter10));
  nor2  gate810(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate811(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate812(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1471(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1472(.a(gate33inter0), .b(s_132), .O(gate33inter1));
  and2  gate1473(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1474(.a(s_132), .O(gate33inter3));
  inv1  gate1475(.a(s_133), .O(gate33inter4));
  nand2 gate1476(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1477(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1478(.a(G17), .O(gate33inter7));
  inv1  gate1479(.a(G21), .O(gate33inter8));
  nand2 gate1480(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1481(.a(s_133), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1482(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1483(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1484(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate2339(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2340(.a(gate34inter0), .b(s_256), .O(gate34inter1));
  and2  gate2341(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2342(.a(s_256), .O(gate34inter3));
  inv1  gate2343(.a(s_257), .O(gate34inter4));
  nand2 gate2344(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2345(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2346(.a(G25), .O(gate34inter7));
  inv1  gate2347(.a(G29), .O(gate34inter8));
  nand2 gate2348(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2349(.a(s_257), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2350(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2351(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2352(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate3333(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate3334(.a(gate36inter0), .b(s_398), .O(gate36inter1));
  and2  gate3335(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate3336(.a(s_398), .O(gate36inter3));
  inv1  gate3337(.a(s_399), .O(gate36inter4));
  nand2 gate3338(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate3339(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate3340(.a(G26), .O(gate36inter7));
  inv1  gate3341(.a(G30), .O(gate36inter8));
  nand2 gate3342(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate3343(.a(s_399), .b(gate36inter3), .O(gate36inter10));
  nor2  gate3344(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate3345(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate3346(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate939(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate940(.a(gate37inter0), .b(s_56), .O(gate37inter1));
  and2  gate941(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate942(.a(s_56), .O(gate37inter3));
  inv1  gate943(.a(s_57), .O(gate37inter4));
  nand2 gate944(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate945(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate946(.a(G19), .O(gate37inter7));
  inv1  gate947(.a(G23), .O(gate37inter8));
  nand2 gate948(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate949(.a(s_57), .b(gate37inter3), .O(gate37inter10));
  nor2  gate950(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate951(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate952(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate3095(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate3096(.a(gate38inter0), .b(s_364), .O(gate38inter1));
  and2  gate3097(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate3098(.a(s_364), .O(gate38inter3));
  inv1  gate3099(.a(s_365), .O(gate38inter4));
  nand2 gate3100(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate3101(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate3102(.a(G27), .O(gate38inter7));
  inv1  gate3103(.a(G31), .O(gate38inter8));
  nand2 gate3104(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate3105(.a(s_365), .b(gate38inter3), .O(gate38inter10));
  nor2  gate3106(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate3107(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate3108(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1751(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1752(.a(gate39inter0), .b(s_172), .O(gate39inter1));
  and2  gate1753(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1754(.a(s_172), .O(gate39inter3));
  inv1  gate1755(.a(s_173), .O(gate39inter4));
  nand2 gate1756(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1757(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1758(.a(G20), .O(gate39inter7));
  inv1  gate1759(.a(G24), .O(gate39inter8));
  nand2 gate1760(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1761(.a(s_173), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1762(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1763(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1764(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2857(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2858(.a(gate43inter0), .b(s_330), .O(gate43inter1));
  and2  gate2859(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2860(.a(s_330), .O(gate43inter3));
  inv1  gate2861(.a(s_331), .O(gate43inter4));
  nand2 gate2862(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2863(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2864(.a(G3), .O(gate43inter7));
  inv1  gate2865(.a(G269), .O(gate43inter8));
  nand2 gate2866(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2867(.a(s_331), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2868(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2869(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2870(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate659(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate660(.a(gate45inter0), .b(s_16), .O(gate45inter1));
  and2  gate661(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate662(.a(s_16), .O(gate45inter3));
  inv1  gate663(.a(s_17), .O(gate45inter4));
  nand2 gate664(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate665(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate666(.a(G5), .O(gate45inter7));
  inv1  gate667(.a(G272), .O(gate45inter8));
  nand2 gate668(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate669(.a(s_17), .b(gate45inter3), .O(gate45inter10));
  nor2  gate670(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate671(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate672(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1793(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1794(.a(gate46inter0), .b(s_178), .O(gate46inter1));
  and2  gate1795(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1796(.a(s_178), .O(gate46inter3));
  inv1  gate1797(.a(s_179), .O(gate46inter4));
  nand2 gate1798(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1799(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1800(.a(G6), .O(gate46inter7));
  inv1  gate1801(.a(G272), .O(gate46inter8));
  nand2 gate1802(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1803(.a(s_179), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1804(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1805(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1806(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1065(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1066(.a(gate53inter0), .b(s_74), .O(gate53inter1));
  and2  gate1067(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1068(.a(s_74), .O(gate53inter3));
  inv1  gate1069(.a(s_75), .O(gate53inter4));
  nand2 gate1070(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1071(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1072(.a(G13), .O(gate53inter7));
  inv1  gate1073(.a(G284), .O(gate53inter8));
  nand2 gate1074(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1075(.a(s_75), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1076(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1077(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1078(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate687(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate688(.a(gate55inter0), .b(s_20), .O(gate55inter1));
  and2  gate689(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate690(.a(s_20), .O(gate55inter3));
  inv1  gate691(.a(s_21), .O(gate55inter4));
  nand2 gate692(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate693(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate694(.a(G15), .O(gate55inter7));
  inv1  gate695(.a(G287), .O(gate55inter8));
  nand2 gate696(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate697(.a(s_21), .b(gate55inter3), .O(gate55inter10));
  nor2  gate698(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate699(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate700(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1541(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1542(.a(gate57inter0), .b(s_142), .O(gate57inter1));
  and2  gate1543(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1544(.a(s_142), .O(gate57inter3));
  inv1  gate1545(.a(s_143), .O(gate57inter4));
  nand2 gate1546(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1547(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1548(.a(G17), .O(gate57inter7));
  inv1  gate1549(.a(G290), .O(gate57inter8));
  nand2 gate1550(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1551(.a(s_143), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1552(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1553(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1554(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate2255(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2256(.a(gate58inter0), .b(s_244), .O(gate58inter1));
  and2  gate2257(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2258(.a(s_244), .O(gate58inter3));
  inv1  gate2259(.a(s_245), .O(gate58inter4));
  nand2 gate2260(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2261(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2262(.a(G18), .O(gate58inter7));
  inv1  gate2263(.a(G290), .O(gate58inter8));
  nand2 gate2264(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2265(.a(s_245), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2266(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2267(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2268(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate813(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate814(.a(gate60inter0), .b(s_38), .O(gate60inter1));
  and2  gate815(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate816(.a(s_38), .O(gate60inter3));
  inv1  gate817(.a(s_39), .O(gate60inter4));
  nand2 gate818(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate819(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate820(.a(G20), .O(gate60inter7));
  inv1  gate821(.a(G293), .O(gate60inter8));
  nand2 gate822(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate823(.a(s_39), .b(gate60inter3), .O(gate60inter10));
  nor2  gate824(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate825(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate826(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2241(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2242(.a(gate62inter0), .b(s_242), .O(gate62inter1));
  and2  gate2243(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2244(.a(s_242), .O(gate62inter3));
  inv1  gate2245(.a(s_243), .O(gate62inter4));
  nand2 gate2246(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2247(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2248(.a(G22), .O(gate62inter7));
  inv1  gate2249(.a(G296), .O(gate62inter8));
  nand2 gate2250(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2251(.a(s_243), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2252(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2253(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2254(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2073(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2074(.a(gate63inter0), .b(s_218), .O(gate63inter1));
  and2  gate2075(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2076(.a(s_218), .O(gate63inter3));
  inv1  gate2077(.a(s_219), .O(gate63inter4));
  nand2 gate2078(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2079(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2080(.a(G23), .O(gate63inter7));
  inv1  gate2081(.a(G299), .O(gate63inter8));
  nand2 gate2082(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2083(.a(s_219), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2084(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2085(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2086(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1457(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1458(.a(gate65inter0), .b(s_130), .O(gate65inter1));
  and2  gate1459(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1460(.a(s_130), .O(gate65inter3));
  inv1  gate1461(.a(s_131), .O(gate65inter4));
  nand2 gate1462(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1463(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1464(.a(G25), .O(gate65inter7));
  inv1  gate1465(.a(G302), .O(gate65inter8));
  nand2 gate1466(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1467(.a(s_131), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1468(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1469(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1470(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2171(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2172(.a(gate68inter0), .b(s_232), .O(gate68inter1));
  and2  gate2173(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2174(.a(s_232), .O(gate68inter3));
  inv1  gate2175(.a(s_233), .O(gate68inter4));
  nand2 gate2176(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2177(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2178(.a(G28), .O(gate68inter7));
  inv1  gate2179(.a(G305), .O(gate68inter8));
  nand2 gate2180(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2181(.a(s_233), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2182(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2183(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2184(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate3249(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate3250(.a(gate70inter0), .b(s_386), .O(gate70inter1));
  and2  gate3251(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate3252(.a(s_386), .O(gate70inter3));
  inv1  gate3253(.a(s_387), .O(gate70inter4));
  nand2 gate3254(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate3255(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate3256(.a(G30), .O(gate70inter7));
  inv1  gate3257(.a(G308), .O(gate70inter8));
  nand2 gate3258(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate3259(.a(s_387), .b(gate70inter3), .O(gate70inter10));
  nor2  gate3260(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate3261(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate3262(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate3025(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate3026(.a(gate72inter0), .b(s_354), .O(gate72inter1));
  and2  gate3027(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate3028(.a(s_354), .O(gate72inter3));
  inv1  gate3029(.a(s_355), .O(gate72inter4));
  nand2 gate3030(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate3031(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate3032(.a(G32), .O(gate72inter7));
  inv1  gate3033(.a(G311), .O(gate72inter8));
  nand2 gate3034(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate3035(.a(s_355), .b(gate72inter3), .O(gate72inter10));
  nor2  gate3036(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate3037(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate3038(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate2899(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate2900(.a(gate73inter0), .b(s_336), .O(gate73inter1));
  and2  gate2901(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate2902(.a(s_336), .O(gate73inter3));
  inv1  gate2903(.a(s_337), .O(gate73inter4));
  nand2 gate2904(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate2905(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate2906(.a(G1), .O(gate73inter7));
  inv1  gate2907(.a(G314), .O(gate73inter8));
  nand2 gate2908(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate2909(.a(s_337), .b(gate73inter3), .O(gate73inter10));
  nor2  gate2910(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate2911(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate2912(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate2437(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2438(.a(gate74inter0), .b(s_270), .O(gate74inter1));
  and2  gate2439(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2440(.a(s_270), .O(gate74inter3));
  inv1  gate2441(.a(s_271), .O(gate74inter4));
  nand2 gate2442(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2443(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2444(.a(G5), .O(gate74inter7));
  inv1  gate2445(.a(G314), .O(gate74inter8));
  nand2 gate2446(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2447(.a(s_271), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2448(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2449(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2450(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate729(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate730(.a(gate75inter0), .b(s_26), .O(gate75inter1));
  and2  gate731(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate732(.a(s_26), .O(gate75inter3));
  inv1  gate733(.a(s_27), .O(gate75inter4));
  nand2 gate734(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate735(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate736(.a(G9), .O(gate75inter7));
  inv1  gate737(.a(G317), .O(gate75inter8));
  nand2 gate738(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate739(.a(s_27), .b(gate75inter3), .O(gate75inter10));
  nor2  gate740(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate741(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate742(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate2283(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2284(.a(gate76inter0), .b(s_248), .O(gate76inter1));
  and2  gate2285(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2286(.a(s_248), .O(gate76inter3));
  inv1  gate2287(.a(s_249), .O(gate76inter4));
  nand2 gate2288(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2289(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2290(.a(G13), .O(gate76inter7));
  inv1  gate2291(.a(G317), .O(gate76inter8));
  nand2 gate2292(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2293(.a(s_249), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2294(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2295(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2296(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2605(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2606(.a(gate78inter0), .b(s_294), .O(gate78inter1));
  and2  gate2607(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2608(.a(s_294), .O(gate78inter3));
  inv1  gate2609(.a(s_295), .O(gate78inter4));
  nand2 gate2610(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2611(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2612(.a(G6), .O(gate78inter7));
  inv1  gate2613(.a(G320), .O(gate78inter8));
  nand2 gate2614(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2615(.a(s_295), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2616(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2617(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2618(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate1849(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1850(.a(gate79inter0), .b(s_186), .O(gate79inter1));
  and2  gate1851(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1852(.a(s_186), .O(gate79inter3));
  inv1  gate1853(.a(s_187), .O(gate79inter4));
  nand2 gate1854(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1855(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1856(.a(G10), .O(gate79inter7));
  inv1  gate1857(.a(G323), .O(gate79inter8));
  nand2 gate1858(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1859(.a(s_187), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1860(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1861(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1862(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate2591(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2592(.a(gate80inter0), .b(s_292), .O(gate80inter1));
  and2  gate2593(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2594(.a(s_292), .O(gate80inter3));
  inv1  gate2595(.a(s_293), .O(gate80inter4));
  nand2 gate2596(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2597(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2598(.a(G14), .O(gate80inter7));
  inv1  gate2599(.a(G323), .O(gate80inter8));
  nand2 gate2600(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2601(.a(s_293), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2602(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2603(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2604(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1037(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1038(.a(gate82inter0), .b(s_70), .O(gate82inter1));
  and2  gate1039(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1040(.a(s_70), .O(gate82inter3));
  inv1  gate1041(.a(s_71), .O(gate82inter4));
  nand2 gate1042(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1043(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1044(.a(G7), .O(gate82inter7));
  inv1  gate1045(.a(G326), .O(gate82inter8));
  nand2 gate1046(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1047(.a(s_71), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1048(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1049(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1050(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1821(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1822(.a(gate84inter0), .b(s_182), .O(gate84inter1));
  and2  gate1823(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1824(.a(s_182), .O(gate84inter3));
  inv1  gate1825(.a(s_183), .O(gate84inter4));
  nand2 gate1826(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1827(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1828(.a(G15), .O(gate84inter7));
  inv1  gate1829(.a(G329), .O(gate84inter8));
  nand2 gate1830(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1831(.a(s_183), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1832(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1833(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1834(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1205(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1206(.a(gate85inter0), .b(s_94), .O(gate85inter1));
  and2  gate1207(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1208(.a(s_94), .O(gate85inter3));
  inv1  gate1209(.a(s_95), .O(gate85inter4));
  nand2 gate1210(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1211(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1212(.a(G4), .O(gate85inter7));
  inv1  gate1213(.a(G332), .O(gate85inter8));
  nand2 gate1214(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1215(.a(s_95), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1216(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1217(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1218(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate3011(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate3012(.a(gate89inter0), .b(s_352), .O(gate89inter1));
  and2  gate3013(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate3014(.a(s_352), .O(gate89inter3));
  inv1  gate3015(.a(s_353), .O(gate89inter4));
  nand2 gate3016(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate3017(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate3018(.a(G17), .O(gate89inter7));
  inv1  gate3019(.a(G338), .O(gate89inter8));
  nand2 gate3020(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate3021(.a(s_353), .b(gate89inter3), .O(gate89inter10));
  nor2  gate3022(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate3023(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate3024(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate2773(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2774(.a(gate92inter0), .b(s_318), .O(gate92inter1));
  and2  gate2775(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2776(.a(s_318), .O(gate92inter3));
  inv1  gate2777(.a(s_319), .O(gate92inter4));
  nand2 gate2778(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2779(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2780(.a(G29), .O(gate92inter7));
  inv1  gate2781(.a(G341), .O(gate92inter8));
  nand2 gate2782(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2783(.a(s_319), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2784(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2785(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2786(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1611(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1612(.a(gate95inter0), .b(s_152), .O(gate95inter1));
  and2  gate1613(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1614(.a(s_152), .O(gate95inter3));
  inv1  gate1615(.a(s_153), .O(gate95inter4));
  nand2 gate1616(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1617(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1618(.a(G26), .O(gate95inter7));
  inv1  gate1619(.a(G347), .O(gate95inter8));
  nand2 gate1620(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1621(.a(s_153), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1622(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1623(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1624(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate981(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate982(.a(gate96inter0), .b(s_62), .O(gate96inter1));
  and2  gate983(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate984(.a(s_62), .O(gate96inter3));
  inv1  gate985(.a(s_63), .O(gate96inter4));
  nand2 gate986(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate987(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate988(.a(G30), .O(gate96inter7));
  inv1  gate989(.a(G347), .O(gate96inter8));
  nand2 gate990(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate991(.a(s_63), .b(gate96inter3), .O(gate96inter10));
  nor2  gate992(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate993(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate994(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate2381(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate2382(.a(gate97inter0), .b(s_262), .O(gate97inter1));
  and2  gate2383(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate2384(.a(s_262), .O(gate97inter3));
  inv1  gate2385(.a(s_263), .O(gate97inter4));
  nand2 gate2386(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate2387(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate2388(.a(G19), .O(gate97inter7));
  inv1  gate2389(.a(G350), .O(gate97inter8));
  nand2 gate2390(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate2391(.a(s_263), .b(gate97inter3), .O(gate97inter10));
  nor2  gate2392(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate2393(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate2394(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate3081(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate3082(.a(gate100inter0), .b(s_362), .O(gate100inter1));
  and2  gate3083(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate3084(.a(s_362), .O(gate100inter3));
  inv1  gate3085(.a(s_363), .O(gate100inter4));
  nand2 gate3086(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate3087(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate3088(.a(G31), .O(gate100inter7));
  inv1  gate3089(.a(G353), .O(gate100inter8));
  nand2 gate3090(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate3091(.a(s_363), .b(gate100inter3), .O(gate100inter10));
  nor2  gate3092(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate3093(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate3094(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2871(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2872(.a(gate102inter0), .b(s_332), .O(gate102inter1));
  and2  gate2873(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2874(.a(s_332), .O(gate102inter3));
  inv1  gate2875(.a(s_333), .O(gate102inter4));
  nand2 gate2876(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2877(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2878(.a(G24), .O(gate102inter7));
  inv1  gate2879(.a(G356), .O(gate102inter8));
  nand2 gate2880(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2881(.a(s_333), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2882(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2883(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2884(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1443(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1444(.a(gate103inter0), .b(s_128), .O(gate103inter1));
  and2  gate1445(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1446(.a(s_128), .O(gate103inter3));
  inv1  gate1447(.a(s_129), .O(gate103inter4));
  nand2 gate1448(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1449(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1450(.a(G28), .O(gate103inter7));
  inv1  gate1451(.a(G359), .O(gate103inter8));
  nand2 gate1452(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1453(.a(s_129), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1454(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1455(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1456(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1975(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1976(.a(gate104inter0), .b(s_204), .O(gate104inter1));
  and2  gate1977(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1978(.a(s_204), .O(gate104inter3));
  inv1  gate1979(.a(s_205), .O(gate104inter4));
  nand2 gate1980(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1981(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1982(.a(G32), .O(gate104inter7));
  inv1  gate1983(.a(G359), .O(gate104inter8));
  nand2 gate1984(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1985(.a(s_205), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1986(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1987(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1988(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate2465(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2466(.a(gate105inter0), .b(s_274), .O(gate105inter1));
  and2  gate2467(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2468(.a(s_274), .O(gate105inter3));
  inv1  gate2469(.a(s_275), .O(gate105inter4));
  nand2 gate2470(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2471(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2472(.a(G362), .O(gate105inter7));
  inv1  gate2473(.a(G363), .O(gate105inter8));
  nand2 gate2474(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2475(.a(s_275), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2476(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2477(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2478(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate3179(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate3180(.a(gate106inter0), .b(s_376), .O(gate106inter1));
  and2  gate3181(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate3182(.a(s_376), .O(gate106inter3));
  inv1  gate3183(.a(s_377), .O(gate106inter4));
  nand2 gate3184(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate3185(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate3186(.a(G364), .O(gate106inter7));
  inv1  gate3187(.a(G365), .O(gate106inter8));
  nand2 gate3188(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate3189(.a(s_377), .b(gate106inter3), .O(gate106inter10));
  nor2  gate3190(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate3191(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate3192(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate631(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate632(.a(gate108inter0), .b(s_12), .O(gate108inter1));
  and2  gate633(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate634(.a(s_12), .O(gate108inter3));
  inv1  gate635(.a(s_13), .O(gate108inter4));
  nand2 gate636(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate637(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate638(.a(G368), .O(gate108inter7));
  inv1  gate639(.a(G369), .O(gate108inter8));
  nand2 gate640(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate641(.a(s_13), .b(gate108inter3), .O(gate108inter10));
  nor2  gate642(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate643(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate644(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate2913(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2914(.a(gate109inter0), .b(s_338), .O(gate109inter1));
  and2  gate2915(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2916(.a(s_338), .O(gate109inter3));
  inv1  gate2917(.a(s_339), .O(gate109inter4));
  nand2 gate2918(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2919(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2920(.a(G370), .O(gate109inter7));
  inv1  gate2921(.a(G371), .O(gate109inter8));
  nand2 gate2922(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2923(.a(s_339), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2924(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2925(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2926(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2983(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2984(.a(gate111inter0), .b(s_348), .O(gate111inter1));
  and2  gate2985(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2986(.a(s_348), .O(gate111inter3));
  inv1  gate2987(.a(s_349), .O(gate111inter4));
  nand2 gate2988(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2989(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2990(.a(G374), .O(gate111inter7));
  inv1  gate2991(.a(G375), .O(gate111inter8));
  nand2 gate2992(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2993(.a(s_349), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2994(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2995(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2996(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate757(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate758(.a(gate115inter0), .b(s_30), .O(gate115inter1));
  and2  gate759(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate760(.a(s_30), .O(gate115inter3));
  inv1  gate761(.a(s_31), .O(gate115inter4));
  nand2 gate762(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate763(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate764(.a(G382), .O(gate115inter7));
  inv1  gate765(.a(G383), .O(gate115inter8));
  nand2 gate766(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate767(.a(s_31), .b(gate115inter3), .O(gate115inter10));
  nor2  gate768(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate769(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate770(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate561(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate562(.a(gate116inter0), .b(s_2), .O(gate116inter1));
  and2  gate563(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate564(.a(s_2), .O(gate116inter3));
  inv1  gate565(.a(s_3), .O(gate116inter4));
  nand2 gate566(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate567(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate568(.a(G384), .O(gate116inter7));
  inv1  gate569(.a(G385), .O(gate116inter8));
  nand2 gate570(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate571(.a(s_3), .b(gate116inter3), .O(gate116inter10));
  nor2  gate572(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate573(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate574(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate2969(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2970(.a(gate117inter0), .b(s_346), .O(gate117inter1));
  and2  gate2971(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2972(.a(s_346), .O(gate117inter3));
  inv1  gate2973(.a(s_347), .O(gate117inter4));
  nand2 gate2974(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2975(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2976(.a(G386), .O(gate117inter7));
  inv1  gate2977(.a(G387), .O(gate117inter8));
  nand2 gate2978(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2979(.a(s_347), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2980(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2981(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2982(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate3067(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate3068(.a(gate118inter0), .b(s_360), .O(gate118inter1));
  and2  gate3069(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate3070(.a(s_360), .O(gate118inter3));
  inv1  gate3071(.a(s_361), .O(gate118inter4));
  nand2 gate3072(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate3073(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate3074(.a(G388), .O(gate118inter7));
  inv1  gate3075(.a(G389), .O(gate118inter8));
  nand2 gate3076(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate3077(.a(s_361), .b(gate118inter3), .O(gate118inter10));
  nor2  gate3078(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate3079(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate3080(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2647(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2648(.a(gate122inter0), .b(s_300), .O(gate122inter1));
  and2  gate2649(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2650(.a(s_300), .O(gate122inter3));
  inv1  gate2651(.a(s_301), .O(gate122inter4));
  nand2 gate2652(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2653(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2654(.a(G396), .O(gate122inter7));
  inv1  gate2655(.a(G397), .O(gate122inter8));
  nand2 gate2656(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2657(.a(s_301), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2658(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2659(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2660(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1947(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1948(.a(gate125inter0), .b(s_200), .O(gate125inter1));
  and2  gate1949(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1950(.a(s_200), .O(gate125inter3));
  inv1  gate1951(.a(s_201), .O(gate125inter4));
  nand2 gate1952(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1953(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1954(.a(G402), .O(gate125inter7));
  inv1  gate1955(.a(G403), .O(gate125inter8));
  nand2 gate1956(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1957(.a(s_201), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1958(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1959(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1960(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2017(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2018(.a(gate127inter0), .b(s_210), .O(gate127inter1));
  and2  gate2019(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2020(.a(s_210), .O(gate127inter3));
  inv1  gate2021(.a(s_211), .O(gate127inter4));
  nand2 gate2022(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2023(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2024(.a(G406), .O(gate127inter7));
  inv1  gate2025(.a(G407), .O(gate127inter8));
  nand2 gate2026(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2027(.a(s_211), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2028(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2029(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2030(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1317(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1318(.a(gate128inter0), .b(s_110), .O(gate128inter1));
  and2  gate1319(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1320(.a(s_110), .O(gate128inter3));
  inv1  gate1321(.a(s_111), .O(gate128inter4));
  nand2 gate1322(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1323(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1324(.a(G408), .O(gate128inter7));
  inv1  gate1325(.a(G409), .O(gate128inter8));
  nand2 gate1326(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1327(.a(s_111), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1328(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1329(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1330(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1261(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1262(.a(gate129inter0), .b(s_102), .O(gate129inter1));
  and2  gate1263(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1264(.a(s_102), .O(gate129inter3));
  inv1  gate1265(.a(s_103), .O(gate129inter4));
  nand2 gate1266(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1267(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1268(.a(G410), .O(gate129inter7));
  inv1  gate1269(.a(G411), .O(gate129inter8));
  nand2 gate1270(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1271(.a(s_103), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1272(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1273(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1274(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate967(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate968(.a(gate130inter0), .b(s_60), .O(gate130inter1));
  and2  gate969(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate970(.a(s_60), .O(gate130inter3));
  inv1  gate971(.a(s_61), .O(gate130inter4));
  nand2 gate972(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate973(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate974(.a(G412), .O(gate130inter7));
  inv1  gate975(.a(G413), .O(gate130inter8));
  nand2 gate976(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate977(.a(s_61), .b(gate130inter3), .O(gate130inter10));
  nor2  gate978(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate979(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate980(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate3039(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate3040(.a(gate131inter0), .b(s_356), .O(gate131inter1));
  and2  gate3041(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate3042(.a(s_356), .O(gate131inter3));
  inv1  gate3043(.a(s_357), .O(gate131inter4));
  nand2 gate3044(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate3045(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate3046(.a(G414), .O(gate131inter7));
  inv1  gate3047(.a(G415), .O(gate131inter8));
  nand2 gate3048(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate3049(.a(s_357), .b(gate131inter3), .O(gate131inter10));
  nor2  gate3050(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate3051(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate3052(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate1331(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1332(.a(gate132inter0), .b(s_112), .O(gate132inter1));
  and2  gate1333(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1334(.a(s_112), .O(gate132inter3));
  inv1  gate1335(.a(s_113), .O(gate132inter4));
  nand2 gate1336(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1337(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1338(.a(G416), .O(gate132inter7));
  inv1  gate1339(.a(G417), .O(gate132inter8));
  nand2 gate1340(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1341(.a(s_113), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1342(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1343(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1344(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2633(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2634(.a(gate135inter0), .b(s_298), .O(gate135inter1));
  and2  gate2635(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2636(.a(s_298), .O(gate135inter3));
  inv1  gate2637(.a(s_299), .O(gate135inter4));
  nand2 gate2638(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2639(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2640(.a(G422), .O(gate135inter7));
  inv1  gate2641(.a(G423), .O(gate135inter8));
  nand2 gate2642(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2643(.a(s_299), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2644(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2645(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2646(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate603(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate604(.a(gate139inter0), .b(s_8), .O(gate139inter1));
  and2  gate605(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate606(.a(s_8), .O(gate139inter3));
  inv1  gate607(.a(s_9), .O(gate139inter4));
  nand2 gate608(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate609(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate610(.a(G438), .O(gate139inter7));
  inv1  gate611(.a(G441), .O(gate139inter8));
  nand2 gate612(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate613(.a(s_9), .b(gate139inter3), .O(gate139inter10));
  nor2  gate614(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate615(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate616(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1163(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1164(.a(gate140inter0), .b(s_88), .O(gate140inter1));
  and2  gate1165(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1166(.a(s_88), .O(gate140inter3));
  inv1  gate1167(.a(s_89), .O(gate140inter4));
  nand2 gate1168(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1169(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1170(.a(G444), .O(gate140inter7));
  inv1  gate1171(.a(G447), .O(gate140inter8));
  nand2 gate1172(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1173(.a(s_89), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1174(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1175(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1176(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate1891(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1892(.a(gate141inter0), .b(s_192), .O(gate141inter1));
  and2  gate1893(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1894(.a(s_192), .O(gate141inter3));
  inv1  gate1895(.a(s_193), .O(gate141inter4));
  nand2 gate1896(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1897(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1898(.a(G450), .O(gate141inter7));
  inv1  gate1899(.a(G453), .O(gate141inter8));
  nand2 gate1900(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1901(.a(s_193), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1902(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1903(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1904(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2269(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2270(.a(gate143inter0), .b(s_246), .O(gate143inter1));
  and2  gate2271(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2272(.a(s_246), .O(gate143inter3));
  inv1  gate2273(.a(s_247), .O(gate143inter4));
  nand2 gate2274(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2275(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2276(.a(G462), .O(gate143inter7));
  inv1  gate2277(.a(G465), .O(gate143inter8));
  nand2 gate2278(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2279(.a(s_247), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2280(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2281(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2282(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1135(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1136(.a(gate149inter0), .b(s_84), .O(gate149inter1));
  and2  gate1137(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1138(.a(s_84), .O(gate149inter3));
  inv1  gate1139(.a(s_85), .O(gate149inter4));
  nand2 gate1140(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1141(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1142(.a(G498), .O(gate149inter7));
  inv1  gate1143(.a(G501), .O(gate149inter8));
  nand2 gate1144(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1145(.a(s_85), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1146(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1147(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1148(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate827(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate828(.a(gate150inter0), .b(s_40), .O(gate150inter1));
  and2  gate829(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate830(.a(s_40), .O(gate150inter3));
  inv1  gate831(.a(s_41), .O(gate150inter4));
  nand2 gate832(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate833(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate834(.a(G504), .O(gate150inter7));
  inv1  gate835(.a(G507), .O(gate150inter8));
  nand2 gate836(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate837(.a(s_41), .b(gate150inter3), .O(gate150inter10));
  nor2  gate838(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate839(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate840(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate2675(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2676(.a(gate151inter0), .b(s_304), .O(gate151inter1));
  and2  gate2677(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2678(.a(s_304), .O(gate151inter3));
  inv1  gate2679(.a(s_305), .O(gate151inter4));
  nand2 gate2680(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2681(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2682(.a(G510), .O(gate151inter7));
  inv1  gate2683(.a(G513), .O(gate151inter8));
  nand2 gate2684(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2685(.a(s_305), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2686(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2687(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2688(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate2787(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2788(.a(gate152inter0), .b(s_320), .O(gate152inter1));
  and2  gate2789(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2790(.a(s_320), .O(gate152inter3));
  inv1  gate2791(.a(s_321), .O(gate152inter4));
  nand2 gate2792(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2793(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2794(.a(G516), .O(gate152inter7));
  inv1  gate2795(.a(G519), .O(gate152inter8));
  nand2 gate2796(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2797(.a(s_321), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2798(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2799(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2800(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2563(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2564(.a(gate155inter0), .b(s_288), .O(gate155inter1));
  and2  gate2565(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2566(.a(s_288), .O(gate155inter3));
  inv1  gate2567(.a(s_289), .O(gate155inter4));
  nand2 gate2568(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2569(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2570(.a(G432), .O(gate155inter7));
  inv1  gate2571(.a(G525), .O(gate155inter8));
  nand2 gate2572(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2573(.a(s_289), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2574(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2575(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2576(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2353(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2354(.a(gate157inter0), .b(s_258), .O(gate157inter1));
  and2  gate2355(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2356(.a(s_258), .O(gate157inter3));
  inv1  gate2357(.a(s_259), .O(gate157inter4));
  nand2 gate2358(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2359(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2360(.a(G438), .O(gate157inter7));
  inv1  gate2361(.a(G528), .O(gate157inter8));
  nand2 gate2362(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2363(.a(s_259), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2364(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2365(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2366(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2423(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2424(.a(gate158inter0), .b(s_268), .O(gate158inter1));
  and2  gate2425(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2426(.a(s_268), .O(gate158inter3));
  inv1  gate2427(.a(s_269), .O(gate158inter4));
  nand2 gate2428(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2429(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2430(.a(G441), .O(gate158inter7));
  inv1  gate2431(.a(G528), .O(gate158inter8));
  nand2 gate2432(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2433(.a(s_269), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2434(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2435(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2436(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2479(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2480(.a(gate159inter0), .b(s_276), .O(gate159inter1));
  and2  gate2481(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2482(.a(s_276), .O(gate159inter3));
  inv1  gate2483(.a(s_277), .O(gate159inter4));
  nand2 gate2484(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2485(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2486(.a(G444), .O(gate159inter7));
  inv1  gate2487(.a(G531), .O(gate159inter8));
  nand2 gate2488(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2489(.a(s_277), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2490(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2491(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2492(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2549(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2550(.a(gate160inter0), .b(s_286), .O(gate160inter1));
  and2  gate2551(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2552(.a(s_286), .O(gate160inter3));
  inv1  gate2553(.a(s_287), .O(gate160inter4));
  nand2 gate2554(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2555(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2556(.a(G447), .O(gate160inter7));
  inv1  gate2557(.a(G531), .O(gate160inter8));
  nand2 gate2558(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2559(.a(s_287), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2560(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2561(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2562(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate2493(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2494(.a(gate163inter0), .b(s_278), .O(gate163inter1));
  and2  gate2495(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2496(.a(s_278), .O(gate163inter3));
  inv1  gate2497(.a(s_279), .O(gate163inter4));
  nand2 gate2498(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2499(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2500(.a(G456), .O(gate163inter7));
  inv1  gate2501(.a(G537), .O(gate163inter8));
  nand2 gate2502(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2503(.a(s_279), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2504(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2505(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2506(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2367(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2368(.a(gate165inter0), .b(s_260), .O(gate165inter1));
  and2  gate2369(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2370(.a(s_260), .O(gate165inter3));
  inv1  gate2371(.a(s_261), .O(gate165inter4));
  nand2 gate2372(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2373(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2374(.a(G462), .O(gate165inter7));
  inv1  gate2375(.a(G540), .O(gate165inter8));
  nand2 gate2376(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2377(.a(s_261), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2378(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2379(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2380(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1835(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1836(.a(gate166inter0), .b(s_184), .O(gate166inter1));
  and2  gate1837(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1838(.a(s_184), .O(gate166inter3));
  inv1  gate1839(.a(s_185), .O(gate166inter4));
  nand2 gate1840(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1841(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1842(.a(G465), .O(gate166inter7));
  inv1  gate1843(.a(G540), .O(gate166inter8));
  nand2 gate1844(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1845(.a(s_185), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1846(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1847(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1848(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate3151(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate3152(.a(gate167inter0), .b(s_372), .O(gate167inter1));
  and2  gate3153(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate3154(.a(s_372), .O(gate167inter3));
  inv1  gate3155(.a(s_373), .O(gate167inter4));
  nand2 gate3156(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate3157(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate3158(.a(G468), .O(gate167inter7));
  inv1  gate3159(.a(G543), .O(gate167inter8));
  nand2 gate3160(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate3161(.a(s_373), .b(gate167inter3), .O(gate167inter10));
  nor2  gate3162(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate3163(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate3164(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate2227(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate2228(.a(gate168inter0), .b(s_240), .O(gate168inter1));
  and2  gate2229(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate2230(.a(s_240), .O(gate168inter3));
  inv1  gate2231(.a(s_241), .O(gate168inter4));
  nand2 gate2232(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate2233(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate2234(.a(G471), .O(gate168inter7));
  inv1  gate2235(.a(G543), .O(gate168inter8));
  nand2 gate2236(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate2237(.a(s_241), .b(gate168inter3), .O(gate168inter10));
  nor2  gate2238(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate2239(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate2240(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1401(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1402(.a(gate169inter0), .b(s_122), .O(gate169inter1));
  and2  gate1403(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1404(.a(s_122), .O(gate169inter3));
  inv1  gate1405(.a(s_123), .O(gate169inter4));
  nand2 gate1406(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1407(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1408(.a(G474), .O(gate169inter7));
  inv1  gate1409(.a(G546), .O(gate169inter8));
  nand2 gate1410(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1411(.a(s_123), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1412(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1413(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1414(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2087(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2088(.a(gate170inter0), .b(s_220), .O(gate170inter1));
  and2  gate2089(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2090(.a(s_220), .O(gate170inter3));
  inv1  gate2091(.a(s_221), .O(gate170inter4));
  nand2 gate2092(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2093(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2094(.a(G477), .O(gate170inter7));
  inv1  gate2095(.a(G546), .O(gate170inter8));
  nand2 gate2096(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2097(.a(s_221), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2098(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2099(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2100(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1583(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1584(.a(gate171inter0), .b(s_148), .O(gate171inter1));
  and2  gate1585(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1586(.a(s_148), .O(gate171inter3));
  inv1  gate1587(.a(s_149), .O(gate171inter4));
  nand2 gate1588(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1589(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1590(.a(G480), .O(gate171inter7));
  inv1  gate1591(.a(G549), .O(gate171inter8));
  nand2 gate1592(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1593(.a(s_149), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1594(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1595(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1596(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1737(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1738(.a(gate173inter0), .b(s_170), .O(gate173inter1));
  and2  gate1739(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1740(.a(s_170), .O(gate173inter3));
  inv1  gate1741(.a(s_171), .O(gate173inter4));
  nand2 gate1742(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1743(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1744(.a(G486), .O(gate173inter7));
  inv1  gate1745(.a(G552), .O(gate173inter8));
  nand2 gate1746(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1747(.a(s_171), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1748(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1749(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1750(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2661(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2662(.a(gate176inter0), .b(s_302), .O(gate176inter1));
  and2  gate2663(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2664(.a(s_302), .O(gate176inter3));
  inv1  gate2665(.a(s_303), .O(gate176inter4));
  nand2 gate2666(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2667(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2668(.a(G495), .O(gate176inter7));
  inv1  gate2669(.a(G555), .O(gate176inter8));
  nand2 gate2670(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2671(.a(s_303), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2672(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2673(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2674(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate617(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate618(.a(gate177inter0), .b(s_10), .O(gate177inter1));
  and2  gate619(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate620(.a(s_10), .O(gate177inter3));
  inv1  gate621(.a(s_11), .O(gate177inter4));
  nand2 gate622(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate623(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate624(.a(G498), .O(gate177inter7));
  inv1  gate625(.a(G558), .O(gate177inter8));
  nand2 gate626(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate627(.a(s_11), .b(gate177inter3), .O(gate177inter10));
  nor2  gate628(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate629(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate630(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1093(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1094(.a(gate178inter0), .b(s_78), .O(gate178inter1));
  and2  gate1095(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1096(.a(s_78), .O(gate178inter3));
  inv1  gate1097(.a(s_79), .O(gate178inter4));
  nand2 gate1098(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1099(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1100(.a(G501), .O(gate178inter7));
  inv1  gate1101(.a(G558), .O(gate178inter8));
  nand2 gate1102(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1103(.a(s_79), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1104(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1105(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1106(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate3263(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate3264(.a(gate179inter0), .b(s_388), .O(gate179inter1));
  and2  gate3265(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate3266(.a(s_388), .O(gate179inter3));
  inv1  gate3267(.a(s_389), .O(gate179inter4));
  nand2 gate3268(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate3269(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate3270(.a(G504), .O(gate179inter7));
  inv1  gate3271(.a(G561), .O(gate179inter8));
  nand2 gate3272(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate3273(.a(s_389), .b(gate179inter3), .O(gate179inter10));
  nor2  gate3274(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate3275(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate3276(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1149(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1150(.a(gate182inter0), .b(s_86), .O(gate182inter1));
  and2  gate1151(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1152(.a(s_86), .O(gate182inter3));
  inv1  gate1153(.a(s_87), .O(gate182inter4));
  nand2 gate1154(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1155(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1156(.a(G513), .O(gate182inter7));
  inv1  gate1157(.a(G564), .O(gate182inter8));
  nand2 gate1158(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1159(.a(s_87), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1160(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1161(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1162(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate2451(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2452(.a(gate183inter0), .b(s_272), .O(gate183inter1));
  and2  gate2453(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2454(.a(s_272), .O(gate183inter3));
  inv1  gate2455(.a(s_273), .O(gate183inter4));
  nand2 gate2456(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2457(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2458(.a(G516), .O(gate183inter7));
  inv1  gate2459(.a(G567), .O(gate183inter8));
  nand2 gate2460(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2461(.a(s_273), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2462(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2463(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2464(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate3053(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate3054(.a(gate185inter0), .b(s_358), .O(gate185inter1));
  and2  gate3055(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate3056(.a(s_358), .O(gate185inter3));
  inv1  gate3057(.a(s_359), .O(gate185inter4));
  nand2 gate3058(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate3059(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate3060(.a(G570), .O(gate185inter7));
  inv1  gate3061(.a(G571), .O(gate185inter8));
  nand2 gate3062(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate3063(.a(s_359), .b(gate185inter3), .O(gate185inter10));
  nor2  gate3064(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate3065(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate3066(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate3347(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate3348(.a(gate186inter0), .b(s_400), .O(gate186inter1));
  and2  gate3349(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate3350(.a(s_400), .O(gate186inter3));
  inv1  gate3351(.a(s_401), .O(gate186inter4));
  nand2 gate3352(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate3353(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate3354(.a(G572), .O(gate186inter7));
  inv1  gate3355(.a(G573), .O(gate186inter8));
  nand2 gate3356(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate3357(.a(s_401), .b(gate186inter3), .O(gate186inter10));
  nor2  gate3358(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate3359(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate3360(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1485(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1486(.a(gate188inter0), .b(s_134), .O(gate188inter1));
  and2  gate1487(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1488(.a(s_134), .O(gate188inter3));
  inv1  gate1489(.a(s_135), .O(gate188inter4));
  nand2 gate1490(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1491(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1492(.a(G576), .O(gate188inter7));
  inv1  gate1493(.a(G577), .O(gate188inter8));
  nand2 gate1494(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1495(.a(s_135), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1496(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1497(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1498(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate771(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate772(.a(gate191inter0), .b(s_32), .O(gate191inter1));
  and2  gate773(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate774(.a(s_32), .O(gate191inter3));
  inv1  gate775(.a(s_33), .O(gate191inter4));
  nand2 gate776(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate777(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate778(.a(G582), .O(gate191inter7));
  inv1  gate779(.a(G583), .O(gate191inter8));
  nand2 gate780(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate781(.a(s_33), .b(gate191inter3), .O(gate191inter10));
  nor2  gate782(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate783(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate784(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1429(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1430(.a(gate193inter0), .b(s_126), .O(gate193inter1));
  and2  gate1431(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1432(.a(s_126), .O(gate193inter3));
  inv1  gate1433(.a(s_127), .O(gate193inter4));
  nand2 gate1434(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1435(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1436(.a(G586), .O(gate193inter7));
  inv1  gate1437(.a(G587), .O(gate193inter8));
  nand2 gate1438(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1439(.a(s_127), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1440(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1441(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1442(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate2129(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2130(.a(gate194inter0), .b(s_226), .O(gate194inter1));
  and2  gate2131(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2132(.a(s_226), .O(gate194inter3));
  inv1  gate2133(.a(s_227), .O(gate194inter4));
  nand2 gate2134(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2135(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2136(.a(G588), .O(gate194inter7));
  inv1  gate2137(.a(G589), .O(gate194inter8));
  nand2 gate2138(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2139(.a(s_227), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2140(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2141(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2142(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2927(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2928(.a(gate198inter0), .b(s_340), .O(gate198inter1));
  and2  gate2929(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2930(.a(s_340), .O(gate198inter3));
  inv1  gate2931(.a(s_341), .O(gate198inter4));
  nand2 gate2932(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2933(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2934(.a(G596), .O(gate198inter7));
  inv1  gate2935(.a(G597), .O(gate198inter8));
  nand2 gate2936(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2937(.a(s_341), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2938(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2939(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2940(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1121(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1122(.a(gate200inter0), .b(s_82), .O(gate200inter1));
  and2  gate1123(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1124(.a(s_82), .O(gate200inter3));
  inv1  gate1125(.a(s_83), .O(gate200inter4));
  nand2 gate1126(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1127(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1128(.a(G600), .O(gate200inter7));
  inv1  gate1129(.a(G601), .O(gate200inter8));
  nand2 gate1130(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1131(.a(s_83), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1132(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1133(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1134(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1905(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1906(.a(gate201inter0), .b(s_194), .O(gate201inter1));
  and2  gate1907(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1908(.a(s_194), .O(gate201inter3));
  inv1  gate1909(.a(s_195), .O(gate201inter4));
  nand2 gate1910(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1911(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1912(.a(G602), .O(gate201inter7));
  inv1  gate1913(.a(G607), .O(gate201inter8));
  nand2 gate1914(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1915(.a(s_195), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1916(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1917(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1918(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate2521(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate2522(.a(gate202inter0), .b(s_282), .O(gate202inter1));
  and2  gate2523(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate2524(.a(s_282), .O(gate202inter3));
  inv1  gate2525(.a(s_283), .O(gate202inter4));
  nand2 gate2526(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate2527(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate2528(.a(G612), .O(gate202inter7));
  inv1  gate2529(.a(G617), .O(gate202inter8));
  nand2 gate2530(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate2531(.a(s_283), .b(gate202inter3), .O(gate202inter10));
  nor2  gate2532(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate2533(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate2534(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate3221(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate3222(.a(gate205inter0), .b(s_382), .O(gate205inter1));
  and2  gate3223(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate3224(.a(s_382), .O(gate205inter3));
  inv1  gate3225(.a(s_383), .O(gate205inter4));
  nand2 gate3226(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate3227(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate3228(.a(G622), .O(gate205inter7));
  inv1  gate3229(.a(G627), .O(gate205inter8));
  nand2 gate3230(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate3231(.a(s_383), .b(gate205inter3), .O(gate205inter10));
  nor2  gate3232(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate3233(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate3234(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2115(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2116(.a(gate206inter0), .b(s_224), .O(gate206inter1));
  and2  gate2117(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2118(.a(s_224), .O(gate206inter3));
  inv1  gate2119(.a(s_225), .O(gate206inter4));
  nand2 gate2120(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2121(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2122(.a(G632), .O(gate206inter7));
  inv1  gate2123(.a(G637), .O(gate206inter8));
  nand2 gate2124(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2125(.a(s_225), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2126(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2127(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2128(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1695(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1696(.a(gate207inter0), .b(s_164), .O(gate207inter1));
  and2  gate1697(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1698(.a(s_164), .O(gate207inter3));
  inv1  gate1699(.a(s_165), .O(gate207inter4));
  nand2 gate1700(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1701(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1702(.a(G622), .O(gate207inter7));
  inv1  gate1703(.a(G632), .O(gate207inter8));
  nand2 gate1704(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1705(.a(s_165), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1706(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1707(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1708(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate743(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate744(.a(gate208inter0), .b(s_28), .O(gate208inter1));
  and2  gate745(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate746(.a(s_28), .O(gate208inter3));
  inv1  gate747(.a(s_29), .O(gate208inter4));
  nand2 gate748(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate749(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate750(.a(G627), .O(gate208inter7));
  inv1  gate751(.a(G637), .O(gate208inter8));
  nand2 gate752(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate753(.a(s_29), .b(gate208inter3), .O(gate208inter10));
  nor2  gate754(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate755(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate756(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1275(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1276(.a(gate209inter0), .b(s_104), .O(gate209inter1));
  and2  gate1277(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1278(.a(s_104), .O(gate209inter3));
  inv1  gate1279(.a(s_105), .O(gate209inter4));
  nand2 gate1280(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1281(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1282(.a(G602), .O(gate209inter7));
  inv1  gate1283(.a(G666), .O(gate209inter8));
  nand2 gate1284(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1285(.a(s_105), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1286(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1287(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1288(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1051(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1052(.a(gate210inter0), .b(s_72), .O(gate210inter1));
  and2  gate1053(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1054(.a(s_72), .O(gate210inter3));
  inv1  gate1055(.a(s_73), .O(gate210inter4));
  nand2 gate1056(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1057(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1058(.a(G607), .O(gate210inter7));
  inv1  gate1059(.a(G666), .O(gate210inter8));
  nand2 gate1060(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1061(.a(s_73), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1062(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1063(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1064(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate2101(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2102(.a(gate211inter0), .b(s_222), .O(gate211inter1));
  and2  gate2103(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2104(.a(s_222), .O(gate211inter3));
  inv1  gate2105(.a(s_223), .O(gate211inter4));
  nand2 gate2106(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2107(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2108(.a(G612), .O(gate211inter7));
  inv1  gate2109(.a(G669), .O(gate211inter8));
  nand2 gate2110(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2111(.a(s_223), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2112(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2113(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2114(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1765(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1766(.a(gate214inter0), .b(s_174), .O(gate214inter1));
  and2  gate1767(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1768(.a(s_174), .O(gate214inter3));
  inv1  gate1769(.a(s_175), .O(gate214inter4));
  nand2 gate1770(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1771(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1772(.a(G612), .O(gate214inter7));
  inv1  gate1773(.a(G672), .O(gate214inter8));
  nand2 gate1774(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1775(.a(s_175), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1776(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1777(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1778(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1345(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1346(.a(gate219inter0), .b(s_114), .O(gate219inter1));
  and2  gate1347(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1348(.a(s_114), .O(gate219inter3));
  inv1  gate1349(.a(s_115), .O(gate219inter4));
  nand2 gate1350(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1351(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1352(.a(G632), .O(gate219inter7));
  inv1  gate1353(.a(G681), .O(gate219inter8));
  nand2 gate1354(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1355(.a(s_115), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1356(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1357(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1358(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate575(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate576(.a(gate222inter0), .b(s_4), .O(gate222inter1));
  and2  gate577(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate578(.a(s_4), .O(gate222inter3));
  inv1  gate579(.a(s_5), .O(gate222inter4));
  nand2 gate580(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate581(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate582(.a(G632), .O(gate222inter7));
  inv1  gate583(.a(G684), .O(gate222inter8));
  nand2 gate584(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate585(.a(s_5), .b(gate222inter3), .O(gate222inter10));
  nor2  gate586(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate587(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate588(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2759(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2760(.a(gate223inter0), .b(s_316), .O(gate223inter1));
  and2  gate2761(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2762(.a(s_316), .O(gate223inter3));
  inv1  gate2763(.a(s_317), .O(gate223inter4));
  nand2 gate2764(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2765(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2766(.a(G627), .O(gate223inter7));
  inv1  gate2767(.a(G687), .O(gate223inter8));
  nand2 gate2768(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2769(.a(s_317), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2770(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2771(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2772(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1303(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1304(.a(gate226inter0), .b(s_108), .O(gate226inter1));
  and2  gate1305(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1306(.a(s_108), .O(gate226inter3));
  inv1  gate1307(.a(s_109), .O(gate226inter4));
  nand2 gate1308(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1309(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1310(.a(G692), .O(gate226inter7));
  inv1  gate1311(.a(G693), .O(gate226inter8));
  nand2 gate1312(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1313(.a(s_109), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1314(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1315(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1316(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1597(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1598(.a(gate229inter0), .b(s_150), .O(gate229inter1));
  and2  gate1599(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1600(.a(s_150), .O(gate229inter3));
  inv1  gate1601(.a(s_151), .O(gate229inter4));
  nand2 gate1602(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1603(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1604(.a(G698), .O(gate229inter7));
  inv1  gate1605(.a(G699), .O(gate229inter8));
  nand2 gate1606(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1607(.a(s_151), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1608(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1609(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1610(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate2143(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2144(.a(gate230inter0), .b(s_228), .O(gate230inter1));
  and2  gate2145(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2146(.a(s_228), .O(gate230inter3));
  inv1  gate2147(.a(s_229), .O(gate230inter4));
  nand2 gate2148(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2149(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2150(.a(G700), .O(gate230inter7));
  inv1  gate2151(.a(G701), .O(gate230inter8));
  nand2 gate2152(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2153(.a(s_229), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2154(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2155(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2156(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1723(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1724(.a(gate231inter0), .b(s_168), .O(gate231inter1));
  and2  gate1725(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1726(.a(s_168), .O(gate231inter3));
  inv1  gate1727(.a(s_169), .O(gate231inter4));
  nand2 gate1728(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1729(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1730(.a(G702), .O(gate231inter7));
  inv1  gate1731(.a(G703), .O(gate231inter8));
  nand2 gate1732(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1733(.a(s_169), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1734(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1735(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1736(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate2885(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2886(.a(gate235inter0), .b(s_334), .O(gate235inter1));
  and2  gate2887(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2888(.a(s_334), .O(gate235inter3));
  inv1  gate2889(.a(s_335), .O(gate235inter4));
  nand2 gate2890(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2891(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2892(.a(G248), .O(gate235inter7));
  inv1  gate2893(.a(G724), .O(gate235inter8));
  nand2 gate2894(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2895(.a(s_335), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2896(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2897(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2898(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate1023(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1024(.a(gate236inter0), .b(s_68), .O(gate236inter1));
  and2  gate1025(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1026(.a(s_68), .O(gate236inter3));
  inv1  gate1027(.a(s_69), .O(gate236inter4));
  nand2 gate1028(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1029(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1030(.a(G251), .O(gate236inter7));
  inv1  gate1031(.a(G727), .O(gate236inter8));
  nand2 gate1032(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1033(.a(s_69), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1034(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1035(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1036(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate841(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate842(.a(gate238inter0), .b(s_42), .O(gate238inter1));
  and2  gate843(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate844(.a(s_42), .O(gate238inter3));
  inv1  gate845(.a(s_43), .O(gate238inter4));
  nand2 gate846(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate847(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate848(.a(G257), .O(gate238inter7));
  inv1  gate849(.a(G709), .O(gate238inter8));
  nand2 gate850(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate851(.a(s_43), .b(gate238inter3), .O(gate238inter10));
  nor2  gate852(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate853(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate854(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1247(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1248(.a(gate240inter0), .b(s_100), .O(gate240inter1));
  and2  gate1249(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1250(.a(s_100), .O(gate240inter3));
  inv1  gate1251(.a(s_101), .O(gate240inter4));
  nand2 gate1252(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1253(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1254(.a(G263), .O(gate240inter7));
  inv1  gate1255(.a(G715), .O(gate240inter8));
  nand2 gate1256(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1257(.a(s_101), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1258(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1259(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1260(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate3165(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate3166(.a(gate242inter0), .b(s_374), .O(gate242inter1));
  and2  gate3167(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate3168(.a(s_374), .O(gate242inter3));
  inv1  gate3169(.a(s_375), .O(gate242inter4));
  nand2 gate3170(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate3171(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate3172(.a(G718), .O(gate242inter7));
  inv1  gate3173(.a(G730), .O(gate242inter8));
  nand2 gate3174(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate3175(.a(s_375), .b(gate242inter3), .O(gate242inter10));
  nor2  gate3176(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate3177(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate3178(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate3319(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate3320(.a(gate246inter0), .b(s_396), .O(gate246inter1));
  and2  gate3321(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate3322(.a(s_396), .O(gate246inter3));
  inv1  gate3323(.a(s_397), .O(gate246inter4));
  nand2 gate3324(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate3325(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate3326(.a(G724), .O(gate246inter7));
  inv1  gate3327(.a(G736), .O(gate246inter8));
  nand2 gate3328(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate3329(.a(s_397), .b(gate246inter3), .O(gate246inter10));
  nor2  gate3330(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate3331(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate3332(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1681(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1682(.a(gate250inter0), .b(s_162), .O(gate250inter1));
  and2  gate1683(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1684(.a(s_162), .O(gate250inter3));
  inv1  gate1685(.a(s_163), .O(gate250inter4));
  nand2 gate1686(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1687(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1688(.a(G706), .O(gate250inter7));
  inv1  gate1689(.a(G742), .O(gate250inter8));
  nand2 gate1690(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1691(.a(s_163), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1692(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1693(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1694(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2801(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2802(.a(gate256inter0), .b(s_322), .O(gate256inter1));
  and2  gate2803(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2804(.a(s_322), .O(gate256inter3));
  inv1  gate2805(.a(s_323), .O(gate256inter4));
  nand2 gate2806(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2807(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2808(.a(G715), .O(gate256inter7));
  inv1  gate2809(.a(G751), .O(gate256inter8));
  nand2 gate2810(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2811(.a(s_323), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2812(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2813(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2814(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1513(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1514(.a(gate257inter0), .b(s_138), .O(gate257inter1));
  and2  gate1515(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1516(.a(s_138), .O(gate257inter3));
  inv1  gate1517(.a(s_139), .O(gate257inter4));
  nand2 gate1518(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1519(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1520(.a(G754), .O(gate257inter7));
  inv1  gate1521(.a(G755), .O(gate257inter8));
  nand2 gate1522(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1523(.a(s_139), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1524(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1525(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1526(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate3305(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate3306(.a(gate258inter0), .b(s_394), .O(gate258inter1));
  and2  gate3307(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate3308(.a(s_394), .O(gate258inter3));
  inv1  gate3309(.a(s_395), .O(gate258inter4));
  nand2 gate3310(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate3311(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate3312(.a(G756), .O(gate258inter7));
  inv1  gate3313(.a(G757), .O(gate258inter8));
  nand2 gate3314(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate3315(.a(s_395), .b(gate258inter3), .O(gate258inter10));
  nor2  gate3316(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate3317(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate3318(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1863(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1864(.a(gate262inter0), .b(s_188), .O(gate262inter1));
  and2  gate1865(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1866(.a(s_188), .O(gate262inter3));
  inv1  gate1867(.a(s_189), .O(gate262inter4));
  nand2 gate1868(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1869(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1870(.a(G764), .O(gate262inter7));
  inv1  gate1871(.a(G765), .O(gate262inter8));
  nand2 gate1872(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1873(.a(s_189), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1874(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1875(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1876(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate883(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate884(.a(gate263inter0), .b(s_48), .O(gate263inter1));
  and2  gate885(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate886(.a(s_48), .O(gate263inter3));
  inv1  gate887(.a(s_49), .O(gate263inter4));
  nand2 gate888(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate889(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate890(.a(G766), .O(gate263inter7));
  inv1  gate891(.a(G767), .O(gate263inter8));
  nand2 gate892(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate893(.a(s_49), .b(gate263inter3), .O(gate263inter10));
  nor2  gate894(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate895(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate896(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1779(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1780(.a(gate264inter0), .b(s_176), .O(gate264inter1));
  and2  gate1781(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1782(.a(s_176), .O(gate264inter3));
  inv1  gate1783(.a(s_177), .O(gate264inter4));
  nand2 gate1784(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1785(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1786(.a(G768), .O(gate264inter7));
  inv1  gate1787(.a(G769), .O(gate264inter8));
  nand2 gate1788(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1789(.a(s_177), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1790(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1791(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1792(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate547(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate548(.a(gate265inter0), .b(s_0), .O(gate265inter1));
  and2  gate549(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate550(.a(s_0), .O(gate265inter3));
  inv1  gate551(.a(s_1), .O(gate265inter4));
  nand2 gate552(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate553(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate554(.a(G642), .O(gate265inter7));
  inv1  gate555(.a(G770), .O(gate265inter8));
  nand2 gate556(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate557(.a(s_1), .b(gate265inter3), .O(gate265inter10));
  nor2  gate558(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate559(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate560(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2997(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2998(.a(gate267inter0), .b(s_350), .O(gate267inter1));
  and2  gate2999(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate3000(.a(s_350), .O(gate267inter3));
  inv1  gate3001(.a(s_351), .O(gate267inter4));
  nand2 gate3002(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate3003(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate3004(.a(G648), .O(gate267inter7));
  inv1  gate3005(.a(G776), .O(gate267inter8));
  nand2 gate3006(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate3007(.a(s_351), .b(gate267inter3), .O(gate267inter10));
  nor2  gate3008(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate3009(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate3010(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate2213(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2214(.a(gate272inter0), .b(s_238), .O(gate272inter1));
  and2  gate2215(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2216(.a(s_238), .O(gate272inter3));
  inv1  gate2217(.a(s_239), .O(gate272inter4));
  nand2 gate2218(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2219(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2220(.a(G663), .O(gate272inter7));
  inv1  gate2221(.a(G791), .O(gate272inter8));
  nand2 gate2222(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2223(.a(s_239), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2224(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2225(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2226(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate3207(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate3208(.a(gate273inter0), .b(s_380), .O(gate273inter1));
  and2  gate3209(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate3210(.a(s_380), .O(gate273inter3));
  inv1  gate3211(.a(s_381), .O(gate273inter4));
  nand2 gate3212(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate3213(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate3214(.a(G642), .O(gate273inter7));
  inv1  gate3215(.a(G794), .O(gate273inter8));
  nand2 gate3216(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate3217(.a(s_381), .b(gate273inter3), .O(gate273inter10));
  nor2  gate3218(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate3219(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate3220(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2325(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2326(.a(gate274inter0), .b(s_254), .O(gate274inter1));
  and2  gate2327(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2328(.a(s_254), .O(gate274inter3));
  inv1  gate2329(.a(s_255), .O(gate274inter4));
  nand2 gate2330(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2331(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2332(.a(G770), .O(gate274inter7));
  inv1  gate2333(.a(G794), .O(gate274inter8));
  nand2 gate2334(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2335(.a(s_255), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2336(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2337(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2338(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate785(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate786(.a(gate276inter0), .b(s_34), .O(gate276inter1));
  and2  gate787(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate788(.a(s_34), .O(gate276inter3));
  inv1  gate789(.a(s_35), .O(gate276inter4));
  nand2 gate790(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate791(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate792(.a(G773), .O(gate276inter7));
  inv1  gate793(.a(G797), .O(gate276inter8));
  nand2 gate794(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate795(.a(s_35), .b(gate276inter3), .O(gate276inter10));
  nor2  gate796(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate797(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate798(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate2185(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2186(.a(gate277inter0), .b(s_234), .O(gate277inter1));
  and2  gate2187(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2188(.a(s_234), .O(gate277inter3));
  inv1  gate2189(.a(s_235), .O(gate277inter4));
  nand2 gate2190(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2191(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2192(.a(G648), .O(gate277inter7));
  inv1  gate2193(.a(G800), .O(gate277inter8));
  nand2 gate2194(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2195(.a(s_235), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2196(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2197(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2198(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate855(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate856(.a(gate281inter0), .b(s_44), .O(gate281inter1));
  and2  gate857(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate858(.a(s_44), .O(gate281inter3));
  inv1  gate859(.a(s_45), .O(gate281inter4));
  nand2 gate860(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate861(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate862(.a(G654), .O(gate281inter7));
  inv1  gate863(.a(G806), .O(gate281inter8));
  nand2 gate864(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate865(.a(s_45), .b(gate281inter3), .O(gate281inter10));
  nor2  gate866(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate867(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate868(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1387(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1388(.a(gate283inter0), .b(s_120), .O(gate283inter1));
  and2  gate1389(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1390(.a(s_120), .O(gate283inter3));
  inv1  gate1391(.a(s_121), .O(gate283inter4));
  nand2 gate1392(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1393(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1394(.a(G657), .O(gate283inter7));
  inv1  gate1395(.a(G809), .O(gate283inter8));
  nand2 gate1396(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1397(.a(s_121), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1398(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1399(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1400(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate673(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate674(.a(gate293inter0), .b(s_18), .O(gate293inter1));
  and2  gate675(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate676(.a(s_18), .O(gate293inter3));
  inv1  gate677(.a(s_19), .O(gate293inter4));
  nand2 gate678(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate679(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate680(.a(G828), .O(gate293inter7));
  inv1  gate681(.a(G829), .O(gate293inter8));
  nand2 gate682(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate683(.a(s_19), .b(gate293inter3), .O(gate293inter10));
  nor2  gate684(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate685(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate686(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate2045(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2046(.a(gate294inter0), .b(s_214), .O(gate294inter1));
  and2  gate2047(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2048(.a(s_214), .O(gate294inter3));
  inv1  gate2049(.a(s_215), .O(gate294inter4));
  nand2 gate2050(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2051(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2052(.a(G832), .O(gate294inter7));
  inv1  gate2053(.a(G833), .O(gate294inter8));
  nand2 gate2054(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2055(.a(s_215), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2056(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2057(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2058(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate3291(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate3292(.a(gate296inter0), .b(s_392), .O(gate296inter1));
  and2  gate3293(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate3294(.a(s_392), .O(gate296inter3));
  inv1  gate3295(.a(s_393), .O(gate296inter4));
  nand2 gate3296(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate3297(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate3298(.a(G826), .O(gate296inter7));
  inv1  gate3299(.a(G827), .O(gate296inter8));
  nand2 gate3300(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate3301(.a(s_393), .b(gate296inter3), .O(gate296inter10));
  nor2  gate3302(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate3303(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate3304(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate3235(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate3236(.a(gate389inter0), .b(s_384), .O(gate389inter1));
  and2  gate3237(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate3238(.a(s_384), .O(gate389inter3));
  inv1  gate3239(.a(s_385), .O(gate389inter4));
  nand2 gate3240(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate3241(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate3242(.a(G3), .O(gate389inter7));
  inv1  gate3243(.a(G1042), .O(gate389inter8));
  nand2 gate3244(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate3245(.a(s_385), .b(gate389inter3), .O(gate389inter10));
  nor2  gate3246(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate3247(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate3248(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1009(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1010(.a(gate394inter0), .b(s_66), .O(gate394inter1));
  and2  gate1011(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1012(.a(s_66), .O(gate394inter3));
  inv1  gate1013(.a(s_67), .O(gate394inter4));
  nand2 gate1014(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1015(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1016(.a(G8), .O(gate394inter7));
  inv1  gate1017(.a(G1057), .O(gate394inter8));
  nand2 gate1018(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1019(.a(s_67), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1020(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1021(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1022(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate869(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate870(.a(gate399inter0), .b(s_46), .O(gate399inter1));
  and2  gate871(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate872(.a(s_46), .O(gate399inter3));
  inv1  gate873(.a(s_47), .O(gate399inter4));
  nand2 gate874(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate875(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate876(.a(G13), .O(gate399inter7));
  inv1  gate877(.a(G1072), .O(gate399inter8));
  nand2 gate878(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate879(.a(s_47), .b(gate399inter3), .O(gate399inter10));
  nor2  gate880(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate881(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate882(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1639(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1640(.a(gate400inter0), .b(s_156), .O(gate400inter1));
  and2  gate1641(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1642(.a(s_156), .O(gate400inter3));
  inv1  gate1643(.a(s_157), .O(gate400inter4));
  nand2 gate1644(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1645(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1646(.a(G14), .O(gate400inter7));
  inv1  gate1647(.a(G1075), .O(gate400inter8));
  nand2 gate1648(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1649(.a(s_157), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1650(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1651(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1652(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1989(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1990(.a(gate402inter0), .b(s_206), .O(gate402inter1));
  and2  gate1991(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1992(.a(s_206), .O(gate402inter3));
  inv1  gate1993(.a(s_207), .O(gate402inter4));
  nand2 gate1994(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1995(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1996(.a(G16), .O(gate402inter7));
  inv1  gate1997(.a(G1081), .O(gate402inter8));
  nand2 gate1998(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1999(.a(s_207), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2000(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2001(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2002(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1107(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1108(.a(gate405inter0), .b(s_80), .O(gate405inter1));
  and2  gate1109(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1110(.a(s_80), .O(gate405inter3));
  inv1  gate1111(.a(s_81), .O(gate405inter4));
  nand2 gate1112(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1113(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1114(.a(G19), .O(gate405inter7));
  inv1  gate1115(.a(G1090), .O(gate405inter8));
  nand2 gate1116(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1117(.a(s_81), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1118(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1119(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1120(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1933(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1934(.a(gate407inter0), .b(s_198), .O(gate407inter1));
  and2  gate1935(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1936(.a(s_198), .O(gate407inter3));
  inv1  gate1937(.a(s_199), .O(gate407inter4));
  nand2 gate1938(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1939(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1940(.a(G21), .O(gate407inter7));
  inv1  gate1941(.a(G1096), .O(gate407inter8));
  nand2 gate1942(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1943(.a(s_199), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1944(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1945(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1946(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate3137(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate3138(.a(gate408inter0), .b(s_370), .O(gate408inter1));
  and2  gate3139(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate3140(.a(s_370), .O(gate408inter3));
  inv1  gate3141(.a(s_371), .O(gate408inter4));
  nand2 gate3142(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate3143(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate3144(.a(G22), .O(gate408inter7));
  inv1  gate3145(.a(G1099), .O(gate408inter8));
  nand2 gate3146(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate3147(.a(s_371), .b(gate408inter3), .O(gate408inter10));
  nor2  gate3148(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate3149(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate3150(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2689(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2690(.a(gate410inter0), .b(s_306), .O(gate410inter1));
  and2  gate2691(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2692(.a(s_306), .O(gate410inter3));
  inv1  gate2693(.a(s_307), .O(gate410inter4));
  nand2 gate2694(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2695(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2696(.a(G24), .O(gate410inter7));
  inv1  gate2697(.a(G1105), .O(gate410inter8));
  nand2 gate2698(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2699(.a(s_307), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2700(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2701(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2702(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate2703(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2704(.a(gate411inter0), .b(s_308), .O(gate411inter1));
  and2  gate2705(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2706(.a(s_308), .O(gate411inter3));
  inv1  gate2707(.a(s_309), .O(gate411inter4));
  nand2 gate2708(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2709(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2710(.a(G25), .O(gate411inter7));
  inv1  gate2711(.a(G1108), .O(gate411inter8));
  nand2 gate2712(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2713(.a(s_309), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2714(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2715(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2716(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate645(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate646(.a(gate412inter0), .b(s_14), .O(gate412inter1));
  and2  gate647(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate648(.a(s_14), .O(gate412inter3));
  inv1  gate649(.a(s_15), .O(gate412inter4));
  nand2 gate650(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate651(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate652(.a(G26), .O(gate412inter7));
  inv1  gate653(.a(G1111), .O(gate412inter8));
  nand2 gate654(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate655(.a(s_15), .b(gate412inter3), .O(gate412inter10));
  nor2  gate656(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate657(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate658(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1191(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1192(.a(gate417inter0), .b(s_92), .O(gate417inter1));
  and2  gate1193(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1194(.a(s_92), .O(gate417inter3));
  inv1  gate1195(.a(s_93), .O(gate417inter4));
  nand2 gate1196(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1197(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1198(.a(G31), .O(gate417inter7));
  inv1  gate1199(.a(G1126), .O(gate417inter8));
  nand2 gate1200(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1201(.a(s_93), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1202(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1203(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1204(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1625(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1626(.a(gate418inter0), .b(s_154), .O(gate418inter1));
  and2  gate1627(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1628(.a(s_154), .O(gate418inter3));
  inv1  gate1629(.a(s_155), .O(gate418inter4));
  nand2 gate1630(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1631(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1632(.a(G32), .O(gate418inter7));
  inv1  gate1633(.a(G1129), .O(gate418inter8));
  nand2 gate1634(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1635(.a(s_155), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1636(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1637(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1638(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2059(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2060(.a(gate421inter0), .b(s_216), .O(gate421inter1));
  and2  gate2061(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2062(.a(s_216), .O(gate421inter3));
  inv1  gate2063(.a(s_217), .O(gate421inter4));
  nand2 gate2064(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2065(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2066(.a(G2), .O(gate421inter7));
  inv1  gate2067(.a(G1135), .O(gate421inter8));
  nand2 gate2068(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2069(.a(s_217), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2070(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2071(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2072(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate1961(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1962(.a(gate422inter0), .b(s_202), .O(gate422inter1));
  and2  gate1963(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1964(.a(s_202), .O(gate422inter3));
  inv1  gate1965(.a(s_203), .O(gate422inter4));
  nand2 gate1966(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1967(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1968(.a(G1039), .O(gate422inter7));
  inv1  gate1969(.a(G1135), .O(gate422inter8));
  nand2 gate1970(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1971(.a(s_203), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1972(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1973(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1974(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1289(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1290(.a(gate423inter0), .b(s_106), .O(gate423inter1));
  and2  gate1291(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1292(.a(s_106), .O(gate423inter3));
  inv1  gate1293(.a(s_107), .O(gate423inter4));
  nand2 gate1294(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1295(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1296(.a(G3), .O(gate423inter7));
  inv1  gate1297(.a(G1138), .O(gate423inter8));
  nand2 gate1298(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1299(.a(s_107), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1300(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1301(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1302(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate2843(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2844(.a(gate424inter0), .b(s_328), .O(gate424inter1));
  and2  gate2845(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2846(.a(s_328), .O(gate424inter3));
  inv1  gate2847(.a(s_329), .O(gate424inter4));
  nand2 gate2848(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2849(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2850(.a(G1042), .O(gate424inter7));
  inv1  gate2851(.a(G1138), .O(gate424inter8));
  nand2 gate2852(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2853(.a(s_329), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2854(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2855(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2856(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate2829(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2830(.a(gate425inter0), .b(s_326), .O(gate425inter1));
  and2  gate2831(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2832(.a(s_326), .O(gate425inter3));
  inv1  gate2833(.a(s_327), .O(gate425inter4));
  nand2 gate2834(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2835(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2836(.a(G4), .O(gate425inter7));
  inv1  gate2837(.a(G1141), .O(gate425inter8));
  nand2 gate2838(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2839(.a(s_327), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2840(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2841(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2842(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate701(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate702(.a(gate427inter0), .b(s_22), .O(gate427inter1));
  and2  gate703(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate704(.a(s_22), .O(gate427inter3));
  inv1  gate705(.a(s_23), .O(gate427inter4));
  nand2 gate706(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate707(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate708(.a(G5), .O(gate427inter7));
  inv1  gate709(.a(G1144), .O(gate427inter8));
  nand2 gate710(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate711(.a(s_23), .b(gate427inter3), .O(gate427inter10));
  nor2  gate712(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate713(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate714(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2619(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2620(.a(gate430inter0), .b(s_296), .O(gate430inter1));
  and2  gate2621(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2622(.a(s_296), .O(gate430inter3));
  inv1  gate2623(.a(s_297), .O(gate430inter4));
  nand2 gate2624(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2625(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2626(.a(G1051), .O(gate430inter7));
  inv1  gate2627(.a(G1147), .O(gate430inter8));
  nand2 gate2628(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2629(.a(s_297), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2630(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2631(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2632(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate911(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate912(.a(gate433inter0), .b(s_52), .O(gate433inter1));
  and2  gate913(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate914(.a(s_52), .O(gate433inter3));
  inv1  gate915(.a(s_53), .O(gate433inter4));
  nand2 gate916(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate917(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate918(.a(G8), .O(gate433inter7));
  inv1  gate919(.a(G1153), .O(gate433inter8));
  nand2 gate920(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate921(.a(s_53), .b(gate433inter3), .O(gate433inter10));
  nor2  gate922(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate923(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate924(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate3109(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate3110(.a(gate434inter0), .b(s_366), .O(gate434inter1));
  and2  gate3111(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate3112(.a(s_366), .O(gate434inter3));
  inv1  gate3113(.a(s_367), .O(gate434inter4));
  nand2 gate3114(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate3115(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate3116(.a(G1057), .O(gate434inter7));
  inv1  gate3117(.a(G1153), .O(gate434inter8));
  nand2 gate3118(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate3119(.a(s_367), .b(gate434inter3), .O(gate434inter10));
  nor2  gate3120(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate3121(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate3122(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1877(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1878(.a(gate435inter0), .b(s_190), .O(gate435inter1));
  and2  gate1879(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1880(.a(s_190), .O(gate435inter3));
  inv1  gate1881(.a(s_191), .O(gate435inter4));
  nand2 gate1882(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1883(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1884(.a(G9), .O(gate435inter7));
  inv1  gate1885(.a(G1156), .O(gate435inter8));
  nand2 gate1886(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1887(.a(s_191), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1888(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1889(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1890(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate925(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate926(.a(gate436inter0), .b(s_54), .O(gate436inter1));
  and2  gate927(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate928(.a(s_54), .O(gate436inter3));
  inv1  gate929(.a(s_55), .O(gate436inter4));
  nand2 gate930(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate931(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate932(.a(G1060), .O(gate436inter7));
  inv1  gate933(.a(G1156), .O(gate436inter8));
  nand2 gate934(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate935(.a(s_55), .b(gate436inter3), .O(gate436inter10));
  nor2  gate936(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate937(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate938(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate2003(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2004(.a(gate437inter0), .b(s_208), .O(gate437inter1));
  and2  gate2005(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2006(.a(s_208), .O(gate437inter3));
  inv1  gate2007(.a(s_209), .O(gate437inter4));
  nand2 gate2008(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2009(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2010(.a(G10), .O(gate437inter7));
  inv1  gate2011(.a(G1159), .O(gate437inter8));
  nand2 gate2012(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2013(.a(s_209), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2014(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2015(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2016(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1359(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1360(.a(gate438inter0), .b(s_116), .O(gate438inter1));
  and2  gate1361(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1362(.a(s_116), .O(gate438inter3));
  inv1  gate1363(.a(s_117), .O(gate438inter4));
  nand2 gate1364(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1365(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1366(.a(G1063), .O(gate438inter7));
  inv1  gate1367(.a(G1159), .O(gate438inter8));
  nand2 gate1368(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1369(.a(s_117), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1370(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1371(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1372(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate3277(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate3278(.a(gate439inter0), .b(s_390), .O(gate439inter1));
  and2  gate3279(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate3280(.a(s_390), .O(gate439inter3));
  inv1  gate3281(.a(s_391), .O(gate439inter4));
  nand2 gate3282(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate3283(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate3284(.a(G11), .O(gate439inter7));
  inv1  gate3285(.a(G1162), .O(gate439inter8));
  nand2 gate3286(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate3287(.a(s_391), .b(gate439inter3), .O(gate439inter10));
  nor2  gate3288(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate3289(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate3290(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate2031(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2032(.a(gate440inter0), .b(s_212), .O(gate440inter1));
  and2  gate2033(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2034(.a(s_212), .O(gate440inter3));
  inv1  gate2035(.a(s_213), .O(gate440inter4));
  nand2 gate2036(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2037(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2038(.a(G1066), .O(gate440inter7));
  inv1  gate2039(.a(G1162), .O(gate440inter8));
  nand2 gate2040(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2041(.a(s_213), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2042(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2043(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2044(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1233(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1234(.a(gate443inter0), .b(s_98), .O(gate443inter1));
  and2  gate1235(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1236(.a(s_98), .O(gate443inter3));
  inv1  gate1237(.a(s_99), .O(gate443inter4));
  nand2 gate1238(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1239(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1240(.a(G13), .O(gate443inter7));
  inv1  gate1241(.a(G1168), .O(gate443inter8));
  nand2 gate1242(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1243(.a(s_99), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1244(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1245(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1246(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1569(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1570(.a(gate445inter0), .b(s_146), .O(gate445inter1));
  and2  gate1571(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1572(.a(s_146), .O(gate445inter3));
  inv1  gate1573(.a(s_147), .O(gate445inter4));
  nand2 gate1574(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1575(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1576(.a(G14), .O(gate445inter7));
  inv1  gate1577(.a(G1171), .O(gate445inter8));
  nand2 gate1578(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1579(.a(s_147), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1580(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1581(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1582(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate2507(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2508(.a(gate447inter0), .b(s_280), .O(gate447inter1));
  and2  gate2509(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2510(.a(s_280), .O(gate447inter3));
  inv1  gate2511(.a(s_281), .O(gate447inter4));
  nand2 gate2512(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2513(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2514(.a(G15), .O(gate447inter7));
  inv1  gate2515(.a(G1174), .O(gate447inter8));
  nand2 gate2516(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2517(.a(s_281), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2518(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2519(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2520(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1527(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1528(.a(gate448inter0), .b(s_140), .O(gate448inter1));
  and2  gate1529(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1530(.a(s_140), .O(gate448inter3));
  inv1  gate1531(.a(s_141), .O(gate448inter4));
  nand2 gate1532(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1533(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1534(.a(G1078), .O(gate448inter7));
  inv1  gate1535(.a(G1174), .O(gate448inter8));
  nand2 gate1536(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1537(.a(s_141), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1538(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1539(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1540(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2395(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2396(.a(gate451inter0), .b(s_264), .O(gate451inter1));
  and2  gate2397(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2398(.a(s_264), .O(gate451inter3));
  inv1  gate2399(.a(s_265), .O(gate451inter4));
  nand2 gate2400(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2401(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2402(.a(G17), .O(gate451inter7));
  inv1  gate2403(.a(G1180), .O(gate451inter8));
  nand2 gate2404(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2405(.a(s_265), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2406(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2407(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2408(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate2535(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate2536(.a(gate454inter0), .b(s_284), .O(gate454inter1));
  and2  gate2537(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate2538(.a(s_284), .O(gate454inter3));
  inv1  gate2539(.a(s_285), .O(gate454inter4));
  nand2 gate2540(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate2541(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate2542(.a(G1087), .O(gate454inter7));
  inv1  gate2543(.a(G1183), .O(gate454inter8));
  nand2 gate2544(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate2545(.a(s_285), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2546(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2547(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2548(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1219(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1220(.a(gate455inter0), .b(s_96), .O(gate455inter1));
  and2  gate1221(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1222(.a(s_96), .O(gate455inter3));
  inv1  gate1223(.a(s_97), .O(gate455inter4));
  nand2 gate1224(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1225(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1226(.a(G19), .O(gate455inter7));
  inv1  gate1227(.a(G1186), .O(gate455inter8));
  nand2 gate1228(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1229(.a(s_97), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1230(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1231(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1232(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1079(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1080(.a(gate456inter0), .b(s_76), .O(gate456inter1));
  and2  gate1081(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1082(.a(s_76), .O(gate456inter3));
  inv1  gate1083(.a(s_77), .O(gate456inter4));
  nand2 gate1084(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1085(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1086(.a(G1090), .O(gate456inter7));
  inv1  gate1087(.a(G1186), .O(gate456inter8));
  nand2 gate1088(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1089(.a(s_77), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1090(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1091(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1092(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate2731(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2732(.a(gate457inter0), .b(s_312), .O(gate457inter1));
  and2  gate2733(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2734(.a(s_312), .O(gate457inter3));
  inv1  gate2735(.a(s_313), .O(gate457inter4));
  nand2 gate2736(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2737(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2738(.a(G20), .O(gate457inter7));
  inv1  gate2739(.a(G1189), .O(gate457inter8));
  nand2 gate2740(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2741(.a(s_313), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2742(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2743(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2744(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1555(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1556(.a(gate464inter0), .b(s_144), .O(gate464inter1));
  and2  gate1557(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1558(.a(s_144), .O(gate464inter3));
  inv1  gate1559(.a(s_145), .O(gate464inter4));
  nand2 gate1560(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1561(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1562(.a(G1102), .O(gate464inter7));
  inv1  gate1563(.a(G1198), .O(gate464inter8));
  nand2 gate1564(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1565(.a(s_145), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1566(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1567(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1568(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate995(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate996(.a(gate466inter0), .b(s_64), .O(gate466inter1));
  and2  gate997(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate998(.a(s_64), .O(gate466inter3));
  inv1  gate999(.a(s_65), .O(gate466inter4));
  nand2 gate1000(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1001(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1002(.a(G1105), .O(gate466inter7));
  inv1  gate1003(.a(G1201), .O(gate466inter8));
  nand2 gate1004(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1005(.a(s_65), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1006(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1007(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1008(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1177(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1178(.a(gate467inter0), .b(s_90), .O(gate467inter1));
  and2  gate1179(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1180(.a(s_90), .O(gate467inter3));
  inv1  gate1181(.a(s_91), .O(gate467inter4));
  nand2 gate1182(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1183(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1184(.a(G25), .O(gate467inter7));
  inv1  gate1185(.a(G1204), .O(gate467inter8));
  nand2 gate1186(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1187(.a(s_91), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1188(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1189(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1190(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2955(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2956(.a(gate470inter0), .b(s_344), .O(gate470inter1));
  and2  gate2957(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2958(.a(s_344), .O(gate470inter3));
  inv1  gate2959(.a(s_345), .O(gate470inter4));
  nand2 gate2960(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2961(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2962(.a(G1111), .O(gate470inter7));
  inv1  gate2963(.a(G1207), .O(gate470inter8));
  nand2 gate2964(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2965(.a(s_345), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2966(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2967(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2968(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2409(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2410(.a(gate475inter0), .b(s_266), .O(gate475inter1));
  and2  gate2411(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2412(.a(s_266), .O(gate475inter3));
  inv1  gate2413(.a(s_267), .O(gate475inter4));
  nand2 gate2414(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2415(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2416(.a(G29), .O(gate475inter7));
  inv1  gate2417(.a(G1216), .O(gate475inter8));
  nand2 gate2418(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2419(.a(s_267), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2420(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2421(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2422(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1807(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1808(.a(gate476inter0), .b(s_180), .O(gate476inter1));
  and2  gate1809(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1810(.a(s_180), .O(gate476inter3));
  inv1  gate1811(.a(s_181), .O(gate476inter4));
  nand2 gate1812(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1813(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1814(.a(G1120), .O(gate476inter7));
  inv1  gate1815(.a(G1216), .O(gate476inter8));
  nand2 gate1816(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1817(.a(s_181), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1818(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1819(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1820(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate589(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate590(.a(gate478inter0), .b(s_6), .O(gate478inter1));
  and2  gate591(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate592(.a(s_6), .O(gate478inter3));
  inv1  gate593(.a(s_7), .O(gate478inter4));
  nand2 gate594(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate595(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate596(.a(G1123), .O(gate478inter7));
  inv1  gate597(.a(G1219), .O(gate478inter8));
  nand2 gate598(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate599(.a(s_7), .b(gate478inter3), .O(gate478inter10));
  nor2  gate600(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate601(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate602(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2745(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2746(.a(gate479inter0), .b(s_314), .O(gate479inter1));
  and2  gate2747(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2748(.a(s_314), .O(gate479inter3));
  inv1  gate2749(.a(s_315), .O(gate479inter4));
  nand2 gate2750(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2751(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2752(.a(G31), .O(gate479inter7));
  inv1  gate2753(.a(G1222), .O(gate479inter8));
  nand2 gate2754(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2755(.a(s_315), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2756(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2757(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2758(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate2577(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2578(.a(gate481inter0), .b(s_290), .O(gate481inter1));
  and2  gate2579(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2580(.a(s_290), .O(gate481inter3));
  inv1  gate2581(.a(s_291), .O(gate481inter4));
  nand2 gate2582(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2583(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2584(.a(G32), .O(gate481inter7));
  inv1  gate2585(.a(G1225), .O(gate481inter8));
  nand2 gate2586(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2587(.a(s_291), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2588(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2589(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2590(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2199(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2200(.a(gate486inter0), .b(s_236), .O(gate486inter1));
  and2  gate2201(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2202(.a(s_236), .O(gate486inter3));
  inv1  gate2203(.a(s_237), .O(gate486inter4));
  nand2 gate2204(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2205(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2206(.a(G1234), .O(gate486inter7));
  inv1  gate2207(.a(G1235), .O(gate486inter8));
  nand2 gate2208(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2209(.a(s_237), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2210(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2211(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2212(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate953(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate954(.a(gate489inter0), .b(s_58), .O(gate489inter1));
  and2  gate955(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate956(.a(s_58), .O(gate489inter3));
  inv1  gate957(.a(s_59), .O(gate489inter4));
  nand2 gate958(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate959(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate960(.a(G1240), .O(gate489inter7));
  inv1  gate961(.a(G1241), .O(gate489inter8));
  nand2 gate962(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate963(.a(s_59), .b(gate489inter3), .O(gate489inter10));
  nor2  gate964(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate965(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate966(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1667(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1668(.a(gate491inter0), .b(s_160), .O(gate491inter1));
  and2  gate1669(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1670(.a(s_160), .O(gate491inter3));
  inv1  gate1671(.a(s_161), .O(gate491inter4));
  nand2 gate1672(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1673(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1674(.a(G1244), .O(gate491inter7));
  inv1  gate1675(.a(G1245), .O(gate491inter8));
  nand2 gate1676(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1677(.a(s_161), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1678(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1679(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1680(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2941(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2942(.a(gate493inter0), .b(s_342), .O(gate493inter1));
  and2  gate2943(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2944(.a(s_342), .O(gate493inter3));
  inv1  gate2945(.a(s_343), .O(gate493inter4));
  nand2 gate2946(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2947(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2948(.a(G1248), .O(gate493inter7));
  inv1  gate2949(.a(G1249), .O(gate493inter8));
  nand2 gate2950(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2951(.a(s_343), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2952(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2953(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2954(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate2717(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2718(.a(gate494inter0), .b(s_310), .O(gate494inter1));
  and2  gate2719(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2720(.a(s_310), .O(gate494inter3));
  inv1  gate2721(.a(s_311), .O(gate494inter4));
  nand2 gate2722(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2723(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2724(.a(G1250), .O(gate494inter7));
  inv1  gate2725(.a(G1251), .O(gate494inter8));
  nand2 gate2726(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2727(.a(s_311), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2728(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2729(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2730(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate897(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate898(.a(gate502inter0), .b(s_50), .O(gate502inter1));
  and2  gate899(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate900(.a(s_50), .O(gate502inter3));
  inv1  gate901(.a(s_51), .O(gate502inter4));
  nand2 gate902(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate903(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate904(.a(G1266), .O(gate502inter7));
  inv1  gate905(.a(G1267), .O(gate502inter8));
  nand2 gate906(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate907(.a(s_51), .b(gate502inter3), .O(gate502inter10));
  nor2  gate908(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate909(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate910(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate3193(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate3194(.a(gate505inter0), .b(s_378), .O(gate505inter1));
  and2  gate3195(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate3196(.a(s_378), .O(gate505inter3));
  inv1  gate3197(.a(s_379), .O(gate505inter4));
  nand2 gate3198(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate3199(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate3200(.a(G1272), .O(gate505inter7));
  inv1  gate3201(.a(G1273), .O(gate505inter8));
  nand2 gate3202(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate3203(.a(s_379), .b(gate505inter3), .O(gate505inter10));
  nor2  gate3204(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate3205(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate3206(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate2815(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate2816(.a(gate506inter0), .b(s_324), .O(gate506inter1));
  and2  gate2817(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate2818(.a(s_324), .O(gate506inter3));
  inv1  gate2819(.a(s_325), .O(gate506inter4));
  nand2 gate2820(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate2821(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate2822(.a(G1274), .O(gate506inter7));
  inv1  gate2823(.a(G1275), .O(gate506inter8));
  nand2 gate2824(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate2825(.a(s_325), .b(gate506inter3), .O(gate506inter10));
  nor2  gate2826(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate2827(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate2828(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1499(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1500(.a(gate509inter0), .b(s_136), .O(gate509inter1));
  and2  gate1501(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1502(.a(s_136), .O(gate509inter3));
  inv1  gate1503(.a(s_137), .O(gate509inter4));
  nand2 gate1504(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1505(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1506(.a(G1280), .O(gate509inter7));
  inv1  gate1507(.a(G1281), .O(gate509inter8));
  nand2 gate1508(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1509(.a(s_137), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1510(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1511(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1512(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate3123(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate3124(.a(gate510inter0), .b(s_368), .O(gate510inter1));
  and2  gate3125(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate3126(.a(s_368), .O(gate510inter3));
  inv1  gate3127(.a(s_369), .O(gate510inter4));
  nand2 gate3128(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate3129(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate3130(.a(G1282), .O(gate510inter7));
  inv1  gate3131(.a(G1283), .O(gate510inter8));
  nand2 gate3132(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate3133(.a(s_369), .b(gate510inter3), .O(gate510inter10));
  nor2  gate3134(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate3135(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate3136(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule