module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2717(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2718(.a(gate13inter0), .b(s_310), .O(gate13inter1));
  and2  gate2719(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2720(.a(s_310), .O(gate13inter3));
  inv1  gate2721(.a(s_311), .O(gate13inter4));
  nand2 gate2722(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2723(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2724(.a(G9), .O(gate13inter7));
  inv1  gate2725(.a(G10), .O(gate13inter8));
  nand2 gate2726(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2727(.a(s_311), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2728(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2729(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2730(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1751(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1752(.a(gate20inter0), .b(s_172), .O(gate20inter1));
  and2  gate1753(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1754(.a(s_172), .O(gate20inter3));
  inv1  gate1755(.a(s_173), .O(gate20inter4));
  nand2 gate1756(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1757(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1758(.a(G23), .O(gate20inter7));
  inv1  gate1759(.a(G24), .O(gate20inter8));
  nand2 gate1760(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1761(.a(s_173), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1762(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1763(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1764(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1933(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1934(.a(gate22inter0), .b(s_198), .O(gate22inter1));
  and2  gate1935(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1936(.a(s_198), .O(gate22inter3));
  inv1  gate1937(.a(s_199), .O(gate22inter4));
  nand2 gate1938(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1939(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1940(.a(G27), .O(gate22inter7));
  inv1  gate1941(.a(G28), .O(gate22inter8));
  nand2 gate1942(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1943(.a(s_199), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1944(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1945(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1946(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1065(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1066(.a(gate23inter0), .b(s_74), .O(gate23inter1));
  and2  gate1067(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1068(.a(s_74), .O(gate23inter3));
  inv1  gate1069(.a(s_75), .O(gate23inter4));
  nand2 gate1070(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1071(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1072(.a(G29), .O(gate23inter7));
  inv1  gate1073(.a(G30), .O(gate23inter8));
  nand2 gate1074(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1075(.a(s_75), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1076(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1077(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1078(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1975(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1976(.a(gate24inter0), .b(s_204), .O(gate24inter1));
  and2  gate1977(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1978(.a(s_204), .O(gate24inter3));
  inv1  gate1979(.a(s_205), .O(gate24inter4));
  nand2 gate1980(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1981(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1982(.a(G31), .O(gate24inter7));
  inv1  gate1983(.a(G32), .O(gate24inter8));
  nand2 gate1984(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1985(.a(s_205), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1986(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1987(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1988(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1247(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1248(.a(gate25inter0), .b(s_100), .O(gate25inter1));
  and2  gate1249(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1250(.a(s_100), .O(gate25inter3));
  inv1  gate1251(.a(s_101), .O(gate25inter4));
  nand2 gate1252(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1253(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1254(.a(G1), .O(gate25inter7));
  inv1  gate1255(.a(G5), .O(gate25inter8));
  nand2 gate1256(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1257(.a(s_101), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1258(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1259(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1260(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate2801(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2802(.a(gate26inter0), .b(s_322), .O(gate26inter1));
  and2  gate2803(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2804(.a(s_322), .O(gate26inter3));
  inv1  gate2805(.a(s_323), .O(gate26inter4));
  nand2 gate2806(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2807(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2808(.a(G9), .O(gate26inter7));
  inv1  gate2809(.a(G13), .O(gate26inter8));
  nand2 gate2810(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2811(.a(s_323), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2812(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2813(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2814(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2885(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2886(.a(gate29inter0), .b(s_334), .O(gate29inter1));
  and2  gate2887(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2888(.a(s_334), .O(gate29inter3));
  inv1  gate2889(.a(s_335), .O(gate29inter4));
  nand2 gate2890(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2891(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2892(.a(G3), .O(gate29inter7));
  inv1  gate2893(.a(G7), .O(gate29inter8));
  nand2 gate2894(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2895(.a(s_335), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2896(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2897(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2898(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate939(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate940(.a(gate30inter0), .b(s_56), .O(gate30inter1));
  and2  gate941(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate942(.a(s_56), .O(gate30inter3));
  inv1  gate943(.a(s_57), .O(gate30inter4));
  nand2 gate944(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate945(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate946(.a(G11), .O(gate30inter7));
  inv1  gate947(.a(G15), .O(gate30inter8));
  nand2 gate948(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate949(.a(s_57), .b(gate30inter3), .O(gate30inter10));
  nor2  gate950(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate951(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate952(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1359(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1360(.a(gate32inter0), .b(s_116), .O(gate32inter1));
  and2  gate1361(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1362(.a(s_116), .O(gate32inter3));
  inv1  gate1363(.a(s_117), .O(gate32inter4));
  nand2 gate1364(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1365(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1366(.a(G12), .O(gate32inter7));
  inv1  gate1367(.a(G16), .O(gate32inter8));
  nand2 gate1368(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1369(.a(s_117), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1370(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1371(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1372(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate2549(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2550(.a(gate33inter0), .b(s_286), .O(gate33inter1));
  and2  gate2551(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2552(.a(s_286), .O(gate33inter3));
  inv1  gate2553(.a(s_287), .O(gate33inter4));
  nand2 gate2554(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2555(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2556(.a(G17), .O(gate33inter7));
  inv1  gate2557(.a(G21), .O(gate33inter8));
  nand2 gate2558(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2559(.a(s_287), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2560(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2561(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2562(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1093(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1094(.a(gate35inter0), .b(s_78), .O(gate35inter1));
  and2  gate1095(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1096(.a(s_78), .O(gate35inter3));
  inv1  gate1097(.a(s_79), .O(gate35inter4));
  nand2 gate1098(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1099(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1100(.a(G18), .O(gate35inter7));
  inv1  gate1101(.a(G22), .O(gate35inter8));
  nand2 gate1102(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1103(.a(s_79), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1104(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1105(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1106(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1485(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1486(.a(gate38inter0), .b(s_134), .O(gate38inter1));
  and2  gate1487(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1488(.a(s_134), .O(gate38inter3));
  inv1  gate1489(.a(s_135), .O(gate38inter4));
  nand2 gate1490(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1491(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1492(.a(G27), .O(gate38inter7));
  inv1  gate1493(.a(G31), .O(gate38inter8));
  nand2 gate1494(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1495(.a(s_135), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1496(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1497(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1498(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate3137(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate3138(.a(gate39inter0), .b(s_370), .O(gate39inter1));
  and2  gate3139(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate3140(.a(s_370), .O(gate39inter3));
  inv1  gate3141(.a(s_371), .O(gate39inter4));
  nand2 gate3142(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate3143(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate3144(.a(G20), .O(gate39inter7));
  inv1  gate3145(.a(G24), .O(gate39inter8));
  nand2 gate3146(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate3147(.a(s_371), .b(gate39inter3), .O(gate39inter10));
  nor2  gate3148(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate3149(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate3150(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1821(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1822(.a(gate41inter0), .b(s_182), .O(gate41inter1));
  and2  gate1823(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1824(.a(s_182), .O(gate41inter3));
  inv1  gate1825(.a(s_183), .O(gate41inter4));
  nand2 gate1826(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1827(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1828(.a(G1), .O(gate41inter7));
  inv1  gate1829(.a(G266), .O(gate41inter8));
  nand2 gate1830(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1831(.a(s_183), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1832(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1833(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1834(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1611(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1612(.a(gate42inter0), .b(s_152), .O(gate42inter1));
  and2  gate1613(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1614(.a(s_152), .O(gate42inter3));
  inv1  gate1615(.a(s_153), .O(gate42inter4));
  nand2 gate1616(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1617(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1618(.a(G2), .O(gate42inter7));
  inv1  gate1619(.a(G266), .O(gate42inter8));
  nand2 gate1620(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1621(.a(s_153), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1622(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1623(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1624(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1989(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1990(.a(gate45inter0), .b(s_206), .O(gate45inter1));
  and2  gate1991(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1992(.a(s_206), .O(gate45inter3));
  inv1  gate1993(.a(s_207), .O(gate45inter4));
  nand2 gate1994(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1995(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1996(.a(G5), .O(gate45inter7));
  inv1  gate1997(.a(G272), .O(gate45inter8));
  nand2 gate1998(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1999(.a(s_207), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2000(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2001(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2002(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2003(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2004(.a(gate47inter0), .b(s_208), .O(gate47inter1));
  and2  gate2005(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2006(.a(s_208), .O(gate47inter3));
  inv1  gate2007(.a(s_209), .O(gate47inter4));
  nand2 gate2008(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2009(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2010(.a(G7), .O(gate47inter7));
  inv1  gate2011(.a(G275), .O(gate47inter8));
  nand2 gate2012(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2013(.a(s_209), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2014(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2015(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2016(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1555(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1556(.a(gate48inter0), .b(s_144), .O(gate48inter1));
  and2  gate1557(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1558(.a(s_144), .O(gate48inter3));
  inv1  gate1559(.a(s_145), .O(gate48inter4));
  nand2 gate1560(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1561(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1562(.a(G8), .O(gate48inter7));
  inv1  gate1563(.a(G275), .O(gate48inter8));
  nand2 gate1564(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1565(.a(s_145), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1566(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1567(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1568(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2563(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2564(.a(gate50inter0), .b(s_288), .O(gate50inter1));
  and2  gate2565(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2566(.a(s_288), .O(gate50inter3));
  inv1  gate2567(.a(s_289), .O(gate50inter4));
  nand2 gate2568(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2569(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2570(.a(G10), .O(gate50inter7));
  inv1  gate2571(.a(G278), .O(gate50inter8));
  nand2 gate2572(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2573(.a(s_289), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2574(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2575(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2576(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1023(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1024(.a(gate51inter0), .b(s_68), .O(gate51inter1));
  and2  gate1025(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1026(.a(s_68), .O(gate51inter3));
  inv1  gate1027(.a(s_69), .O(gate51inter4));
  nand2 gate1028(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1029(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1030(.a(G11), .O(gate51inter7));
  inv1  gate1031(.a(G281), .O(gate51inter8));
  nand2 gate1032(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1033(.a(s_69), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1034(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1035(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1036(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1079(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1080(.a(gate56inter0), .b(s_76), .O(gate56inter1));
  and2  gate1081(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1082(.a(s_76), .O(gate56inter3));
  inv1  gate1083(.a(s_77), .O(gate56inter4));
  nand2 gate1084(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1085(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1086(.a(G16), .O(gate56inter7));
  inv1  gate1087(.a(G287), .O(gate56inter8));
  nand2 gate1088(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1089(.a(s_77), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1090(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1091(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1092(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2325(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2326(.a(gate66inter0), .b(s_254), .O(gate66inter1));
  and2  gate2327(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2328(.a(s_254), .O(gate66inter3));
  inv1  gate2329(.a(s_255), .O(gate66inter4));
  nand2 gate2330(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2331(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2332(.a(G26), .O(gate66inter7));
  inv1  gate2333(.a(G302), .O(gate66inter8));
  nand2 gate2334(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2335(.a(s_255), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2336(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2337(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2338(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate981(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate982(.a(gate69inter0), .b(s_62), .O(gate69inter1));
  and2  gate983(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate984(.a(s_62), .O(gate69inter3));
  inv1  gate985(.a(s_63), .O(gate69inter4));
  nand2 gate986(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate987(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate988(.a(G29), .O(gate69inter7));
  inv1  gate989(.a(G308), .O(gate69inter8));
  nand2 gate990(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate991(.a(s_63), .b(gate69inter3), .O(gate69inter10));
  nor2  gate992(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate993(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate994(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate2857(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate2858(.a(gate71inter0), .b(s_330), .O(gate71inter1));
  and2  gate2859(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate2860(.a(s_330), .O(gate71inter3));
  inv1  gate2861(.a(s_331), .O(gate71inter4));
  nand2 gate2862(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate2863(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate2864(.a(G31), .O(gate71inter7));
  inv1  gate2865(.a(G311), .O(gate71inter8));
  nand2 gate2866(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate2867(.a(s_331), .b(gate71inter3), .O(gate71inter10));
  nor2  gate2868(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate2869(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate2870(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate2927(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2928(.a(gate75inter0), .b(s_340), .O(gate75inter1));
  and2  gate2929(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2930(.a(s_340), .O(gate75inter3));
  inv1  gate2931(.a(s_341), .O(gate75inter4));
  nand2 gate2932(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2933(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2934(.a(G9), .O(gate75inter7));
  inv1  gate2935(.a(G317), .O(gate75inter8));
  nand2 gate2936(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2937(.a(s_341), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2938(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2939(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2940(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate2185(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2186(.a(gate76inter0), .b(s_234), .O(gate76inter1));
  and2  gate2187(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2188(.a(s_234), .O(gate76inter3));
  inv1  gate2189(.a(s_235), .O(gate76inter4));
  nand2 gate2190(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2191(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2192(.a(G13), .O(gate76inter7));
  inv1  gate2193(.a(G317), .O(gate76inter8));
  nand2 gate2194(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2195(.a(s_235), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2196(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2197(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2198(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate2101(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2102(.a(gate77inter0), .b(s_222), .O(gate77inter1));
  and2  gate2103(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2104(.a(s_222), .O(gate77inter3));
  inv1  gate2105(.a(s_223), .O(gate77inter4));
  nand2 gate2106(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2107(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2108(.a(G2), .O(gate77inter7));
  inv1  gate2109(.a(G320), .O(gate77inter8));
  nand2 gate2110(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2111(.a(s_223), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2112(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2113(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2114(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate1681(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate1682(.a(gate78inter0), .b(s_162), .O(gate78inter1));
  and2  gate1683(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate1684(.a(s_162), .O(gate78inter3));
  inv1  gate1685(.a(s_163), .O(gate78inter4));
  nand2 gate1686(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate1687(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate1688(.a(G6), .O(gate78inter7));
  inv1  gate1689(.a(G320), .O(gate78inter8));
  nand2 gate1690(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate1691(.a(s_163), .b(gate78inter3), .O(gate78inter10));
  nor2  gate1692(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate1693(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate1694(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate645(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate646(.a(gate79inter0), .b(s_14), .O(gate79inter1));
  and2  gate647(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate648(.a(s_14), .O(gate79inter3));
  inv1  gate649(.a(s_15), .O(gate79inter4));
  nand2 gate650(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate651(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate652(.a(G10), .O(gate79inter7));
  inv1  gate653(.a(G323), .O(gate79inter8));
  nand2 gate654(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate655(.a(s_15), .b(gate79inter3), .O(gate79inter10));
  nor2  gate656(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate657(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate658(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate2731(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2732(.a(gate80inter0), .b(s_312), .O(gate80inter1));
  and2  gate2733(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2734(.a(s_312), .O(gate80inter3));
  inv1  gate2735(.a(s_313), .O(gate80inter4));
  nand2 gate2736(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2737(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2738(.a(G14), .O(gate80inter7));
  inv1  gate2739(.a(G323), .O(gate80inter8));
  nand2 gate2740(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2741(.a(s_313), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2742(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2743(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2744(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1625(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1626(.a(gate81inter0), .b(s_154), .O(gate81inter1));
  and2  gate1627(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1628(.a(s_154), .O(gate81inter3));
  inv1  gate1629(.a(s_155), .O(gate81inter4));
  nand2 gate1630(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1631(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1632(.a(G3), .O(gate81inter7));
  inv1  gate1633(.a(G326), .O(gate81inter8));
  nand2 gate1634(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1635(.a(s_155), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1636(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1637(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1638(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1723(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1724(.a(gate83inter0), .b(s_168), .O(gate83inter1));
  and2  gate1725(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1726(.a(s_168), .O(gate83inter3));
  inv1  gate1727(.a(s_169), .O(gate83inter4));
  nand2 gate1728(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1729(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1730(.a(G11), .O(gate83inter7));
  inv1  gate1731(.a(G329), .O(gate83inter8));
  nand2 gate1732(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1733(.a(s_169), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1734(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1735(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1736(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate687(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate688(.a(gate86inter0), .b(s_20), .O(gate86inter1));
  and2  gate689(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate690(.a(s_20), .O(gate86inter3));
  inv1  gate691(.a(s_21), .O(gate86inter4));
  nand2 gate692(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate693(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate694(.a(G8), .O(gate86inter7));
  inv1  gate695(.a(G332), .O(gate86inter8));
  nand2 gate696(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate697(.a(s_21), .b(gate86inter3), .O(gate86inter10));
  nor2  gate698(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate699(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate700(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate841(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate842(.a(gate88inter0), .b(s_42), .O(gate88inter1));
  and2  gate843(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate844(.a(s_42), .O(gate88inter3));
  inv1  gate845(.a(s_43), .O(gate88inter4));
  nand2 gate846(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate847(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate848(.a(G16), .O(gate88inter7));
  inv1  gate849(.a(G335), .O(gate88inter8));
  nand2 gate850(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate851(.a(s_43), .b(gate88inter3), .O(gate88inter10));
  nor2  gate852(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate853(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate854(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1541(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1542(.a(gate91inter0), .b(s_142), .O(gate91inter1));
  and2  gate1543(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1544(.a(s_142), .O(gate91inter3));
  inv1  gate1545(.a(s_143), .O(gate91inter4));
  nand2 gate1546(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1547(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1548(.a(G25), .O(gate91inter7));
  inv1  gate1549(.a(G341), .O(gate91inter8));
  nand2 gate1550(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1551(.a(s_143), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1552(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1553(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1554(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2983(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2984(.a(gate92inter0), .b(s_348), .O(gate92inter1));
  and2  gate2985(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2986(.a(s_348), .O(gate92inter3));
  inv1  gate2987(.a(s_349), .O(gate92inter4));
  nand2 gate2988(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2989(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2990(.a(G29), .O(gate92inter7));
  inv1  gate2991(.a(G341), .O(gate92inter8));
  nand2 gate2992(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2993(.a(s_349), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2994(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2995(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2996(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate729(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate730(.a(gate93inter0), .b(s_26), .O(gate93inter1));
  and2  gate731(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate732(.a(s_26), .O(gate93inter3));
  inv1  gate733(.a(s_27), .O(gate93inter4));
  nand2 gate734(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate735(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate736(.a(G18), .O(gate93inter7));
  inv1  gate737(.a(G344), .O(gate93inter8));
  nand2 gate738(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate739(.a(s_27), .b(gate93inter3), .O(gate93inter10));
  nor2  gate740(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate741(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate742(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate855(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate856(.a(gate95inter0), .b(s_44), .O(gate95inter1));
  and2  gate857(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate858(.a(s_44), .O(gate95inter3));
  inv1  gate859(.a(s_45), .O(gate95inter4));
  nand2 gate860(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate861(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate862(.a(G26), .O(gate95inter7));
  inv1  gate863(.a(G347), .O(gate95inter8));
  nand2 gate864(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate865(.a(s_45), .b(gate95inter3), .O(gate95inter10));
  nor2  gate866(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate867(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate868(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2157(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2158(.a(gate105inter0), .b(s_230), .O(gate105inter1));
  and2  gate2159(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2160(.a(s_230), .O(gate105inter3));
  inv1  gate2161(.a(s_231), .O(gate105inter4));
  nand2 gate2162(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2163(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2164(.a(G362), .O(gate105inter7));
  inv1  gate2165(.a(G363), .O(gate105inter8));
  nand2 gate2166(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2167(.a(s_231), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2168(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2169(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2170(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1863(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1864(.a(gate108inter0), .b(s_188), .O(gate108inter1));
  and2  gate1865(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1866(.a(s_188), .O(gate108inter3));
  inv1  gate1867(.a(s_189), .O(gate108inter4));
  nand2 gate1868(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1869(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1870(.a(G368), .O(gate108inter7));
  inv1  gate1871(.a(G369), .O(gate108inter8));
  nand2 gate1872(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1873(.a(s_189), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1874(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1875(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1876(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate953(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate954(.a(gate109inter0), .b(s_58), .O(gate109inter1));
  and2  gate955(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate956(.a(s_58), .O(gate109inter3));
  inv1  gate957(.a(s_59), .O(gate109inter4));
  nand2 gate958(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate959(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate960(.a(G370), .O(gate109inter7));
  inv1  gate961(.a(G371), .O(gate109inter8));
  nand2 gate962(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate963(.a(s_59), .b(gate109inter3), .O(gate109inter10));
  nor2  gate964(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate965(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate966(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate1779(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1780(.a(gate110inter0), .b(s_176), .O(gate110inter1));
  and2  gate1781(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1782(.a(s_176), .O(gate110inter3));
  inv1  gate1783(.a(s_177), .O(gate110inter4));
  nand2 gate1784(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1785(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1786(.a(G372), .O(gate110inter7));
  inv1  gate1787(.a(G373), .O(gate110inter8));
  nand2 gate1788(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1789(.a(s_177), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1790(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1791(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1792(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate575(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate576(.a(gate112inter0), .b(s_4), .O(gate112inter1));
  and2  gate577(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate578(.a(s_4), .O(gate112inter3));
  inv1  gate579(.a(s_5), .O(gate112inter4));
  nand2 gate580(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate581(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate582(.a(G376), .O(gate112inter7));
  inv1  gate583(.a(G377), .O(gate112inter8));
  nand2 gate584(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate585(.a(s_5), .b(gate112inter3), .O(gate112inter10));
  nor2  gate586(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate587(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate588(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate3123(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate3124(.a(gate115inter0), .b(s_368), .O(gate115inter1));
  and2  gate3125(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate3126(.a(s_368), .O(gate115inter3));
  inv1  gate3127(.a(s_369), .O(gate115inter4));
  nand2 gate3128(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate3129(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate3130(.a(G382), .O(gate115inter7));
  inv1  gate3131(.a(G383), .O(gate115inter8));
  nand2 gate3132(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate3133(.a(s_369), .b(gate115inter3), .O(gate115inter10));
  nor2  gate3134(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate3135(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate3136(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate869(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate870(.a(gate117inter0), .b(s_46), .O(gate117inter1));
  and2  gate871(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate872(.a(s_46), .O(gate117inter3));
  inv1  gate873(.a(s_47), .O(gate117inter4));
  nand2 gate874(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate875(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate876(.a(G386), .O(gate117inter7));
  inv1  gate877(.a(G387), .O(gate117inter8));
  nand2 gate878(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate879(.a(s_47), .b(gate117inter3), .O(gate117inter10));
  nor2  gate880(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate881(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate882(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate2087(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2088(.a(gate118inter0), .b(s_220), .O(gate118inter1));
  and2  gate2089(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2090(.a(s_220), .O(gate118inter3));
  inv1  gate2091(.a(s_221), .O(gate118inter4));
  nand2 gate2092(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2093(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2094(.a(G388), .O(gate118inter7));
  inv1  gate2095(.a(G389), .O(gate118inter8));
  nand2 gate2096(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2097(.a(s_221), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2098(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2099(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2100(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate911(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate912(.a(gate119inter0), .b(s_52), .O(gate119inter1));
  and2  gate913(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate914(.a(s_52), .O(gate119inter3));
  inv1  gate915(.a(s_53), .O(gate119inter4));
  nand2 gate916(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate917(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate918(.a(G390), .O(gate119inter7));
  inv1  gate919(.a(G391), .O(gate119inter8));
  nand2 gate920(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate921(.a(s_53), .b(gate119inter3), .O(gate119inter10));
  nor2  gate922(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate923(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate924(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate603(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate604(.a(gate121inter0), .b(s_8), .O(gate121inter1));
  and2  gate605(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate606(.a(s_8), .O(gate121inter3));
  inv1  gate607(.a(s_9), .O(gate121inter4));
  nand2 gate608(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate609(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate610(.a(G394), .O(gate121inter7));
  inv1  gate611(.a(G395), .O(gate121inter8));
  nand2 gate612(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate613(.a(s_9), .b(gate121inter3), .O(gate121inter10));
  nor2  gate614(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate615(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate616(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate2073(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2074(.a(gate122inter0), .b(s_218), .O(gate122inter1));
  and2  gate2075(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2076(.a(s_218), .O(gate122inter3));
  inv1  gate2077(.a(s_219), .O(gate122inter4));
  nand2 gate2078(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2079(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2080(.a(G396), .O(gate122inter7));
  inv1  gate2081(.a(G397), .O(gate122inter8));
  nand2 gate2082(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2083(.a(s_219), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2084(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2085(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2086(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1205(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1206(.a(gate126inter0), .b(s_94), .O(gate126inter1));
  and2  gate1207(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1208(.a(s_94), .O(gate126inter3));
  inv1  gate1209(.a(s_95), .O(gate126inter4));
  nand2 gate1210(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1211(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1212(.a(G404), .O(gate126inter7));
  inv1  gate1213(.a(G405), .O(gate126inter8));
  nand2 gate1214(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1215(.a(s_95), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1216(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1217(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1218(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate2577(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2578(.a(gate127inter0), .b(s_290), .O(gate127inter1));
  and2  gate2579(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2580(.a(s_290), .O(gate127inter3));
  inv1  gate2581(.a(s_291), .O(gate127inter4));
  nand2 gate2582(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2583(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2584(.a(G406), .O(gate127inter7));
  inv1  gate2585(.a(G407), .O(gate127inter8));
  nand2 gate2586(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2587(.a(s_291), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2588(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2589(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2590(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate2017(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2018(.a(gate128inter0), .b(s_210), .O(gate128inter1));
  and2  gate2019(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2020(.a(s_210), .O(gate128inter3));
  inv1  gate2021(.a(s_211), .O(gate128inter4));
  nand2 gate2022(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2023(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2024(.a(G408), .O(gate128inter7));
  inv1  gate2025(.a(G409), .O(gate128inter8));
  nand2 gate2026(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2027(.a(s_211), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2028(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2029(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2030(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1947(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1948(.a(gate130inter0), .b(s_200), .O(gate130inter1));
  and2  gate1949(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1950(.a(s_200), .O(gate130inter3));
  inv1  gate1951(.a(s_201), .O(gate130inter4));
  nand2 gate1952(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1953(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1954(.a(G412), .O(gate130inter7));
  inv1  gate1955(.a(G413), .O(gate130inter8));
  nand2 gate1956(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1957(.a(s_201), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1958(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1959(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1960(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2199(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2200(.a(gate132inter0), .b(s_236), .O(gate132inter1));
  and2  gate2201(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2202(.a(s_236), .O(gate132inter3));
  inv1  gate2203(.a(s_237), .O(gate132inter4));
  nand2 gate2204(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2205(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2206(.a(G416), .O(gate132inter7));
  inv1  gate2207(.a(G417), .O(gate132inter8));
  nand2 gate2208(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2209(.a(s_237), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2210(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2211(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2212(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2647(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2648(.a(gate135inter0), .b(s_300), .O(gate135inter1));
  and2  gate2649(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2650(.a(s_300), .O(gate135inter3));
  inv1  gate2651(.a(s_301), .O(gate135inter4));
  nand2 gate2652(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2653(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2654(.a(G422), .O(gate135inter7));
  inv1  gate2655(.a(G423), .O(gate135inter8));
  nand2 gate2656(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2657(.a(s_301), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2658(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2659(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2660(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1009(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1010(.a(gate139inter0), .b(s_66), .O(gate139inter1));
  and2  gate1011(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1012(.a(s_66), .O(gate139inter3));
  inv1  gate1013(.a(s_67), .O(gate139inter4));
  nand2 gate1014(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1015(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1016(.a(G438), .O(gate139inter7));
  inv1  gate1017(.a(G441), .O(gate139inter8));
  nand2 gate1018(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1019(.a(s_67), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1020(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1021(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1022(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1275(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1276(.a(gate141inter0), .b(s_104), .O(gate141inter1));
  and2  gate1277(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1278(.a(s_104), .O(gate141inter3));
  inv1  gate1279(.a(s_105), .O(gate141inter4));
  nand2 gate1280(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1281(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1282(.a(G450), .O(gate141inter7));
  inv1  gate1283(.a(G453), .O(gate141inter8));
  nand2 gate1284(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1285(.a(s_105), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1286(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1287(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1288(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate2871(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2872(.a(gate142inter0), .b(s_332), .O(gate142inter1));
  and2  gate2873(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2874(.a(s_332), .O(gate142inter3));
  inv1  gate2875(.a(s_333), .O(gate142inter4));
  nand2 gate2876(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2877(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2878(.a(G456), .O(gate142inter7));
  inv1  gate2879(.a(G459), .O(gate142inter8));
  nand2 gate2880(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2881(.a(s_333), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2882(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2883(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2884(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate2059(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2060(.a(gate143inter0), .b(s_216), .O(gate143inter1));
  and2  gate2061(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2062(.a(s_216), .O(gate143inter3));
  inv1  gate2063(.a(s_217), .O(gate143inter4));
  nand2 gate2064(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2065(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2066(.a(G462), .O(gate143inter7));
  inv1  gate2067(.a(G465), .O(gate143inter8));
  nand2 gate2068(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2069(.a(s_217), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2070(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2071(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2072(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate2353(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2354(.a(gate144inter0), .b(s_258), .O(gate144inter1));
  and2  gate2355(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2356(.a(s_258), .O(gate144inter3));
  inv1  gate2357(.a(s_259), .O(gate144inter4));
  nand2 gate2358(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2359(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2360(.a(G468), .O(gate144inter7));
  inv1  gate2361(.a(G471), .O(gate144inter8));
  nand2 gate2362(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2363(.a(s_259), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2364(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2365(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2366(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2661(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2662(.a(gate146inter0), .b(s_302), .O(gate146inter1));
  and2  gate2663(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2664(.a(s_302), .O(gate146inter3));
  inv1  gate2665(.a(s_303), .O(gate146inter4));
  nand2 gate2666(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2667(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2668(.a(G480), .O(gate146inter7));
  inv1  gate2669(.a(G483), .O(gate146inter8));
  nand2 gate2670(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2671(.a(s_303), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2672(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2673(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2674(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2773(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2774(.a(gate150inter0), .b(s_318), .O(gate150inter1));
  and2  gate2775(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2776(.a(s_318), .O(gate150inter3));
  inv1  gate2777(.a(s_319), .O(gate150inter4));
  nand2 gate2778(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2779(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2780(.a(G504), .O(gate150inter7));
  inv1  gate2781(.a(G507), .O(gate150inter8));
  nand2 gate2782(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2783(.a(s_319), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2784(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2785(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2786(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1331(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1332(.a(gate151inter0), .b(s_112), .O(gate151inter1));
  and2  gate1333(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1334(.a(s_112), .O(gate151inter3));
  inv1  gate1335(.a(s_113), .O(gate151inter4));
  nand2 gate1336(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1337(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1338(.a(G510), .O(gate151inter7));
  inv1  gate1339(.a(G513), .O(gate151inter8));
  nand2 gate1340(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1341(.a(s_113), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1342(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1343(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1344(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate617(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate618(.a(gate152inter0), .b(s_10), .O(gate152inter1));
  and2  gate619(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate620(.a(s_10), .O(gate152inter3));
  inv1  gate621(.a(s_11), .O(gate152inter4));
  nand2 gate622(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate623(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate624(.a(G516), .O(gate152inter7));
  inv1  gate625(.a(G519), .O(gate152inter8));
  nand2 gate626(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate627(.a(s_11), .b(gate152inter3), .O(gate152inter10));
  nor2  gate628(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate629(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate630(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate2395(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2396(.a(gate154inter0), .b(s_264), .O(gate154inter1));
  and2  gate2397(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2398(.a(s_264), .O(gate154inter3));
  inv1  gate2399(.a(s_265), .O(gate154inter4));
  nand2 gate2400(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2401(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2402(.a(G429), .O(gate154inter7));
  inv1  gate2403(.a(G522), .O(gate154inter8));
  nand2 gate2404(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2405(.a(s_265), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2406(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2407(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2408(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1401(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1402(.a(gate157inter0), .b(s_122), .O(gate157inter1));
  and2  gate1403(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1404(.a(s_122), .O(gate157inter3));
  inv1  gate1405(.a(s_123), .O(gate157inter4));
  nand2 gate1406(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1407(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1408(.a(G438), .O(gate157inter7));
  inv1  gate1409(.a(G528), .O(gate157inter8));
  nand2 gate1410(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1411(.a(s_123), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1412(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1413(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1414(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1737(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1738(.a(gate160inter0), .b(s_170), .O(gate160inter1));
  and2  gate1739(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1740(.a(s_170), .O(gate160inter3));
  inv1  gate1741(.a(s_171), .O(gate160inter4));
  nand2 gate1742(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1743(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1744(.a(G447), .O(gate160inter7));
  inv1  gate1745(.a(G531), .O(gate160inter8));
  nand2 gate1746(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1747(.a(s_171), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1748(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1749(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1750(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate813(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate814(.a(gate161inter0), .b(s_38), .O(gate161inter1));
  and2  gate815(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate816(.a(s_38), .O(gate161inter3));
  inv1  gate817(.a(s_39), .O(gate161inter4));
  nand2 gate818(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate819(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate820(.a(G450), .O(gate161inter7));
  inv1  gate821(.a(G534), .O(gate161inter8));
  nand2 gate822(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate823(.a(s_39), .b(gate161inter3), .O(gate161inter10));
  nor2  gate824(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate825(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate826(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate701(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate702(.a(gate166inter0), .b(s_22), .O(gate166inter1));
  and2  gate703(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate704(.a(s_22), .O(gate166inter3));
  inv1  gate705(.a(s_23), .O(gate166inter4));
  nand2 gate706(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate707(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate708(.a(G465), .O(gate166inter7));
  inv1  gate709(.a(G540), .O(gate166inter8));
  nand2 gate710(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate711(.a(s_23), .b(gate166inter3), .O(gate166inter10));
  nor2  gate712(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate713(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate714(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1919(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1920(.a(gate171inter0), .b(s_196), .O(gate171inter1));
  and2  gate1921(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1922(.a(s_196), .O(gate171inter3));
  inv1  gate1923(.a(s_197), .O(gate171inter4));
  nand2 gate1924(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1925(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1926(.a(G480), .O(gate171inter7));
  inv1  gate1927(.a(G549), .O(gate171inter8));
  nand2 gate1928(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1929(.a(s_197), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1930(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1931(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1932(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1569(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1570(.a(gate181inter0), .b(s_146), .O(gate181inter1));
  and2  gate1571(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1572(.a(s_146), .O(gate181inter3));
  inv1  gate1573(.a(s_147), .O(gate181inter4));
  nand2 gate1574(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1575(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1576(.a(G510), .O(gate181inter7));
  inv1  gate1577(.a(G564), .O(gate181inter8));
  nand2 gate1578(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1579(.a(s_147), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1580(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1581(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1582(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1443(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1444(.a(gate183inter0), .b(s_128), .O(gate183inter1));
  and2  gate1445(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1446(.a(s_128), .O(gate183inter3));
  inv1  gate1447(.a(s_129), .O(gate183inter4));
  nand2 gate1448(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1449(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1450(.a(G516), .O(gate183inter7));
  inv1  gate1451(.a(G567), .O(gate183inter8));
  nand2 gate1452(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1453(.a(s_129), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1454(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1455(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1456(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1835(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1836(.a(gate185inter0), .b(s_184), .O(gate185inter1));
  and2  gate1837(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1838(.a(s_184), .O(gate185inter3));
  inv1  gate1839(.a(s_185), .O(gate185inter4));
  nand2 gate1840(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1841(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1842(.a(G570), .O(gate185inter7));
  inv1  gate1843(.a(G571), .O(gate185inter8));
  nand2 gate1844(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1845(.a(s_185), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1846(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1847(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1848(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1163(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1164(.a(gate189inter0), .b(s_88), .O(gate189inter1));
  and2  gate1165(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1166(.a(s_88), .O(gate189inter3));
  inv1  gate1167(.a(s_89), .O(gate189inter4));
  nand2 gate1168(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1169(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1170(.a(G578), .O(gate189inter7));
  inv1  gate1171(.a(G579), .O(gate189inter8));
  nand2 gate1172(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1173(.a(s_89), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1174(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1175(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1176(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate631(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate632(.a(gate191inter0), .b(s_12), .O(gate191inter1));
  and2  gate633(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate634(.a(s_12), .O(gate191inter3));
  inv1  gate635(.a(s_13), .O(gate191inter4));
  nand2 gate636(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate637(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate638(.a(G582), .O(gate191inter7));
  inv1  gate639(.a(G583), .O(gate191inter8));
  nand2 gate640(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate641(.a(s_13), .b(gate191inter3), .O(gate191inter10));
  nor2  gate642(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate643(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate644(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate799(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate800(.a(gate192inter0), .b(s_36), .O(gate192inter1));
  and2  gate801(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate802(.a(s_36), .O(gate192inter3));
  inv1  gate803(.a(s_37), .O(gate192inter4));
  nand2 gate804(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate805(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate806(.a(G584), .O(gate192inter7));
  inv1  gate807(.a(G585), .O(gate192inter8));
  nand2 gate808(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate809(.a(s_37), .b(gate192inter3), .O(gate192inter10));
  nor2  gate810(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate811(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate812(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2423(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2424(.a(gate193inter0), .b(s_268), .O(gate193inter1));
  and2  gate2425(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2426(.a(s_268), .O(gate193inter3));
  inv1  gate2427(.a(s_269), .O(gate193inter4));
  nand2 gate2428(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2429(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2430(.a(G586), .O(gate193inter7));
  inv1  gate2431(.a(G587), .O(gate193inter8));
  nand2 gate2432(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2433(.a(s_269), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2434(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2435(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2436(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2535(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2536(.a(gate200inter0), .b(s_284), .O(gate200inter1));
  and2  gate2537(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2538(.a(s_284), .O(gate200inter3));
  inv1  gate2539(.a(s_285), .O(gate200inter4));
  nand2 gate2540(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2541(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2542(.a(G600), .O(gate200inter7));
  inv1  gate2543(.a(G601), .O(gate200inter8));
  nand2 gate2544(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2545(.a(s_285), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2546(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2547(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2548(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2913(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2914(.a(gate204inter0), .b(s_338), .O(gate204inter1));
  and2  gate2915(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2916(.a(s_338), .O(gate204inter3));
  inv1  gate2917(.a(s_339), .O(gate204inter4));
  nand2 gate2918(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2919(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2920(.a(G607), .O(gate204inter7));
  inv1  gate2921(.a(G617), .O(gate204inter8));
  nand2 gate2922(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2923(.a(s_339), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2924(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2925(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2926(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate757(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate758(.a(gate205inter0), .b(s_30), .O(gate205inter1));
  and2  gate759(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate760(.a(s_30), .O(gate205inter3));
  inv1  gate761(.a(s_31), .O(gate205inter4));
  nand2 gate762(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate763(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate764(.a(G622), .O(gate205inter7));
  inv1  gate765(.a(G627), .O(gate205inter8));
  nand2 gate766(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate767(.a(s_31), .b(gate205inter3), .O(gate205inter10));
  nor2  gate768(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate769(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate770(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2129(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2130(.a(gate207inter0), .b(s_226), .O(gate207inter1));
  and2  gate2131(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2132(.a(s_226), .O(gate207inter3));
  inv1  gate2133(.a(s_227), .O(gate207inter4));
  nand2 gate2134(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2135(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2136(.a(G622), .O(gate207inter7));
  inv1  gate2137(.a(G632), .O(gate207inter8));
  nand2 gate2138(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2139(.a(s_227), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2140(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2141(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2142(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate2045(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2046(.a(gate208inter0), .b(s_214), .O(gate208inter1));
  and2  gate2047(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2048(.a(s_214), .O(gate208inter3));
  inv1  gate2049(.a(s_215), .O(gate208inter4));
  nand2 gate2050(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2051(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2052(.a(G627), .O(gate208inter7));
  inv1  gate2053(.a(G637), .O(gate208inter8));
  nand2 gate2054(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2055(.a(s_215), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2056(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2057(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2058(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2703(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2704(.a(gate210inter0), .b(s_308), .O(gate210inter1));
  and2  gate2705(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2706(.a(s_308), .O(gate210inter3));
  inv1  gate2707(.a(s_309), .O(gate210inter4));
  nand2 gate2708(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2709(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2710(.a(G607), .O(gate210inter7));
  inv1  gate2711(.a(G666), .O(gate210inter8));
  nand2 gate2712(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2713(.a(s_309), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2714(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2715(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2716(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate3095(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate3096(.a(gate213inter0), .b(s_364), .O(gate213inter1));
  and2  gate3097(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate3098(.a(s_364), .O(gate213inter3));
  inv1  gate3099(.a(s_365), .O(gate213inter4));
  nand2 gate3100(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate3101(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate3102(.a(G602), .O(gate213inter7));
  inv1  gate3103(.a(G672), .O(gate213inter8));
  nand2 gate3104(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate3105(.a(s_365), .b(gate213inter3), .O(gate213inter10));
  nor2  gate3106(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate3107(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate3108(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1667(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1668(.a(gate214inter0), .b(s_160), .O(gate214inter1));
  and2  gate1669(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1670(.a(s_160), .O(gate214inter3));
  inv1  gate1671(.a(s_161), .O(gate214inter4));
  nand2 gate1672(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1673(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1674(.a(G612), .O(gate214inter7));
  inv1  gate1675(.a(G672), .O(gate214inter8));
  nand2 gate1676(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1677(.a(s_161), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1678(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1679(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1680(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2227(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2228(.a(gate215inter0), .b(s_240), .O(gate215inter1));
  and2  gate2229(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2230(.a(s_240), .O(gate215inter3));
  inv1  gate2231(.a(s_241), .O(gate215inter4));
  nand2 gate2232(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2233(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2234(.a(G607), .O(gate215inter7));
  inv1  gate2235(.a(G675), .O(gate215inter8));
  nand2 gate2236(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2237(.a(s_241), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2238(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2239(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2240(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1191(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1192(.a(gate216inter0), .b(s_92), .O(gate216inter1));
  and2  gate1193(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1194(.a(s_92), .O(gate216inter3));
  inv1  gate1195(.a(s_93), .O(gate216inter4));
  nand2 gate1196(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1197(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1198(.a(G617), .O(gate216inter7));
  inv1  gate1199(.a(G675), .O(gate216inter8));
  nand2 gate1200(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1201(.a(s_93), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1202(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1203(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1204(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate2899(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2900(.a(gate217inter0), .b(s_336), .O(gate217inter1));
  and2  gate2901(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2902(.a(s_336), .O(gate217inter3));
  inv1  gate2903(.a(s_337), .O(gate217inter4));
  nand2 gate2904(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2905(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2906(.a(G622), .O(gate217inter7));
  inv1  gate2907(.a(G678), .O(gate217inter8));
  nand2 gate2908(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2909(.a(s_337), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2910(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2911(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2912(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2367(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2368(.a(gate220inter0), .b(s_260), .O(gate220inter1));
  and2  gate2369(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2370(.a(s_260), .O(gate220inter3));
  inv1  gate2371(.a(s_261), .O(gate220inter4));
  nand2 gate2372(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2373(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2374(.a(G637), .O(gate220inter7));
  inv1  gate2375(.a(G681), .O(gate220inter8));
  nand2 gate2376(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2377(.a(s_261), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2378(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2379(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2380(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate897(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate898(.a(gate221inter0), .b(s_50), .O(gate221inter1));
  and2  gate899(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate900(.a(s_50), .O(gate221inter3));
  inv1  gate901(.a(s_51), .O(gate221inter4));
  nand2 gate902(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate903(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate904(.a(G622), .O(gate221inter7));
  inv1  gate905(.a(G684), .O(gate221inter8));
  nand2 gate906(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate907(.a(s_51), .b(gate221inter3), .O(gate221inter10));
  nor2  gate908(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate909(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate910(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1373(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1374(.a(gate222inter0), .b(s_118), .O(gate222inter1));
  and2  gate1375(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1376(.a(s_118), .O(gate222inter3));
  inv1  gate1377(.a(s_119), .O(gate222inter4));
  nand2 gate1378(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1379(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1380(.a(G632), .O(gate222inter7));
  inv1  gate1381(.a(G684), .O(gate222inter8));
  nand2 gate1382(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1383(.a(s_119), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1384(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1385(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1386(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2815(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2816(.a(gate223inter0), .b(s_324), .O(gate223inter1));
  and2  gate2817(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2818(.a(s_324), .O(gate223inter3));
  inv1  gate2819(.a(s_325), .O(gate223inter4));
  nand2 gate2820(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2821(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2822(.a(G627), .O(gate223inter7));
  inv1  gate2823(.a(G687), .O(gate223inter8));
  nand2 gate2824(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2825(.a(s_325), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2826(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2827(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2828(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2605(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2606(.a(gate229inter0), .b(s_294), .O(gate229inter1));
  and2  gate2607(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2608(.a(s_294), .O(gate229inter3));
  inv1  gate2609(.a(s_295), .O(gate229inter4));
  nand2 gate2610(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2611(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2612(.a(G698), .O(gate229inter7));
  inv1  gate2613(.a(G699), .O(gate229inter8));
  nand2 gate2614(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2615(.a(s_295), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2616(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2617(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2618(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1429(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1430(.a(gate230inter0), .b(s_126), .O(gate230inter1));
  and2  gate1431(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1432(.a(s_126), .O(gate230inter3));
  inv1  gate1433(.a(s_127), .O(gate230inter4));
  nand2 gate1434(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1435(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1436(.a(G700), .O(gate230inter7));
  inv1  gate1437(.a(G701), .O(gate230inter8));
  nand2 gate1438(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1439(.a(s_127), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1440(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1441(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1442(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate3025(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate3026(.a(gate232inter0), .b(s_354), .O(gate232inter1));
  and2  gate3027(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate3028(.a(s_354), .O(gate232inter3));
  inv1  gate3029(.a(s_355), .O(gate232inter4));
  nand2 gate3030(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate3031(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate3032(.a(G704), .O(gate232inter7));
  inv1  gate3033(.a(G705), .O(gate232inter8));
  nand2 gate3034(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate3035(.a(s_355), .b(gate232inter3), .O(gate232inter10));
  nor2  gate3036(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate3037(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate3038(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1121(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1122(.a(gate233inter0), .b(s_82), .O(gate233inter1));
  and2  gate1123(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1124(.a(s_82), .O(gate233inter3));
  inv1  gate1125(.a(s_83), .O(gate233inter4));
  nand2 gate1126(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1127(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1128(.a(G242), .O(gate233inter7));
  inv1  gate1129(.a(G718), .O(gate233inter8));
  nand2 gate1130(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1131(.a(s_83), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1132(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1133(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1134(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2997(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2998(.a(gate236inter0), .b(s_350), .O(gate236inter1));
  and2  gate2999(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate3000(.a(s_350), .O(gate236inter3));
  inv1  gate3001(.a(s_351), .O(gate236inter4));
  nand2 gate3002(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate3003(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate3004(.a(G251), .O(gate236inter7));
  inv1  gate3005(.a(G727), .O(gate236inter8));
  nand2 gate3006(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate3007(.a(s_351), .b(gate236inter3), .O(gate236inter10));
  nor2  gate3008(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate3009(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate3010(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1457(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1458(.a(gate241inter0), .b(s_130), .O(gate241inter1));
  and2  gate1459(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1460(.a(s_130), .O(gate241inter3));
  inv1  gate1461(.a(s_131), .O(gate241inter4));
  nand2 gate1462(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1463(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1464(.a(G242), .O(gate241inter7));
  inv1  gate1465(.a(G730), .O(gate241inter8));
  nand2 gate1466(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1467(.a(s_131), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1468(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1469(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1470(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate883(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate884(.a(gate243inter0), .b(s_48), .O(gate243inter1));
  and2  gate885(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate886(.a(s_48), .O(gate243inter3));
  inv1  gate887(.a(s_49), .O(gate243inter4));
  nand2 gate888(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate889(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate890(.a(G245), .O(gate243inter7));
  inv1  gate891(.a(G733), .O(gate243inter8));
  nand2 gate892(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate893(.a(s_49), .b(gate243inter3), .O(gate243inter10));
  nor2  gate894(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate895(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate896(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2745(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2746(.a(gate245inter0), .b(s_314), .O(gate245inter1));
  and2  gate2747(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2748(.a(s_314), .O(gate245inter3));
  inv1  gate2749(.a(s_315), .O(gate245inter4));
  nand2 gate2750(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2751(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2752(.a(G248), .O(gate245inter7));
  inv1  gate2753(.a(G736), .O(gate245inter8));
  nand2 gate2754(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2755(.a(s_315), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2756(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2757(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2758(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1387(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1388(.a(gate246inter0), .b(s_120), .O(gate246inter1));
  and2  gate1389(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1390(.a(s_120), .O(gate246inter3));
  inv1  gate1391(.a(s_121), .O(gate246inter4));
  nand2 gate1392(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1393(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1394(.a(G724), .O(gate246inter7));
  inv1  gate1395(.a(G736), .O(gate246inter8));
  nand2 gate1396(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1397(.a(s_121), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1398(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1399(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1400(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1709(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1710(.a(gate247inter0), .b(s_166), .O(gate247inter1));
  and2  gate1711(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1712(.a(s_166), .O(gate247inter3));
  inv1  gate1713(.a(s_167), .O(gate247inter4));
  nand2 gate1714(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1715(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1716(.a(G251), .O(gate247inter7));
  inv1  gate1717(.a(G739), .O(gate247inter8));
  nand2 gate1718(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1719(.a(s_167), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1720(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1721(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1722(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2591(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2592(.a(gate248inter0), .b(s_292), .O(gate248inter1));
  and2  gate2593(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2594(.a(s_292), .O(gate248inter3));
  inv1  gate2595(.a(s_293), .O(gate248inter4));
  nand2 gate2596(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2597(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2598(.a(G727), .O(gate248inter7));
  inv1  gate2599(.a(G739), .O(gate248inter8));
  nand2 gate2600(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2601(.a(s_293), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2602(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2603(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2604(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2465(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2466(.a(gate252inter0), .b(s_274), .O(gate252inter1));
  and2  gate2467(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2468(.a(s_274), .O(gate252inter3));
  inv1  gate2469(.a(s_275), .O(gate252inter4));
  nand2 gate2470(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2471(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2472(.a(G709), .O(gate252inter7));
  inv1  gate2473(.a(G745), .O(gate252inter8));
  nand2 gate2474(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2475(.a(s_275), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2476(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2477(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2478(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate659(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate660(.a(gate253inter0), .b(s_16), .O(gate253inter1));
  and2  gate661(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate662(.a(s_16), .O(gate253inter3));
  inv1  gate663(.a(s_17), .O(gate253inter4));
  nand2 gate664(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate665(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate666(.a(G260), .O(gate253inter7));
  inv1  gate667(.a(G748), .O(gate253inter8));
  nand2 gate668(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate669(.a(s_17), .b(gate253inter3), .O(gate253inter10));
  nor2  gate670(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate671(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate672(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2941(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2942(.a(gate257inter0), .b(s_342), .O(gate257inter1));
  and2  gate2943(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2944(.a(s_342), .O(gate257inter3));
  inv1  gate2945(.a(s_343), .O(gate257inter4));
  nand2 gate2946(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2947(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2948(.a(G754), .O(gate257inter7));
  inv1  gate2949(.a(G755), .O(gate257inter8));
  nand2 gate2950(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2951(.a(s_343), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2952(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2953(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2954(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1471(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1472(.a(gate258inter0), .b(s_132), .O(gate258inter1));
  and2  gate1473(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1474(.a(s_132), .O(gate258inter3));
  inv1  gate1475(.a(s_133), .O(gate258inter4));
  nand2 gate1476(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1477(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1478(.a(G756), .O(gate258inter7));
  inv1  gate1479(.a(G757), .O(gate258inter8));
  nand2 gate1480(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1481(.a(s_133), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1482(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1483(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1484(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate3067(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate3068(.a(gate259inter0), .b(s_360), .O(gate259inter1));
  and2  gate3069(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate3070(.a(s_360), .O(gate259inter3));
  inv1  gate3071(.a(s_361), .O(gate259inter4));
  nand2 gate3072(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate3073(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate3074(.a(G758), .O(gate259inter7));
  inv1  gate3075(.a(G759), .O(gate259inter8));
  nand2 gate3076(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate3077(.a(s_361), .b(gate259inter3), .O(gate259inter10));
  nor2  gate3078(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate3079(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate3080(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate2437(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2438(.a(gate260inter0), .b(s_270), .O(gate260inter1));
  and2  gate2439(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2440(.a(s_270), .O(gate260inter3));
  inv1  gate2441(.a(s_271), .O(gate260inter4));
  nand2 gate2442(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2443(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2444(.a(G760), .O(gate260inter7));
  inv1  gate2445(.a(G761), .O(gate260inter8));
  nand2 gate2446(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2447(.a(s_271), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2448(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2449(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2450(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1233(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1234(.a(gate262inter0), .b(s_98), .O(gate262inter1));
  and2  gate1235(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1236(.a(s_98), .O(gate262inter3));
  inv1  gate1237(.a(s_99), .O(gate262inter4));
  nand2 gate1238(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1239(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1240(.a(G764), .O(gate262inter7));
  inv1  gate1241(.a(G765), .O(gate262inter8));
  nand2 gate1242(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1243(.a(s_99), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1244(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1245(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1246(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate2283(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2284(.a(gate263inter0), .b(s_248), .O(gate263inter1));
  and2  gate2285(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2286(.a(s_248), .O(gate263inter3));
  inv1  gate2287(.a(s_249), .O(gate263inter4));
  nand2 gate2288(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2289(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2290(.a(G766), .O(gate263inter7));
  inv1  gate2291(.a(G767), .O(gate263inter8));
  nand2 gate2292(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2293(.a(s_249), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2294(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2295(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2296(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2241(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2242(.a(gate265inter0), .b(s_242), .O(gate265inter1));
  and2  gate2243(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2244(.a(s_242), .O(gate265inter3));
  inv1  gate2245(.a(s_243), .O(gate265inter4));
  nand2 gate2246(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2247(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2248(.a(G642), .O(gate265inter7));
  inv1  gate2249(.a(G770), .O(gate265inter8));
  nand2 gate2250(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2251(.a(s_243), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2252(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2253(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2254(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate3011(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate3012(.a(gate267inter0), .b(s_352), .O(gate267inter1));
  and2  gate3013(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate3014(.a(s_352), .O(gate267inter3));
  inv1  gate3015(.a(s_353), .O(gate267inter4));
  nand2 gate3016(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate3017(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate3018(.a(G648), .O(gate267inter7));
  inv1  gate3019(.a(G776), .O(gate267inter8));
  nand2 gate3020(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate3021(.a(s_353), .b(gate267inter3), .O(gate267inter10));
  nor2  gate3022(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate3023(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate3024(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1597(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1598(.a(gate269inter0), .b(s_150), .O(gate269inter1));
  and2  gate1599(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1600(.a(s_150), .O(gate269inter3));
  inv1  gate1601(.a(s_151), .O(gate269inter4));
  nand2 gate1602(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1603(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1604(.a(G654), .O(gate269inter7));
  inv1  gate1605(.a(G782), .O(gate269inter8));
  nand2 gate1606(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1607(.a(s_151), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1608(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1609(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1610(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1261(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1262(.a(gate275inter0), .b(s_102), .O(gate275inter1));
  and2  gate1263(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1264(.a(s_102), .O(gate275inter3));
  inv1  gate1265(.a(s_103), .O(gate275inter4));
  nand2 gate1266(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1267(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1268(.a(G645), .O(gate275inter7));
  inv1  gate1269(.a(G797), .O(gate275inter8));
  nand2 gate1270(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1271(.a(s_103), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1272(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1273(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1274(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1177(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1178(.a(gate276inter0), .b(s_90), .O(gate276inter1));
  and2  gate1179(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1180(.a(s_90), .O(gate276inter3));
  inv1  gate1181(.a(s_91), .O(gate276inter4));
  nand2 gate1182(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1183(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1184(.a(G773), .O(gate276inter7));
  inv1  gate1185(.a(G797), .O(gate276inter8));
  nand2 gate1186(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1187(.a(s_91), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1188(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1189(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1190(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1905(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1906(.a(gate279inter0), .b(s_194), .O(gate279inter1));
  and2  gate1907(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1908(.a(s_194), .O(gate279inter3));
  inv1  gate1909(.a(s_195), .O(gate279inter4));
  nand2 gate1910(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1911(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1912(.a(G651), .O(gate279inter7));
  inv1  gate1913(.a(G803), .O(gate279inter8));
  nand2 gate1914(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1915(.a(s_195), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1916(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1917(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1918(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2759(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2760(.a(gate282inter0), .b(s_316), .O(gate282inter1));
  and2  gate2761(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2762(.a(s_316), .O(gate282inter3));
  inv1  gate2763(.a(s_317), .O(gate282inter4));
  nand2 gate2764(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2765(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2766(.a(G782), .O(gate282inter7));
  inv1  gate2767(.a(G806), .O(gate282inter8));
  nand2 gate2768(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2769(.a(s_317), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2770(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2771(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2772(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1037(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1038(.a(gate283inter0), .b(s_70), .O(gate283inter1));
  and2  gate1039(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1040(.a(s_70), .O(gate283inter3));
  inv1  gate1041(.a(s_71), .O(gate283inter4));
  nand2 gate1042(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1043(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1044(.a(G657), .O(gate283inter7));
  inv1  gate1045(.a(G809), .O(gate283inter8));
  nand2 gate1046(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1047(.a(s_71), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1048(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1049(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1050(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1765(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1766(.a(gate288inter0), .b(s_174), .O(gate288inter1));
  and2  gate1767(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1768(.a(s_174), .O(gate288inter3));
  inv1  gate1769(.a(s_175), .O(gate288inter4));
  nand2 gate1770(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1771(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1772(.a(G791), .O(gate288inter7));
  inv1  gate1773(.a(G815), .O(gate288inter8));
  nand2 gate1774(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1775(.a(s_175), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1776(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1777(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1778(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate925(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate926(.a(gate290inter0), .b(s_54), .O(gate290inter1));
  and2  gate927(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate928(.a(s_54), .O(gate290inter3));
  inv1  gate929(.a(s_55), .O(gate290inter4));
  nand2 gate930(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate931(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate932(.a(G820), .O(gate290inter7));
  inv1  gate933(.a(G821), .O(gate290inter8));
  nand2 gate934(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate935(.a(s_55), .b(gate290inter3), .O(gate290inter10));
  nor2  gate936(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate937(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate938(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate1513(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1514(.a(gate291inter0), .b(s_138), .O(gate291inter1));
  and2  gate1515(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1516(.a(s_138), .O(gate291inter3));
  inv1  gate1517(.a(s_139), .O(gate291inter4));
  nand2 gate1518(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1519(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1520(.a(G822), .O(gate291inter7));
  inv1  gate1521(.a(G823), .O(gate291inter8));
  nand2 gate1522(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1523(.a(s_139), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1524(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1525(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1526(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1051(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1052(.a(gate292inter0), .b(s_72), .O(gate292inter1));
  and2  gate1053(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1054(.a(s_72), .O(gate292inter3));
  inv1  gate1055(.a(s_73), .O(gate292inter4));
  nand2 gate1056(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1057(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1058(.a(G824), .O(gate292inter7));
  inv1  gate1059(.a(G825), .O(gate292inter8));
  nand2 gate1060(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1061(.a(s_73), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1062(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1063(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1064(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2493(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2494(.a(gate296inter0), .b(s_278), .O(gate296inter1));
  and2  gate2495(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2496(.a(s_278), .O(gate296inter3));
  inv1  gate2497(.a(s_279), .O(gate296inter4));
  nand2 gate2498(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2499(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2500(.a(G826), .O(gate296inter7));
  inv1  gate2501(.a(G827), .O(gate296inter8));
  nand2 gate2502(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2503(.a(s_279), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2504(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2505(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2506(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate547(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate548(.a(gate390inter0), .b(s_0), .O(gate390inter1));
  and2  gate549(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate550(.a(s_0), .O(gate390inter3));
  inv1  gate551(.a(s_1), .O(gate390inter4));
  nand2 gate552(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate553(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate554(.a(G4), .O(gate390inter7));
  inv1  gate555(.a(G1045), .O(gate390inter8));
  nand2 gate556(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate557(.a(s_1), .b(gate390inter3), .O(gate390inter10));
  nor2  gate558(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate559(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate560(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2031(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2032(.a(gate392inter0), .b(s_212), .O(gate392inter1));
  and2  gate2033(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2034(.a(s_212), .O(gate392inter3));
  inv1  gate2035(.a(s_213), .O(gate392inter4));
  nand2 gate2036(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2037(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2038(.a(G6), .O(gate392inter7));
  inv1  gate2039(.a(G1051), .O(gate392inter8));
  nand2 gate2040(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2041(.a(s_213), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2042(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2043(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2044(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2675(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2676(.a(gate396inter0), .b(s_304), .O(gate396inter1));
  and2  gate2677(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2678(.a(s_304), .O(gate396inter3));
  inv1  gate2679(.a(s_305), .O(gate396inter4));
  nand2 gate2680(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2681(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2682(.a(G10), .O(gate396inter7));
  inv1  gate2683(.a(G1063), .O(gate396inter8));
  nand2 gate2684(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2685(.a(s_305), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2686(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2687(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2688(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1303(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1304(.a(gate398inter0), .b(s_108), .O(gate398inter1));
  and2  gate1305(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1306(.a(s_108), .O(gate398inter3));
  inv1  gate1307(.a(s_109), .O(gate398inter4));
  nand2 gate1308(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1309(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1310(.a(G12), .O(gate398inter7));
  inv1  gate1311(.a(G1069), .O(gate398inter8));
  nand2 gate1312(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1313(.a(s_109), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1314(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1315(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1316(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate2507(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate2508(.a(gate400inter0), .b(s_280), .O(gate400inter1));
  and2  gate2509(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate2510(.a(s_280), .O(gate400inter3));
  inv1  gate2511(.a(s_281), .O(gate400inter4));
  nand2 gate2512(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate2513(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate2514(.a(G14), .O(gate400inter7));
  inv1  gate2515(.a(G1075), .O(gate400inter8));
  nand2 gate2516(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate2517(.a(s_281), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2518(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2519(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2520(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1317(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1318(.a(gate401inter0), .b(s_110), .O(gate401inter1));
  and2  gate1319(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1320(.a(s_110), .O(gate401inter3));
  inv1  gate1321(.a(s_111), .O(gate401inter4));
  nand2 gate1322(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1323(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1324(.a(G15), .O(gate401inter7));
  inv1  gate1325(.a(G1078), .O(gate401inter8));
  nand2 gate1326(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1327(.a(s_111), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1328(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1329(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1330(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2213(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2214(.a(gate403inter0), .b(s_238), .O(gate403inter1));
  and2  gate2215(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2216(.a(s_238), .O(gate403inter3));
  inv1  gate2217(.a(s_239), .O(gate403inter4));
  nand2 gate2218(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2219(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2220(.a(G17), .O(gate403inter7));
  inv1  gate2221(.a(G1084), .O(gate403inter8));
  nand2 gate2222(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2223(.a(s_239), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2224(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2225(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2226(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1653(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1654(.a(gate407inter0), .b(s_158), .O(gate407inter1));
  and2  gate1655(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1656(.a(s_158), .O(gate407inter3));
  inv1  gate1657(.a(s_159), .O(gate407inter4));
  nand2 gate1658(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1659(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1660(.a(G21), .O(gate407inter7));
  inv1  gate1661(.a(G1096), .O(gate407inter8));
  nand2 gate1662(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1663(.a(s_159), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1664(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1665(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1666(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate743(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate744(.a(gate408inter0), .b(s_28), .O(gate408inter1));
  and2  gate745(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate746(.a(s_28), .O(gate408inter3));
  inv1  gate747(.a(s_29), .O(gate408inter4));
  nand2 gate748(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate749(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate750(.a(G22), .O(gate408inter7));
  inv1  gate751(.a(G1099), .O(gate408inter8));
  nand2 gate752(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate753(.a(s_29), .b(gate408inter3), .O(gate408inter10));
  nor2  gate754(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate755(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate756(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate3081(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate3082(.a(gate411inter0), .b(s_362), .O(gate411inter1));
  and2  gate3083(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate3084(.a(s_362), .O(gate411inter3));
  inv1  gate3085(.a(s_363), .O(gate411inter4));
  nand2 gate3086(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate3087(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate3088(.a(G25), .O(gate411inter7));
  inv1  gate3089(.a(G1108), .O(gate411inter8));
  nand2 gate3090(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate3091(.a(s_363), .b(gate411inter3), .O(gate411inter10));
  nor2  gate3092(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate3093(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate3094(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2843(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2844(.a(gate412inter0), .b(s_328), .O(gate412inter1));
  and2  gate2845(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2846(.a(s_328), .O(gate412inter3));
  inv1  gate2847(.a(s_329), .O(gate412inter4));
  nand2 gate2848(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2849(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2850(.a(G26), .O(gate412inter7));
  inv1  gate2851(.a(G1111), .O(gate412inter8));
  nand2 gate2852(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2853(.a(s_329), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2854(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2855(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2856(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2311(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2312(.a(gate415inter0), .b(s_252), .O(gate415inter1));
  and2  gate2313(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2314(.a(s_252), .O(gate415inter3));
  inv1  gate2315(.a(s_253), .O(gate415inter4));
  nand2 gate2316(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2317(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2318(.a(G29), .O(gate415inter7));
  inv1  gate2319(.a(G1120), .O(gate415inter8));
  nand2 gate2320(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2321(.a(s_253), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2322(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2323(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2324(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1583(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1584(.a(gate416inter0), .b(s_148), .O(gate416inter1));
  and2  gate1585(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1586(.a(s_148), .O(gate416inter3));
  inv1  gate1587(.a(s_149), .O(gate416inter4));
  nand2 gate1588(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1589(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1590(.a(G30), .O(gate416inter7));
  inv1  gate1591(.a(G1123), .O(gate416inter8));
  nand2 gate1592(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1593(.a(s_149), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1594(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1595(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1596(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate2479(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2480(.a(gate418inter0), .b(s_276), .O(gate418inter1));
  and2  gate2481(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2482(.a(s_276), .O(gate418inter3));
  inv1  gate2483(.a(s_277), .O(gate418inter4));
  nand2 gate2484(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2485(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2486(.a(G32), .O(gate418inter7));
  inv1  gate2487(.a(G1129), .O(gate418inter8));
  nand2 gate2488(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2489(.a(s_277), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2490(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2491(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2492(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1289(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1290(.a(gate419inter0), .b(s_106), .O(gate419inter1));
  and2  gate1291(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1292(.a(s_106), .O(gate419inter3));
  inv1  gate1293(.a(s_107), .O(gate419inter4));
  nand2 gate1294(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1295(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1296(.a(G1), .O(gate419inter7));
  inv1  gate1297(.a(G1132), .O(gate419inter8));
  nand2 gate1298(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1299(.a(s_107), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1300(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1301(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1302(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1527(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1528(.a(gate420inter0), .b(s_140), .O(gate420inter1));
  and2  gate1529(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1530(.a(s_140), .O(gate420inter3));
  inv1  gate1531(.a(s_141), .O(gate420inter4));
  nand2 gate1532(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1533(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1534(.a(G1036), .O(gate420inter7));
  inv1  gate1535(.a(G1132), .O(gate420inter8));
  nand2 gate1536(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1537(.a(s_141), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1538(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1539(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1540(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1639(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1640(.a(gate421inter0), .b(s_156), .O(gate421inter1));
  and2  gate1641(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1642(.a(s_156), .O(gate421inter3));
  inv1  gate1643(.a(s_157), .O(gate421inter4));
  nand2 gate1644(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1645(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1646(.a(G2), .O(gate421inter7));
  inv1  gate1647(.a(G1135), .O(gate421inter8));
  nand2 gate1648(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1649(.a(s_157), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1650(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1651(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1652(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate995(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate996(.a(gate422inter0), .b(s_64), .O(gate422inter1));
  and2  gate997(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate998(.a(s_64), .O(gate422inter3));
  inv1  gate999(.a(s_65), .O(gate422inter4));
  nand2 gate1000(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1001(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1002(.a(G1039), .O(gate422inter7));
  inv1  gate1003(.a(G1135), .O(gate422inter8));
  nand2 gate1004(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1005(.a(s_65), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1006(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1007(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1008(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate715(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate716(.a(gate423inter0), .b(s_24), .O(gate423inter1));
  and2  gate717(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate718(.a(s_24), .O(gate423inter3));
  inv1  gate719(.a(s_25), .O(gate423inter4));
  nand2 gate720(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate721(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate722(.a(G3), .O(gate423inter7));
  inv1  gate723(.a(G1138), .O(gate423inter8));
  nand2 gate724(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate725(.a(s_25), .b(gate423inter3), .O(gate423inter10));
  nor2  gate726(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate727(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate728(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1499(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1500(.a(gate424inter0), .b(s_136), .O(gate424inter1));
  and2  gate1501(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1502(.a(s_136), .O(gate424inter3));
  inv1  gate1503(.a(s_137), .O(gate424inter4));
  nand2 gate1504(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1505(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1506(.a(G1042), .O(gate424inter7));
  inv1  gate1507(.a(G1138), .O(gate424inter8));
  nand2 gate1508(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1509(.a(s_137), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1510(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1511(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1512(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate2451(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2452(.a(gate425inter0), .b(s_272), .O(gate425inter1));
  and2  gate2453(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2454(.a(s_272), .O(gate425inter3));
  inv1  gate2455(.a(s_273), .O(gate425inter4));
  nand2 gate2456(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2457(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2458(.a(G4), .O(gate425inter7));
  inv1  gate2459(.a(G1141), .O(gate425inter8));
  nand2 gate2460(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2461(.a(s_273), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2462(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2463(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2464(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate3109(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate3110(.a(gate428inter0), .b(s_366), .O(gate428inter1));
  and2  gate3111(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate3112(.a(s_366), .O(gate428inter3));
  inv1  gate3113(.a(s_367), .O(gate428inter4));
  nand2 gate3114(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate3115(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate3116(.a(G1048), .O(gate428inter7));
  inv1  gate3117(.a(G1144), .O(gate428inter8));
  nand2 gate3118(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate3119(.a(s_367), .b(gate428inter3), .O(gate428inter10));
  nor2  gate3120(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate3121(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate3122(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate673(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate674(.a(gate429inter0), .b(s_18), .O(gate429inter1));
  and2  gate675(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate676(.a(s_18), .O(gate429inter3));
  inv1  gate677(.a(s_19), .O(gate429inter4));
  nand2 gate678(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate679(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate680(.a(G6), .O(gate429inter7));
  inv1  gate681(.a(G1147), .O(gate429inter8));
  nand2 gate682(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate683(.a(s_19), .b(gate429inter3), .O(gate429inter10));
  nor2  gate684(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate685(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate686(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate2339(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2340(.a(gate430inter0), .b(s_256), .O(gate430inter1));
  and2  gate2341(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2342(.a(s_256), .O(gate430inter3));
  inv1  gate2343(.a(s_257), .O(gate430inter4));
  nand2 gate2344(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2345(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2346(.a(G1051), .O(gate430inter7));
  inv1  gate2347(.a(G1147), .O(gate430inter8));
  nand2 gate2348(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2349(.a(s_257), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2350(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2351(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2352(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1849(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1850(.a(gate432inter0), .b(s_186), .O(gate432inter1));
  and2  gate1851(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1852(.a(s_186), .O(gate432inter3));
  inv1  gate1853(.a(s_187), .O(gate432inter4));
  nand2 gate1854(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1855(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1856(.a(G1054), .O(gate432inter7));
  inv1  gate1857(.a(G1150), .O(gate432inter8));
  nand2 gate1858(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1859(.a(s_187), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1860(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1861(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1862(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate771(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate772(.a(gate437inter0), .b(s_32), .O(gate437inter1));
  and2  gate773(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate774(.a(s_32), .O(gate437inter3));
  inv1  gate775(.a(s_33), .O(gate437inter4));
  nand2 gate776(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate777(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate778(.a(G10), .O(gate437inter7));
  inv1  gate779(.a(G1159), .O(gate437inter8));
  nand2 gate780(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate781(.a(s_33), .b(gate437inter3), .O(gate437inter10));
  nor2  gate782(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate783(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate784(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2409(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2410(.a(gate438inter0), .b(s_266), .O(gate438inter1));
  and2  gate2411(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2412(.a(s_266), .O(gate438inter3));
  inv1  gate2413(.a(s_267), .O(gate438inter4));
  nand2 gate2414(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2415(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2416(.a(G1063), .O(gate438inter7));
  inv1  gate2417(.a(G1159), .O(gate438inter8));
  nand2 gate2418(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2419(.a(s_267), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2420(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2421(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2422(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate2171(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate2172(.a(gate439inter0), .b(s_232), .O(gate439inter1));
  and2  gate2173(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate2174(.a(s_232), .O(gate439inter3));
  inv1  gate2175(.a(s_233), .O(gate439inter4));
  nand2 gate2176(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate2177(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate2178(.a(G11), .O(gate439inter7));
  inv1  gate2179(.a(G1162), .O(gate439inter8));
  nand2 gate2180(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate2181(.a(s_233), .b(gate439inter3), .O(gate439inter10));
  nor2  gate2182(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate2183(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate2184(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2269(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2270(.a(gate441inter0), .b(s_246), .O(gate441inter1));
  and2  gate2271(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2272(.a(s_246), .O(gate441inter3));
  inv1  gate2273(.a(s_247), .O(gate441inter4));
  nand2 gate2274(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2275(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2276(.a(G12), .O(gate441inter7));
  inv1  gate2277(.a(G1165), .O(gate441inter8));
  nand2 gate2278(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2279(.a(s_247), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2280(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2281(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2282(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2143(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2144(.a(gate442inter0), .b(s_228), .O(gate442inter1));
  and2  gate2145(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2146(.a(s_228), .O(gate442inter3));
  inv1  gate2147(.a(s_229), .O(gate442inter4));
  nand2 gate2148(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2149(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2150(.a(G1069), .O(gate442inter7));
  inv1  gate2151(.a(G1165), .O(gate442inter8));
  nand2 gate2152(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2153(.a(s_229), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2154(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2155(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2156(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1961(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1962(.a(gate445inter0), .b(s_202), .O(gate445inter1));
  and2  gate1963(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1964(.a(s_202), .O(gate445inter3));
  inv1  gate1965(.a(s_203), .O(gate445inter4));
  nand2 gate1966(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1967(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1968(.a(G14), .O(gate445inter7));
  inv1  gate1969(.a(G1171), .O(gate445inter8));
  nand2 gate1970(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1971(.a(s_203), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1972(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1973(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1974(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1877(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1878(.a(gate447inter0), .b(s_190), .O(gate447inter1));
  and2  gate1879(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1880(.a(s_190), .O(gate447inter3));
  inv1  gate1881(.a(s_191), .O(gate447inter4));
  nand2 gate1882(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1883(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1884(.a(G15), .O(gate447inter7));
  inv1  gate1885(.a(G1174), .O(gate447inter8));
  nand2 gate1886(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1887(.a(s_191), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1888(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1889(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1890(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2955(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2956(.a(gate448inter0), .b(s_344), .O(gate448inter1));
  and2  gate2957(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2958(.a(s_344), .O(gate448inter3));
  inv1  gate2959(.a(s_345), .O(gate448inter4));
  nand2 gate2960(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2961(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2962(.a(G1078), .O(gate448inter7));
  inv1  gate2963(.a(G1174), .O(gate448inter8));
  nand2 gate2964(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2965(.a(s_345), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2966(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2967(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2968(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2689(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2690(.a(gate449inter0), .b(s_306), .O(gate449inter1));
  and2  gate2691(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2692(.a(s_306), .O(gate449inter3));
  inv1  gate2693(.a(s_307), .O(gate449inter4));
  nand2 gate2694(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2695(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2696(.a(G16), .O(gate449inter7));
  inv1  gate2697(.a(G1177), .O(gate449inter8));
  nand2 gate2698(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2699(.a(s_307), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2700(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2701(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2702(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2297(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2298(.a(gate451inter0), .b(s_250), .O(gate451inter1));
  and2  gate2299(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2300(.a(s_250), .O(gate451inter3));
  inv1  gate2301(.a(s_251), .O(gate451inter4));
  nand2 gate2302(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2303(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2304(.a(G17), .O(gate451inter7));
  inv1  gate2305(.a(G1180), .O(gate451inter8));
  nand2 gate2306(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2307(.a(s_251), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2308(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2309(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2310(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1135(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1136(.a(gate457inter0), .b(s_84), .O(gate457inter1));
  and2  gate1137(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1138(.a(s_84), .O(gate457inter3));
  inv1  gate1139(.a(s_85), .O(gate457inter4));
  nand2 gate1140(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1141(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1142(.a(G20), .O(gate457inter7));
  inv1  gate1143(.a(G1189), .O(gate457inter8));
  nand2 gate1144(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1145(.a(s_85), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1146(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1147(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1148(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate2521(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2522(.a(gate463inter0), .b(s_282), .O(gate463inter1));
  and2  gate2523(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2524(.a(s_282), .O(gate463inter3));
  inv1  gate2525(.a(s_283), .O(gate463inter4));
  nand2 gate2526(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2527(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2528(.a(G23), .O(gate463inter7));
  inv1  gate2529(.a(G1198), .O(gate463inter8));
  nand2 gate2530(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2531(.a(s_283), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2532(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2533(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2534(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate967(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate968(.a(gate464inter0), .b(s_60), .O(gate464inter1));
  and2  gate969(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate970(.a(s_60), .O(gate464inter3));
  inv1  gate971(.a(s_61), .O(gate464inter4));
  nand2 gate972(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate973(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate974(.a(G1102), .O(gate464inter7));
  inv1  gate975(.a(G1198), .O(gate464inter8));
  nand2 gate976(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate977(.a(s_61), .b(gate464inter3), .O(gate464inter10));
  nor2  gate978(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate979(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate980(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1793(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1794(.a(gate467inter0), .b(s_178), .O(gate467inter1));
  and2  gate1795(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1796(.a(s_178), .O(gate467inter3));
  inv1  gate1797(.a(s_179), .O(gate467inter4));
  nand2 gate1798(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1799(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1800(.a(G25), .O(gate467inter7));
  inv1  gate1801(.a(G1204), .O(gate467inter8));
  nand2 gate1802(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1803(.a(s_179), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1804(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1805(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1806(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1695(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1696(.a(gate471inter0), .b(s_164), .O(gate471inter1));
  and2  gate1697(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1698(.a(s_164), .O(gate471inter3));
  inv1  gate1699(.a(s_165), .O(gate471inter4));
  nand2 gate1700(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1701(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1702(.a(G27), .O(gate471inter7));
  inv1  gate1703(.a(G1210), .O(gate471inter8));
  nand2 gate1704(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1705(.a(s_165), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1706(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1707(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1708(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1345(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1346(.a(gate473inter0), .b(s_114), .O(gate473inter1));
  and2  gate1347(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1348(.a(s_114), .O(gate473inter3));
  inv1  gate1349(.a(s_115), .O(gate473inter4));
  nand2 gate1350(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1351(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1352(.a(G28), .O(gate473inter7));
  inv1  gate1353(.a(G1213), .O(gate473inter8));
  nand2 gate1354(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1355(.a(s_115), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1356(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1357(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1358(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate827(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate828(.a(gate476inter0), .b(s_40), .O(gate476inter1));
  and2  gate829(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate830(.a(s_40), .O(gate476inter3));
  inv1  gate831(.a(s_41), .O(gate476inter4));
  nand2 gate832(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate833(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate834(.a(G1120), .O(gate476inter7));
  inv1  gate835(.a(G1216), .O(gate476inter8));
  nand2 gate836(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate837(.a(s_41), .b(gate476inter3), .O(gate476inter10));
  nor2  gate838(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate839(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate840(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1219(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1220(.a(gate478inter0), .b(s_96), .O(gate478inter1));
  and2  gate1221(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1222(.a(s_96), .O(gate478inter3));
  inv1  gate1223(.a(s_97), .O(gate478inter4));
  nand2 gate1224(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1225(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1226(.a(G1123), .O(gate478inter7));
  inv1  gate1227(.a(G1219), .O(gate478inter8));
  nand2 gate1228(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1229(.a(s_97), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1230(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1231(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1232(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1891(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1892(.a(gate479inter0), .b(s_192), .O(gate479inter1));
  and2  gate1893(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1894(.a(s_192), .O(gate479inter3));
  inv1  gate1895(.a(s_193), .O(gate479inter4));
  nand2 gate1896(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1897(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1898(.a(G31), .O(gate479inter7));
  inv1  gate1899(.a(G1222), .O(gate479inter8));
  nand2 gate1900(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1901(.a(s_193), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1902(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1903(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1904(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate2115(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2116(.a(gate480inter0), .b(s_224), .O(gate480inter1));
  and2  gate2117(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2118(.a(s_224), .O(gate480inter3));
  inv1  gate2119(.a(s_225), .O(gate480inter4));
  nand2 gate2120(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2121(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2122(.a(G1126), .O(gate480inter7));
  inv1  gate2123(.a(G1222), .O(gate480inter8));
  nand2 gate2124(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2125(.a(s_225), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2126(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2127(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2128(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate3053(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate3054(.a(gate481inter0), .b(s_358), .O(gate481inter1));
  and2  gate3055(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate3056(.a(s_358), .O(gate481inter3));
  inv1  gate3057(.a(s_359), .O(gate481inter4));
  nand2 gate3058(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate3059(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate3060(.a(G32), .O(gate481inter7));
  inv1  gate3061(.a(G1225), .O(gate481inter8));
  nand2 gate3062(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate3063(.a(s_359), .b(gate481inter3), .O(gate481inter10));
  nor2  gate3064(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate3065(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate3066(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate2381(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2382(.a(gate482inter0), .b(s_262), .O(gate482inter1));
  and2  gate2383(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2384(.a(s_262), .O(gate482inter3));
  inv1  gate2385(.a(s_263), .O(gate482inter4));
  nand2 gate2386(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2387(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2388(.a(G1129), .O(gate482inter7));
  inv1  gate2389(.a(G1225), .O(gate482inter8));
  nand2 gate2390(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2391(.a(s_263), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2392(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2393(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2394(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate785(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate786(.a(gate483inter0), .b(s_34), .O(gate483inter1));
  and2  gate787(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate788(.a(s_34), .O(gate483inter3));
  inv1  gate789(.a(s_35), .O(gate483inter4));
  nand2 gate790(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate791(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate792(.a(G1228), .O(gate483inter7));
  inv1  gate793(.a(G1229), .O(gate483inter8));
  nand2 gate794(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate795(.a(s_35), .b(gate483inter3), .O(gate483inter10));
  nor2  gate796(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate797(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate798(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2829(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2830(.a(gate485inter0), .b(s_326), .O(gate485inter1));
  and2  gate2831(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2832(.a(s_326), .O(gate485inter3));
  inv1  gate2833(.a(s_327), .O(gate485inter4));
  nand2 gate2834(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2835(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2836(.a(G1232), .O(gate485inter7));
  inv1  gate2837(.a(G1233), .O(gate485inter8));
  nand2 gate2838(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2839(.a(s_327), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2840(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2841(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2842(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate561(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate562(.a(gate487inter0), .b(s_2), .O(gate487inter1));
  and2  gate563(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate564(.a(s_2), .O(gate487inter3));
  inv1  gate565(.a(s_3), .O(gate487inter4));
  nand2 gate566(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate567(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate568(.a(G1236), .O(gate487inter7));
  inv1  gate569(.a(G1237), .O(gate487inter8));
  nand2 gate570(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate571(.a(s_3), .b(gate487inter3), .O(gate487inter10));
  nor2  gate572(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate573(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate574(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate2619(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate2620(.a(gate489inter0), .b(s_296), .O(gate489inter1));
  and2  gate2621(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate2622(.a(s_296), .O(gate489inter3));
  inv1  gate2623(.a(s_297), .O(gate489inter4));
  nand2 gate2624(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate2625(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate2626(.a(G1240), .O(gate489inter7));
  inv1  gate2627(.a(G1241), .O(gate489inter8));
  nand2 gate2628(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate2629(.a(s_297), .b(gate489inter3), .O(gate489inter10));
  nor2  gate2630(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate2631(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate2632(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate589(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate590(.a(gate492inter0), .b(s_6), .O(gate492inter1));
  and2  gate591(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate592(.a(s_6), .O(gate492inter3));
  inv1  gate593(.a(s_7), .O(gate492inter4));
  nand2 gate594(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate595(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate596(.a(G1246), .O(gate492inter7));
  inv1  gate597(.a(G1247), .O(gate492inter8));
  nand2 gate598(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate599(.a(s_7), .b(gate492inter3), .O(gate492inter10));
  nor2  gate600(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate601(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate602(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2633(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2634(.a(gate496inter0), .b(s_298), .O(gate496inter1));
  and2  gate2635(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2636(.a(s_298), .O(gate496inter3));
  inv1  gate2637(.a(s_299), .O(gate496inter4));
  nand2 gate2638(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2639(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2640(.a(G1254), .O(gate496inter7));
  inv1  gate2641(.a(G1255), .O(gate496inter8));
  nand2 gate2642(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2643(.a(s_299), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2644(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2645(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2646(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1107(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1108(.a(gate497inter0), .b(s_80), .O(gate497inter1));
  and2  gate1109(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1110(.a(s_80), .O(gate497inter3));
  inv1  gate1111(.a(s_81), .O(gate497inter4));
  nand2 gate1112(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1113(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1114(.a(G1256), .O(gate497inter7));
  inv1  gate1115(.a(G1257), .O(gate497inter8));
  nand2 gate1116(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1117(.a(s_81), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1118(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1119(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1120(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1415(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1416(.a(gate500inter0), .b(s_124), .O(gate500inter1));
  and2  gate1417(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1418(.a(s_124), .O(gate500inter3));
  inv1  gate1419(.a(s_125), .O(gate500inter4));
  nand2 gate1420(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1421(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1422(.a(G1262), .O(gate500inter7));
  inv1  gate1423(.a(G1263), .O(gate500inter8));
  nand2 gate1424(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1425(.a(s_125), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1426(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1427(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1428(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1807(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1808(.a(gate501inter0), .b(s_180), .O(gate501inter1));
  and2  gate1809(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1810(.a(s_180), .O(gate501inter3));
  inv1  gate1811(.a(s_181), .O(gate501inter4));
  nand2 gate1812(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1813(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1814(.a(G1264), .O(gate501inter7));
  inv1  gate1815(.a(G1265), .O(gate501inter8));
  nand2 gate1816(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1817(.a(s_181), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1818(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1819(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1820(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2255(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2256(.a(gate502inter0), .b(s_244), .O(gate502inter1));
  and2  gate2257(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2258(.a(s_244), .O(gate502inter3));
  inv1  gate2259(.a(s_245), .O(gate502inter4));
  nand2 gate2260(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2261(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2262(.a(G1266), .O(gate502inter7));
  inv1  gate2263(.a(G1267), .O(gate502inter8));
  nand2 gate2264(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2265(.a(s_245), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2266(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2267(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2268(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2787(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2788(.a(gate503inter0), .b(s_320), .O(gate503inter1));
  and2  gate2789(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2790(.a(s_320), .O(gate503inter3));
  inv1  gate2791(.a(s_321), .O(gate503inter4));
  nand2 gate2792(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2793(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2794(.a(G1268), .O(gate503inter7));
  inv1  gate2795(.a(G1269), .O(gate503inter8));
  nand2 gate2796(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2797(.a(s_321), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2798(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2799(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2800(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2969(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2970(.a(gate507inter0), .b(s_346), .O(gate507inter1));
  and2  gate2971(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2972(.a(s_346), .O(gate507inter3));
  inv1  gate2973(.a(s_347), .O(gate507inter4));
  nand2 gate2974(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2975(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2976(.a(G1276), .O(gate507inter7));
  inv1  gate2977(.a(G1277), .O(gate507inter8));
  nand2 gate2978(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2979(.a(s_347), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2980(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2981(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2982(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1149(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1150(.a(gate509inter0), .b(s_86), .O(gate509inter1));
  and2  gate1151(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1152(.a(s_86), .O(gate509inter3));
  inv1  gate1153(.a(s_87), .O(gate509inter4));
  nand2 gate1154(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1155(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1156(.a(G1280), .O(gate509inter7));
  inv1  gate1157(.a(G1281), .O(gate509inter8));
  nand2 gate1158(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1159(.a(s_87), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1160(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1161(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1162(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate3039(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate3040(.a(gate513inter0), .b(s_356), .O(gate513inter1));
  and2  gate3041(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate3042(.a(s_356), .O(gate513inter3));
  inv1  gate3043(.a(s_357), .O(gate513inter4));
  nand2 gate3044(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate3045(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate3046(.a(G1288), .O(gate513inter7));
  inv1  gate3047(.a(G1289), .O(gate513inter8));
  nand2 gate3048(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate3049(.a(s_357), .b(gate513inter3), .O(gate513inter10));
  nor2  gate3050(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate3051(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate3052(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule