module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1163(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1164(.a(gate9inter0), .b(s_88), .O(gate9inter1));
  and2  gate1165(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1166(.a(s_88), .O(gate9inter3));
  inv1  gate1167(.a(s_89), .O(gate9inter4));
  nand2 gate1168(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1169(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1170(.a(G1), .O(gate9inter7));
  inv1  gate1171(.a(G2), .O(gate9inter8));
  nand2 gate1172(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1173(.a(s_89), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1174(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1175(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1176(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate827(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate828(.a(gate15inter0), .b(s_40), .O(gate15inter1));
  and2  gate829(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate830(.a(s_40), .O(gate15inter3));
  inv1  gate831(.a(s_41), .O(gate15inter4));
  nand2 gate832(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate833(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate834(.a(G13), .O(gate15inter7));
  inv1  gate835(.a(G14), .O(gate15inter8));
  nand2 gate836(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate837(.a(s_41), .b(gate15inter3), .O(gate15inter10));
  nor2  gate838(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate839(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate840(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate855(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate856(.a(gate16inter0), .b(s_44), .O(gate16inter1));
  and2  gate857(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate858(.a(s_44), .O(gate16inter3));
  inv1  gate859(.a(s_45), .O(gate16inter4));
  nand2 gate860(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate861(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate862(.a(G15), .O(gate16inter7));
  inv1  gate863(.a(G16), .O(gate16inter8));
  nand2 gate864(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate865(.a(s_45), .b(gate16inter3), .O(gate16inter10));
  nor2  gate866(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate867(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate868(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1359(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1360(.a(gate17inter0), .b(s_116), .O(gate17inter1));
  and2  gate1361(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1362(.a(s_116), .O(gate17inter3));
  inv1  gate1363(.a(s_117), .O(gate17inter4));
  nand2 gate1364(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1365(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1366(.a(G17), .O(gate17inter7));
  inv1  gate1367(.a(G18), .O(gate17inter8));
  nand2 gate1368(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1369(.a(s_117), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1370(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1371(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1372(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1135(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1136(.a(gate26inter0), .b(s_84), .O(gate26inter1));
  and2  gate1137(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1138(.a(s_84), .O(gate26inter3));
  inv1  gate1139(.a(s_85), .O(gate26inter4));
  nand2 gate1140(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1141(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1142(.a(G9), .O(gate26inter7));
  inv1  gate1143(.a(G13), .O(gate26inter8));
  nand2 gate1144(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1145(.a(s_85), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1146(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1147(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1148(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1317(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1318(.a(gate41inter0), .b(s_110), .O(gate41inter1));
  and2  gate1319(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1320(.a(s_110), .O(gate41inter3));
  inv1  gate1321(.a(s_111), .O(gate41inter4));
  nand2 gate1322(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1323(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1324(.a(G1), .O(gate41inter7));
  inv1  gate1325(.a(G266), .O(gate41inter8));
  nand2 gate1326(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1327(.a(s_111), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1328(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1329(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1330(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate575(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate576(.a(gate65inter0), .b(s_4), .O(gate65inter1));
  and2  gate577(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate578(.a(s_4), .O(gate65inter3));
  inv1  gate579(.a(s_5), .O(gate65inter4));
  nand2 gate580(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate581(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate582(.a(G25), .O(gate65inter7));
  inv1  gate583(.a(G302), .O(gate65inter8));
  nand2 gate584(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate585(.a(s_5), .b(gate65inter3), .O(gate65inter10));
  nor2  gate586(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate587(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate588(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate617(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate618(.a(gate71inter0), .b(s_10), .O(gate71inter1));
  and2  gate619(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate620(.a(s_10), .O(gate71inter3));
  inv1  gate621(.a(s_11), .O(gate71inter4));
  nand2 gate622(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate623(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate624(.a(G31), .O(gate71inter7));
  inv1  gate625(.a(G311), .O(gate71inter8));
  nand2 gate626(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate627(.a(s_11), .b(gate71inter3), .O(gate71inter10));
  nor2  gate628(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate629(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate630(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1457(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1458(.a(gate74inter0), .b(s_130), .O(gate74inter1));
  and2  gate1459(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1460(.a(s_130), .O(gate74inter3));
  inv1  gate1461(.a(s_131), .O(gate74inter4));
  nand2 gate1462(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1463(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1464(.a(G5), .O(gate74inter7));
  inv1  gate1465(.a(G314), .O(gate74inter8));
  nand2 gate1466(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1467(.a(s_131), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1468(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1469(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1470(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1345(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1346(.a(gate75inter0), .b(s_114), .O(gate75inter1));
  and2  gate1347(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1348(.a(s_114), .O(gate75inter3));
  inv1  gate1349(.a(s_115), .O(gate75inter4));
  nand2 gate1350(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1351(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1352(.a(G9), .O(gate75inter7));
  inv1  gate1353(.a(G317), .O(gate75inter8));
  nand2 gate1354(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1355(.a(s_115), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1356(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1357(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1358(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1149(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1150(.a(gate81inter0), .b(s_86), .O(gate81inter1));
  and2  gate1151(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1152(.a(s_86), .O(gate81inter3));
  inv1  gate1153(.a(s_87), .O(gate81inter4));
  nand2 gate1154(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1155(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1156(.a(G3), .O(gate81inter7));
  inv1  gate1157(.a(G326), .O(gate81inter8));
  nand2 gate1158(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1159(.a(s_87), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1160(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1161(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1162(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate673(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate674(.a(gate86inter0), .b(s_18), .O(gate86inter1));
  and2  gate675(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate676(.a(s_18), .O(gate86inter3));
  inv1  gate677(.a(s_19), .O(gate86inter4));
  nand2 gate678(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate679(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate680(.a(G8), .O(gate86inter7));
  inv1  gate681(.a(G332), .O(gate86inter8));
  nand2 gate682(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate683(.a(s_19), .b(gate86inter3), .O(gate86inter10));
  nor2  gate684(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate685(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate686(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1443(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1444(.a(gate109inter0), .b(s_128), .O(gate109inter1));
  and2  gate1445(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1446(.a(s_128), .O(gate109inter3));
  inv1  gate1447(.a(s_129), .O(gate109inter4));
  nand2 gate1448(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1449(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1450(.a(G370), .O(gate109inter7));
  inv1  gate1451(.a(G371), .O(gate109inter8));
  nand2 gate1452(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1453(.a(s_129), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1454(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1455(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1456(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1177(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1178(.a(gate115inter0), .b(s_90), .O(gate115inter1));
  and2  gate1179(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1180(.a(s_90), .O(gate115inter3));
  inv1  gate1181(.a(s_91), .O(gate115inter4));
  nand2 gate1182(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1183(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1184(.a(G382), .O(gate115inter7));
  inv1  gate1185(.a(G383), .O(gate115inter8));
  nand2 gate1186(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1187(.a(s_91), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1188(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1189(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1190(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate785(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate786(.a(gate118inter0), .b(s_34), .O(gate118inter1));
  and2  gate787(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate788(.a(s_34), .O(gate118inter3));
  inv1  gate789(.a(s_35), .O(gate118inter4));
  nand2 gate790(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate791(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate792(.a(G388), .O(gate118inter7));
  inv1  gate793(.a(G389), .O(gate118inter8));
  nand2 gate794(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate795(.a(s_35), .b(gate118inter3), .O(gate118inter10));
  nor2  gate796(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate797(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate798(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1051(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1052(.a(gate143inter0), .b(s_72), .O(gate143inter1));
  and2  gate1053(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1054(.a(s_72), .O(gate143inter3));
  inv1  gate1055(.a(s_73), .O(gate143inter4));
  nand2 gate1056(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1057(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1058(.a(G462), .O(gate143inter7));
  inv1  gate1059(.a(G465), .O(gate143inter8));
  nand2 gate1060(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1061(.a(s_73), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1062(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1063(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1064(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1261(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1262(.a(gate144inter0), .b(s_102), .O(gate144inter1));
  and2  gate1263(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1264(.a(s_102), .O(gate144inter3));
  inv1  gate1265(.a(s_103), .O(gate144inter4));
  nand2 gate1266(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1267(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1268(.a(G468), .O(gate144inter7));
  inv1  gate1269(.a(G471), .O(gate144inter8));
  nand2 gate1270(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1271(.a(s_103), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1272(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1273(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1274(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1191(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1192(.a(gate147inter0), .b(s_92), .O(gate147inter1));
  and2  gate1193(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1194(.a(s_92), .O(gate147inter3));
  inv1  gate1195(.a(s_93), .O(gate147inter4));
  nand2 gate1196(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1197(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1198(.a(G486), .O(gate147inter7));
  inv1  gate1199(.a(G489), .O(gate147inter8));
  nand2 gate1200(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1201(.a(s_93), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1202(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1203(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1204(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate547(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate548(.a(gate155inter0), .b(s_0), .O(gate155inter1));
  and2  gate549(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate550(.a(s_0), .O(gate155inter3));
  inv1  gate551(.a(s_1), .O(gate155inter4));
  nand2 gate552(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate553(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate554(.a(G432), .O(gate155inter7));
  inv1  gate555(.a(G525), .O(gate155inter8));
  nand2 gate556(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate557(.a(s_1), .b(gate155inter3), .O(gate155inter10));
  nor2  gate558(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate559(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate560(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate603(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate604(.a(gate167inter0), .b(s_8), .O(gate167inter1));
  and2  gate605(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate606(.a(s_8), .O(gate167inter3));
  inv1  gate607(.a(s_9), .O(gate167inter4));
  nand2 gate608(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate609(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate610(.a(G468), .O(gate167inter7));
  inv1  gate611(.a(G543), .O(gate167inter8));
  nand2 gate612(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate613(.a(s_9), .b(gate167inter3), .O(gate167inter10));
  nor2  gate614(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate615(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate616(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1219(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1220(.a(gate170inter0), .b(s_96), .O(gate170inter1));
  and2  gate1221(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1222(.a(s_96), .O(gate170inter3));
  inv1  gate1223(.a(s_97), .O(gate170inter4));
  nand2 gate1224(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1225(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1226(.a(G477), .O(gate170inter7));
  inv1  gate1227(.a(G546), .O(gate170inter8));
  nand2 gate1228(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1229(.a(s_97), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1230(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1231(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1232(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate589(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate590(.a(gate177inter0), .b(s_6), .O(gate177inter1));
  and2  gate591(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate592(.a(s_6), .O(gate177inter3));
  inv1  gate593(.a(s_7), .O(gate177inter4));
  nand2 gate594(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate595(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate596(.a(G498), .O(gate177inter7));
  inv1  gate597(.a(G558), .O(gate177inter8));
  nand2 gate598(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate599(.a(s_7), .b(gate177inter3), .O(gate177inter10));
  nor2  gate600(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate601(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate602(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate911(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate912(.a(gate178inter0), .b(s_52), .O(gate178inter1));
  and2  gate913(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate914(.a(s_52), .O(gate178inter3));
  inv1  gate915(.a(s_53), .O(gate178inter4));
  nand2 gate916(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate917(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate918(.a(G501), .O(gate178inter7));
  inv1  gate919(.a(G558), .O(gate178inter8));
  nand2 gate920(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate921(.a(s_53), .b(gate178inter3), .O(gate178inter10));
  nor2  gate922(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate923(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate924(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate1387(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1388(.a(gate179inter0), .b(s_120), .O(gate179inter1));
  and2  gate1389(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1390(.a(s_120), .O(gate179inter3));
  inv1  gate1391(.a(s_121), .O(gate179inter4));
  nand2 gate1392(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1393(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1394(.a(G504), .O(gate179inter7));
  inv1  gate1395(.a(G561), .O(gate179inter8));
  nand2 gate1396(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1397(.a(s_121), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1398(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1399(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1400(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1415(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1416(.a(gate188inter0), .b(s_124), .O(gate188inter1));
  and2  gate1417(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1418(.a(s_124), .O(gate188inter3));
  inv1  gate1419(.a(s_125), .O(gate188inter4));
  nand2 gate1420(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1421(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1422(.a(G576), .O(gate188inter7));
  inv1  gate1423(.a(G577), .O(gate188inter8));
  nand2 gate1424(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1425(.a(s_125), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1426(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1427(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1428(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate939(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate940(.a(gate189inter0), .b(s_56), .O(gate189inter1));
  and2  gate941(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate942(.a(s_56), .O(gate189inter3));
  inv1  gate943(.a(s_57), .O(gate189inter4));
  nand2 gate944(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate945(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate946(.a(G578), .O(gate189inter7));
  inv1  gate947(.a(G579), .O(gate189inter8));
  nand2 gate948(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate949(.a(s_57), .b(gate189inter3), .O(gate189inter10));
  nor2  gate950(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate951(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate952(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate841(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate842(.a(gate205inter0), .b(s_42), .O(gate205inter1));
  and2  gate843(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate844(.a(s_42), .O(gate205inter3));
  inv1  gate845(.a(s_43), .O(gate205inter4));
  nand2 gate846(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate847(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate848(.a(G622), .O(gate205inter7));
  inv1  gate849(.a(G627), .O(gate205inter8));
  nand2 gate850(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate851(.a(s_43), .b(gate205inter3), .O(gate205inter10));
  nor2  gate852(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate853(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate854(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate701(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate702(.a(gate208inter0), .b(s_22), .O(gate208inter1));
  and2  gate703(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate704(.a(s_22), .O(gate208inter3));
  inv1  gate705(.a(s_23), .O(gate208inter4));
  nand2 gate706(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate707(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate708(.a(G627), .O(gate208inter7));
  inv1  gate709(.a(G637), .O(gate208inter8));
  nand2 gate710(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate711(.a(s_23), .b(gate208inter3), .O(gate208inter10));
  nor2  gate712(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate713(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate714(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1093(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1094(.a(gate211inter0), .b(s_78), .O(gate211inter1));
  and2  gate1095(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1096(.a(s_78), .O(gate211inter3));
  inv1  gate1097(.a(s_79), .O(gate211inter4));
  nand2 gate1098(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1099(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1100(.a(G612), .O(gate211inter7));
  inv1  gate1101(.a(G669), .O(gate211inter8));
  nand2 gate1102(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1103(.a(s_79), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1104(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1105(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1106(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1275(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1276(.a(gate223inter0), .b(s_104), .O(gate223inter1));
  and2  gate1277(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1278(.a(s_104), .O(gate223inter3));
  inv1  gate1279(.a(s_105), .O(gate223inter4));
  nand2 gate1280(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1281(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1282(.a(G627), .O(gate223inter7));
  inv1  gate1283(.a(G687), .O(gate223inter8));
  nand2 gate1284(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1285(.a(s_105), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1286(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1287(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1288(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate715(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate716(.a(gate224inter0), .b(s_24), .O(gate224inter1));
  and2  gate717(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate718(.a(s_24), .O(gate224inter3));
  inv1  gate719(.a(s_25), .O(gate224inter4));
  nand2 gate720(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate721(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate722(.a(G637), .O(gate224inter7));
  inv1  gate723(.a(G687), .O(gate224inter8));
  nand2 gate724(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate725(.a(s_25), .b(gate224inter3), .O(gate224inter10));
  nor2  gate726(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate727(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate728(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate757(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate758(.a(gate227inter0), .b(s_30), .O(gate227inter1));
  and2  gate759(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate760(.a(s_30), .O(gate227inter3));
  inv1  gate761(.a(s_31), .O(gate227inter4));
  nand2 gate762(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate763(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate764(.a(G694), .O(gate227inter7));
  inv1  gate765(.a(G695), .O(gate227inter8));
  nand2 gate766(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate767(.a(s_31), .b(gate227inter3), .O(gate227inter10));
  nor2  gate768(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate769(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate770(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate729(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate730(.a(gate228inter0), .b(s_26), .O(gate228inter1));
  and2  gate731(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate732(.a(s_26), .O(gate228inter3));
  inv1  gate733(.a(s_27), .O(gate228inter4));
  nand2 gate734(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate735(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate736(.a(G696), .O(gate228inter7));
  inv1  gate737(.a(G697), .O(gate228inter8));
  nand2 gate738(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate739(.a(s_27), .b(gate228inter3), .O(gate228inter10));
  nor2  gate740(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate741(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate742(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1331(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1332(.a(gate229inter0), .b(s_112), .O(gate229inter1));
  and2  gate1333(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1334(.a(s_112), .O(gate229inter3));
  inv1  gate1335(.a(s_113), .O(gate229inter4));
  nand2 gate1336(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1337(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1338(.a(G698), .O(gate229inter7));
  inv1  gate1339(.a(G699), .O(gate229inter8));
  nand2 gate1340(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1341(.a(s_113), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1342(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1343(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1344(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1429(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1430(.a(gate235inter0), .b(s_126), .O(gate235inter1));
  and2  gate1431(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1432(.a(s_126), .O(gate235inter3));
  inv1  gate1433(.a(s_127), .O(gate235inter4));
  nand2 gate1434(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1435(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1436(.a(G248), .O(gate235inter7));
  inv1  gate1437(.a(G724), .O(gate235inter8));
  nand2 gate1438(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1439(.a(s_127), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1440(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1441(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1442(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate771(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate772(.a(gate238inter0), .b(s_32), .O(gate238inter1));
  and2  gate773(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate774(.a(s_32), .O(gate238inter3));
  inv1  gate775(.a(s_33), .O(gate238inter4));
  nand2 gate776(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate777(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate778(.a(G257), .O(gate238inter7));
  inv1  gate779(.a(G709), .O(gate238inter8));
  nand2 gate780(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate781(.a(s_33), .b(gate238inter3), .O(gate238inter10));
  nor2  gate782(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate783(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate784(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1205(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1206(.a(gate240inter0), .b(s_94), .O(gate240inter1));
  and2  gate1207(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1208(.a(s_94), .O(gate240inter3));
  inv1  gate1209(.a(s_95), .O(gate240inter4));
  nand2 gate1210(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1211(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1212(.a(G263), .O(gate240inter7));
  inv1  gate1213(.a(G715), .O(gate240inter8));
  nand2 gate1214(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1215(.a(s_95), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1216(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1217(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1218(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1065(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1066(.a(gate257inter0), .b(s_74), .O(gate257inter1));
  and2  gate1067(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1068(.a(s_74), .O(gate257inter3));
  inv1  gate1069(.a(s_75), .O(gate257inter4));
  nand2 gate1070(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1071(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1072(.a(G754), .O(gate257inter7));
  inv1  gate1073(.a(G755), .O(gate257inter8));
  nand2 gate1074(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1075(.a(s_75), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1076(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1077(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1078(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1107(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1108(.a(gate260inter0), .b(s_80), .O(gate260inter1));
  and2  gate1109(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1110(.a(s_80), .O(gate260inter3));
  inv1  gate1111(.a(s_81), .O(gate260inter4));
  nand2 gate1112(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1113(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1114(.a(G760), .O(gate260inter7));
  inv1  gate1115(.a(G761), .O(gate260inter8));
  nand2 gate1116(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1117(.a(s_81), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1118(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1119(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1120(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate687(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate688(.a(gate263inter0), .b(s_20), .O(gate263inter1));
  and2  gate689(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate690(.a(s_20), .O(gate263inter3));
  inv1  gate691(.a(s_21), .O(gate263inter4));
  nand2 gate692(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate693(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate694(.a(G766), .O(gate263inter7));
  inv1  gate695(.a(G767), .O(gate263inter8));
  nand2 gate696(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate697(.a(s_21), .b(gate263inter3), .O(gate263inter10));
  nor2  gate698(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate699(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate700(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1037(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1038(.a(gate269inter0), .b(s_70), .O(gate269inter1));
  and2  gate1039(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1040(.a(s_70), .O(gate269inter3));
  inv1  gate1041(.a(s_71), .O(gate269inter4));
  nand2 gate1042(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1043(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1044(.a(G654), .O(gate269inter7));
  inv1  gate1045(.a(G782), .O(gate269inter8));
  nand2 gate1046(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1047(.a(s_71), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1048(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1049(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1050(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate869(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate870(.a(gate273inter0), .b(s_46), .O(gate273inter1));
  and2  gate871(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate872(.a(s_46), .O(gate273inter3));
  inv1  gate873(.a(s_47), .O(gate273inter4));
  nand2 gate874(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate875(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate876(.a(G642), .O(gate273inter7));
  inv1  gate877(.a(G794), .O(gate273inter8));
  nand2 gate878(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate879(.a(s_47), .b(gate273inter3), .O(gate273inter10));
  nor2  gate880(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate881(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate882(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate799(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate800(.a(gate276inter0), .b(s_36), .O(gate276inter1));
  and2  gate801(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate802(.a(s_36), .O(gate276inter3));
  inv1  gate803(.a(s_37), .O(gate276inter4));
  nand2 gate804(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate805(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate806(.a(G773), .O(gate276inter7));
  inv1  gate807(.a(G797), .O(gate276inter8));
  nand2 gate808(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate809(.a(s_37), .b(gate276inter3), .O(gate276inter10));
  nor2  gate810(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate811(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate812(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate953(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate954(.a(gate277inter0), .b(s_58), .O(gate277inter1));
  and2  gate955(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate956(.a(s_58), .O(gate277inter3));
  inv1  gate957(.a(s_59), .O(gate277inter4));
  nand2 gate958(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate959(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate960(.a(G648), .O(gate277inter7));
  inv1  gate961(.a(G800), .O(gate277inter8));
  nand2 gate962(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate963(.a(s_59), .b(gate277inter3), .O(gate277inter10));
  nor2  gate964(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate965(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate966(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate995(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate996(.a(gate289inter0), .b(s_64), .O(gate289inter1));
  and2  gate997(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate998(.a(s_64), .O(gate289inter3));
  inv1  gate999(.a(s_65), .O(gate289inter4));
  nand2 gate1000(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1001(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1002(.a(G818), .O(gate289inter7));
  inv1  gate1003(.a(G819), .O(gate289inter8));
  nand2 gate1004(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1005(.a(s_65), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1006(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1007(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1008(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1303(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1304(.a(gate290inter0), .b(s_108), .O(gate290inter1));
  and2  gate1305(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1306(.a(s_108), .O(gate290inter3));
  inv1  gate1307(.a(s_109), .O(gate290inter4));
  nand2 gate1308(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1309(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1310(.a(G820), .O(gate290inter7));
  inv1  gate1311(.a(G821), .O(gate290inter8));
  nand2 gate1312(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1313(.a(s_109), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1314(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1315(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1316(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate631(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate632(.a(gate387inter0), .b(s_12), .O(gate387inter1));
  and2  gate633(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate634(.a(s_12), .O(gate387inter3));
  inv1  gate635(.a(s_13), .O(gate387inter4));
  nand2 gate636(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate637(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate638(.a(G1), .O(gate387inter7));
  inv1  gate639(.a(G1036), .O(gate387inter8));
  nand2 gate640(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate641(.a(s_13), .b(gate387inter3), .O(gate387inter10));
  nor2  gate642(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate643(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate644(.a(gate387inter12), .b(gate387inter1), .O(G1132));

  xor2  gate1009(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1010(.a(gate388inter0), .b(s_66), .O(gate388inter1));
  and2  gate1011(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1012(.a(s_66), .O(gate388inter3));
  inv1  gate1013(.a(s_67), .O(gate388inter4));
  nand2 gate1014(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1015(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1016(.a(G2), .O(gate388inter7));
  inv1  gate1017(.a(G1039), .O(gate388inter8));
  nand2 gate1018(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1019(.a(s_67), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1020(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1021(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1022(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate967(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate968(.a(gate399inter0), .b(s_60), .O(gate399inter1));
  and2  gate969(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate970(.a(s_60), .O(gate399inter3));
  inv1  gate971(.a(s_61), .O(gate399inter4));
  nand2 gate972(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate973(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate974(.a(G13), .O(gate399inter7));
  inv1  gate975(.a(G1072), .O(gate399inter8));
  nand2 gate976(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate977(.a(s_61), .b(gate399inter3), .O(gate399inter10));
  nor2  gate978(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate979(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate980(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1289(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1290(.a(gate412inter0), .b(s_106), .O(gate412inter1));
  and2  gate1291(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1292(.a(s_106), .O(gate412inter3));
  inv1  gate1293(.a(s_107), .O(gate412inter4));
  nand2 gate1294(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1295(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1296(.a(G26), .O(gate412inter7));
  inv1  gate1297(.a(G1111), .O(gate412inter8));
  nand2 gate1298(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1299(.a(s_107), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1300(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1301(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1302(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1079(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1080(.a(gate415inter0), .b(s_76), .O(gate415inter1));
  and2  gate1081(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1082(.a(s_76), .O(gate415inter3));
  inv1  gate1083(.a(s_77), .O(gate415inter4));
  nand2 gate1084(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1085(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1086(.a(G29), .O(gate415inter7));
  inv1  gate1087(.a(G1120), .O(gate415inter8));
  nand2 gate1088(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1089(.a(s_77), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1090(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1091(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1092(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate645(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate646(.a(gate429inter0), .b(s_14), .O(gate429inter1));
  and2  gate647(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate648(.a(s_14), .O(gate429inter3));
  inv1  gate649(.a(s_15), .O(gate429inter4));
  nand2 gate650(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate651(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate652(.a(G6), .O(gate429inter7));
  inv1  gate653(.a(G1147), .O(gate429inter8));
  nand2 gate654(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate655(.a(s_15), .b(gate429inter3), .O(gate429inter10));
  nor2  gate656(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate657(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate658(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate883(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate884(.a(gate432inter0), .b(s_48), .O(gate432inter1));
  and2  gate885(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate886(.a(s_48), .O(gate432inter3));
  inv1  gate887(.a(s_49), .O(gate432inter4));
  nand2 gate888(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate889(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate890(.a(G1054), .O(gate432inter7));
  inv1  gate891(.a(G1150), .O(gate432inter8));
  nand2 gate892(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate893(.a(s_49), .b(gate432inter3), .O(gate432inter10));
  nor2  gate894(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate895(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate896(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate813(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate814(.a(gate451inter0), .b(s_38), .O(gate451inter1));
  and2  gate815(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate816(.a(s_38), .O(gate451inter3));
  inv1  gate817(.a(s_39), .O(gate451inter4));
  nand2 gate818(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate819(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate820(.a(G17), .O(gate451inter7));
  inv1  gate821(.a(G1180), .O(gate451inter8));
  nand2 gate822(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate823(.a(s_39), .b(gate451inter3), .O(gate451inter10));
  nor2  gate824(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate825(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate826(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate743(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate744(.a(gate463inter0), .b(s_28), .O(gate463inter1));
  and2  gate745(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate746(.a(s_28), .O(gate463inter3));
  inv1  gate747(.a(s_29), .O(gate463inter4));
  nand2 gate748(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate749(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate750(.a(G23), .O(gate463inter7));
  inv1  gate751(.a(G1198), .O(gate463inter8));
  nand2 gate752(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate753(.a(s_29), .b(gate463inter3), .O(gate463inter10));
  nor2  gate754(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate755(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate756(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate981(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate982(.a(gate476inter0), .b(s_62), .O(gate476inter1));
  and2  gate983(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate984(.a(s_62), .O(gate476inter3));
  inv1  gate985(.a(s_63), .O(gate476inter4));
  nand2 gate986(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate987(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate988(.a(G1120), .O(gate476inter7));
  inv1  gate989(.a(G1216), .O(gate476inter8));
  nand2 gate990(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate991(.a(s_63), .b(gate476inter3), .O(gate476inter10));
  nor2  gate992(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate993(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate994(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1121(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1122(.a(gate482inter0), .b(s_82), .O(gate482inter1));
  and2  gate1123(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1124(.a(s_82), .O(gate482inter3));
  inv1  gate1125(.a(s_83), .O(gate482inter4));
  nand2 gate1126(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1127(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1128(.a(G1129), .O(gate482inter7));
  inv1  gate1129(.a(G1225), .O(gate482inter8));
  nand2 gate1130(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1131(.a(s_83), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1132(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1133(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1134(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1401(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1402(.a(gate483inter0), .b(s_122), .O(gate483inter1));
  and2  gate1403(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1404(.a(s_122), .O(gate483inter3));
  inv1  gate1405(.a(s_123), .O(gate483inter4));
  nand2 gate1406(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1407(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1408(.a(G1228), .O(gate483inter7));
  inv1  gate1409(.a(G1229), .O(gate483inter8));
  nand2 gate1410(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1411(.a(s_123), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1412(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1413(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1414(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate561(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate562(.a(gate486inter0), .b(s_2), .O(gate486inter1));
  and2  gate563(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate564(.a(s_2), .O(gate486inter3));
  inv1  gate565(.a(s_3), .O(gate486inter4));
  nand2 gate566(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate567(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate568(.a(G1234), .O(gate486inter7));
  inv1  gate569(.a(G1235), .O(gate486inter8));
  nand2 gate570(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate571(.a(s_3), .b(gate486inter3), .O(gate486inter10));
  nor2  gate572(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate573(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate574(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1373(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1374(.a(gate490inter0), .b(s_118), .O(gate490inter1));
  and2  gate1375(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1376(.a(s_118), .O(gate490inter3));
  inv1  gate1377(.a(s_119), .O(gate490inter4));
  nand2 gate1378(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1379(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1380(.a(G1242), .O(gate490inter7));
  inv1  gate1381(.a(G1243), .O(gate490inter8));
  nand2 gate1382(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1383(.a(s_119), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1384(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1385(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1386(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1247(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1248(.a(gate494inter0), .b(s_100), .O(gate494inter1));
  and2  gate1249(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1250(.a(s_100), .O(gate494inter3));
  inv1  gate1251(.a(s_101), .O(gate494inter4));
  nand2 gate1252(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1253(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1254(.a(G1250), .O(gate494inter7));
  inv1  gate1255(.a(G1251), .O(gate494inter8));
  nand2 gate1256(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1257(.a(s_101), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1258(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1259(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1260(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1023(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1024(.a(gate495inter0), .b(s_68), .O(gate495inter1));
  and2  gate1025(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1026(.a(s_68), .O(gate495inter3));
  inv1  gate1027(.a(s_69), .O(gate495inter4));
  nand2 gate1028(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1029(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1030(.a(G1252), .O(gate495inter7));
  inv1  gate1031(.a(G1253), .O(gate495inter8));
  nand2 gate1032(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1033(.a(s_69), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1034(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1035(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1036(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate925(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate926(.a(gate498inter0), .b(s_54), .O(gate498inter1));
  and2  gate927(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate928(.a(s_54), .O(gate498inter3));
  inv1  gate929(.a(s_55), .O(gate498inter4));
  nand2 gate930(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate931(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate932(.a(G1258), .O(gate498inter7));
  inv1  gate933(.a(G1259), .O(gate498inter8));
  nand2 gate934(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate935(.a(s_55), .b(gate498inter3), .O(gate498inter10));
  nor2  gate936(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate937(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate938(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1233(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1234(.a(gate499inter0), .b(s_98), .O(gate499inter1));
  and2  gate1235(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1236(.a(s_98), .O(gate499inter3));
  inv1  gate1237(.a(s_99), .O(gate499inter4));
  nand2 gate1238(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1239(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1240(.a(G1260), .O(gate499inter7));
  inv1  gate1241(.a(G1261), .O(gate499inter8));
  nand2 gate1242(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1243(.a(s_99), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1244(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1245(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1246(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate897(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate898(.a(gate506inter0), .b(s_50), .O(gate506inter1));
  and2  gate899(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate900(.a(s_50), .O(gate506inter3));
  inv1  gate901(.a(s_51), .O(gate506inter4));
  nand2 gate902(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate903(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate904(.a(G1274), .O(gate506inter7));
  inv1  gate905(.a(G1275), .O(gate506inter8));
  nand2 gate906(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate907(.a(s_51), .b(gate506inter3), .O(gate506inter10));
  nor2  gate908(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate909(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate910(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate659(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate660(.a(gate510inter0), .b(s_16), .O(gate510inter1));
  and2  gate661(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate662(.a(s_16), .O(gate510inter3));
  inv1  gate663(.a(s_17), .O(gate510inter4));
  nand2 gate664(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate665(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate666(.a(G1282), .O(gate510inter7));
  inv1  gate667(.a(G1283), .O(gate510inter8));
  nand2 gate668(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate669(.a(s_17), .b(gate510inter3), .O(gate510inter10));
  nor2  gate670(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate671(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate672(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule