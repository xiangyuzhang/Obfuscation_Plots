module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate7inter0, gate7inter1, gate7inter2, gate7inter3, gate7inter4, gate7inter5, gate7inter6, gate7inter7, gate7inter8, gate7inter9, gate7inter10, gate7inter11, gate7inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate5inter0, gate5inter1, gate5inter2, gate5inter3, gate5inter4, gate5inter5, gate5inter6, gate5inter7, gate5inter8, gate5inter9, gate5inter10, gate5inter11, gate5inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );

  xor2  gate539(.a(N37), .b(N33), .O(gate5inter0));
  nand2 gate540(.a(gate5inter0), .b(s_48), .O(gate5inter1));
  and2  gate541(.a(N37), .b(N33), .O(gate5inter2));
  inv1  gate542(.a(s_48), .O(gate5inter3));
  inv1  gate543(.a(s_49), .O(gate5inter4));
  nand2 gate544(.a(gate5inter4), .b(gate5inter3), .O(gate5inter5));
  nor2  gate545(.a(gate5inter5), .b(gate5inter2), .O(gate5inter6));
  inv1  gate546(.a(N33), .O(gate5inter7));
  inv1  gate547(.a(N37), .O(gate5inter8));
  nand2 gate548(.a(gate5inter8), .b(gate5inter7), .O(gate5inter9));
  nand2 gate549(.a(s_49), .b(gate5inter3), .O(gate5inter10));
  nor2  gate550(.a(gate5inter10), .b(gate5inter9), .O(gate5inter11));
  nor2  gate551(.a(gate5inter11), .b(gate5inter6), .O(gate5inter12));
  nand2 gate552(.a(gate5inter12), .b(gate5inter1), .O(N254));
xor2 gate6( .a(N41), .b(N45), .O(N255) );

  xor2  gate301(.a(N53), .b(N49), .O(gate7inter0));
  nand2 gate302(.a(gate7inter0), .b(s_14), .O(gate7inter1));
  and2  gate303(.a(N53), .b(N49), .O(gate7inter2));
  inv1  gate304(.a(s_14), .O(gate7inter3));
  inv1  gate305(.a(s_15), .O(gate7inter4));
  nand2 gate306(.a(gate7inter4), .b(gate7inter3), .O(gate7inter5));
  nor2  gate307(.a(gate7inter5), .b(gate7inter2), .O(gate7inter6));
  inv1  gate308(.a(N49), .O(gate7inter7));
  inv1  gate309(.a(N53), .O(gate7inter8));
  nand2 gate310(.a(gate7inter8), .b(gate7inter7), .O(gate7inter9));
  nand2 gate311(.a(s_15), .b(gate7inter3), .O(gate7inter10));
  nor2  gate312(.a(gate7inter10), .b(gate7inter9), .O(gate7inter11));
  nor2  gate313(.a(gate7inter11), .b(gate7inter6), .O(gate7inter12));
  nand2 gate314(.a(gate7inter12), .b(gate7inter1), .O(N256));
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );

  xor2  gate245(.a(N77), .b(N73), .O(gate10inter0));
  nand2 gate246(.a(gate10inter0), .b(s_6), .O(gate10inter1));
  and2  gate247(.a(N77), .b(N73), .O(gate10inter2));
  inv1  gate248(.a(s_6), .O(gate10inter3));
  inv1  gate249(.a(s_7), .O(gate10inter4));
  nand2 gate250(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate251(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate252(.a(N73), .O(gate10inter7));
  inv1  gate253(.a(N77), .O(gate10inter8));
  nand2 gate254(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate255(.a(s_7), .b(gate10inter3), .O(gate10inter10));
  nor2  gate256(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate257(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate258(.a(gate10inter12), .b(gate10inter1), .O(N259));
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );

  xor2  gate287(.a(N109), .b(N105), .O(gate14inter0));
  nand2 gate288(.a(gate14inter0), .b(s_12), .O(gate14inter1));
  and2  gate289(.a(N109), .b(N105), .O(gate14inter2));
  inv1  gate290(.a(s_12), .O(gate14inter3));
  inv1  gate291(.a(s_13), .O(gate14inter4));
  nand2 gate292(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate293(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate294(.a(N105), .O(gate14inter7));
  inv1  gate295(.a(N109), .O(gate14inter8));
  nand2 gate296(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate297(.a(s_13), .b(gate14inter3), .O(gate14inter10));
  nor2  gate298(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate299(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate300(.a(gate14inter12), .b(gate14inter1), .O(N263));

  xor2  gate483(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate484(.a(gate15inter0), .b(s_40), .O(gate15inter1));
  and2  gate485(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate486(.a(s_40), .O(gate15inter3));
  inv1  gate487(.a(s_41), .O(gate15inter4));
  nand2 gate488(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate489(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate490(.a(N113), .O(gate15inter7));
  inv1  gate491(.a(N117), .O(gate15inter8));
  nand2 gate492(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate493(.a(s_41), .b(gate15inter3), .O(gate15inter10));
  nor2  gate494(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate495(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate496(.a(gate15inter12), .b(gate15inter1), .O(N264));

  xor2  gate469(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate470(.a(gate16inter0), .b(s_38), .O(gate16inter1));
  and2  gate471(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate472(.a(s_38), .O(gate16inter3));
  inv1  gate473(.a(s_39), .O(gate16inter4));
  nand2 gate474(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate475(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate476(.a(N121), .O(gate16inter7));
  inv1  gate477(.a(N125), .O(gate16inter8));
  nand2 gate478(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate479(.a(s_39), .b(gate16inter3), .O(gate16inter10));
  nor2  gate480(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate481(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate482(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate259(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate260(.a(gate30inter0), .b(s_8), .O(gate30inter1));
  and2  gate261(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate262(.a(s_8), .O(gate30inter3));
  inv1  gate263(.a(s_9), .O(gate30inter4));
  nand2 gate264(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate265(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate266(.a(N41), .O(gate30inter7));
  inv1  gate267(.a(N57), .O(gate30inter8));
  nand2 gate268(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate269(.a(s_9), .b(gate30inter3), .O(gate30inter10));
  nor2  gate270(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate271(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate272(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );

  xor2  gate497(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate498(.a(gate32inter0), .b(s_42), .O(gate32inter1));
  and2  gate499(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate500(.a(s_42), .O(gate32inter3));
  inv1  gate501(.a(s_43), .O(gate32inter4));
  nand2 gate502(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate503(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate504(.a(N45), .O(gate32inter7));
  inv1  gate505(.a(N61), .O(gate32inter8));
  nand2 gate506(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate507(.a(s_43), .b(gate32inter3), .O(gate32inter10));
  nor2  gate508(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate509(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate510(.a(gate32inter12), .b(gate32inter1), .O(N281));
xor2 gate33( .a(N65), .b(N81), .O(N282) );

  xor2  gate273(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate274(.a(gate34inter0), .b(s_10), .O(gate34inter1));
  and2  gate275(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate276(.a(s_10), .O(gate34inter3));
  inv1  gate277(.a(s_11), .O(gate34inter4));
  nand2 gate278(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate279(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate280(.a(N97), .O(gate34inter7));
  inv1  gate281(.a(N113), .O(gate34inter8));
  nand2 gate282(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate283(.a(s_11), .b(gate34inter3), .O(gate34inter10));
  nor2  gate284(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate285(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate286(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate511(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate512(.a(gate42inter0), .b(s_44), .O(gate42inter1));
  and2  gate513(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate514(.a(s_44), .O(gate42inter3));
  inv1  gate515(.a(s_45), .O(gate42inter4));
  nand2 gate516(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate517(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate518(.a(N252), .O(gate42inter7));
  inv1  gate519(.a(N253), .O(gate42inter8));
  nand2 gate520(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate521(.a(s_45), .b(gate42inter3), .O(gate42inter10));
  nor2  gate522(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate523(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate524(.a(gate42inter12), .b(gate42inter1), .O(N293));
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );

  xor2  gate455(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate456(.a(gate48inter0), .b(s_36), .O(gate48inter1));
  and2  gate457(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate458(.a(s_36), .O(gate48inter3));
  inv1  gate459(.a(s_37), .O(gate48inter4));
  nand2 gate460(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate461(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate462(.a(N264), .O(gate48inter7));
  inv1  gate463(.a(N265), .O(gate48inter8));
  nand2 gate464(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate465(.a(s_37), .b(gate48inter3), .O(gate48inter10));
  nor2  gate466(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate467(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate468(.a(gate48inter12), .b(gate48inter1), .O(N311));
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate217(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate218(.a(gate50inter0), .b(s_2), .O(gate50inter1));
  and2  gate219(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate220(.a(s_2), .O(gate50inter3));
  inv1  gate221(.a(s_3), .O(gate50inter4));
  nand2 gate222(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate223(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate224(.a(N276), .O(gate50inter7));
  inv1  gate225(.a(N277), .O(gate50inter8));
  nand2 gate226(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate227(.a(s_3), .b(gate50inter3), .O(gate50inter10));
  nor2  gate228(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate229(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate230(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate315(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate316(.a(gate55inter0), .b(s_16), .O(gate55inter1));
  and2  gate317(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate318(.a(s_16), .O(gate55inter3));
  inv1  gate319(.a(s_17), .O(gate55inter4));
  nand2 gate320(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate321(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate322(.a(N286), .O(gate55inter7));
  inv1  gate323(.a(N287), .O(gate55inter8));
  nand2 gate324(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate325(.a(s_17), .b(gate55inter3), .O(gate55inter10));
  nor2  gate326(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate327(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate328(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );

  xor2  gate371(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate372(.a(gate57inter0), .b(s_24), .O(gate57inter1));
  and2  gate373(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate374(.a(s_24), .O(gate57inter3));
  inv1  gate375(.a(s_25), .O(gate57inter4));
  nand2 gate376(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate377(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate378(.a(N290), .O(gate57inter7));
  inv1  gate379(.a(N293), .O(gate57inter8));
  nand2 gate380(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate381(.a(s_25), .b(gate57inter3), .O(gate57inter10));
  nor2  gate382(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate383(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate384(.a(gate57inter12), .b(gate57inter1), .O(N338));
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate441(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate442(.a(gate59inter0), .b(s_34), .O(gate59inter1));
  and2  gate443(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate444(.a(s_34), .O(gate59inter3));
  inv1  gate445(.a(s_35), .O(gate59inter4));
  nand2 gate446(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate447(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate448(.a(N290), .O(gate59inter7));
  inv1  gate449(.a(N296), .O(gate59inter8));
  nand2 gate450(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate451(.a(s_35), .b(gate59inter3), .O(gate59inter10));
  nor2  gate452(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate453(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate454(.a(gate59inter12), .b(gate59inter1), .O(N340));

  xor2  gate413(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate414(.a(gate60inter0), .b(s_30), .O(gate60inter1));
  and2  gate415(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate416(.a(s_30), .O(gate60inter3));
  inv1  gate417(.a(s_31), .O(gate60inter4));
  nand2 gate418(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate419(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate420(.a(N293), .O(gate60inter7));
  inv1  gate421(.a(N299), .O(gate60inter8));
  nand2 gate422(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate423(.a(s_31), .b(gate60inter3), .O(gate60inter10));
  nor2  gate424(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate425(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate426(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );

  xor2  gate385(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate386(.a(gate73inter0), .b(s_26), .O(gate73inter1));
  and2  gate387(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate388(.a(s_26), .O(gate73inter3));
  inv1  gate389(.a(s_27), .O(gate73inter4));
  nand2 gate390(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate391(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate392(.a(N314), .O(gate73inter7));
  inv1  gate393(.a(N346), .O(gate73inter8));
  nand2 gate394(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate395(.a(s_27), .b(gate73inter3), .O(gate73inter10));
  nor2  gate396(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate397(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate398(.a(gate73inter12), .b(gate73inter1), .O(N354));

  xor2  gate203(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate204(.a(gate74inter0), .b(s_0), .O(gate74inter1));
  and2  gate205(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate206(.a(s_0), .O(gate74inter3));
  inv1  gate207(.a(s_1), .O(gate74inter4));
  nand2 gate208(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate209(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate210(.a(N315), .O(gate74inter7));
  inv1  gate211(.a(N347), .O(gate74inter8));
  nand2 gate212(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate213(.a(s_1), .b(gate74inter3), .O(gate74inter10));
  nor2  gate214(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate215(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate216(.a(gate74inter12), .b(gate74inter1), .O(N367));

  xor2  gate231(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate232(.a(gate75inter0), .b(s_4), .O(gate75inter1));
  and2  gate233(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate234(.a(s_4), .O(gate75inter3));
  inv1  gate235(.a(s_5), .O(gate75inter4));
  nand2 gate236(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate237(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate238(.a(N316), .O(gate75inter7));
  inv1  gate239(.a(N348), .O(gate75inter8));
  nand2 gate240(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate241(.a(s_5), .b(gate75inter3), .O(gate75inter10));
  nor2  gate242(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate243(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate244(.a(gate75inter12), .b(gate75inter1), .O(N380));

  xor2  gate329(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate330(.a(gate76inter0), .b(s_18), .O(gate76inter1));
  and2  gate331(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate332(.a(s_18), .O(gate76inter3));
  inv1  gate333(.a(s_19), .O(gate76inter4));
  nand2 gate334(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate335(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate336(.a(N317), .O(gate76inter7));
  inv1  gate337(.a(N349), .O(gate76inter8));
  nand2 gate338(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate339(.a(s_19), .b(gate76inter3), .O(gate76inter10));
  nor2  gate340(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate341(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate342(.a(gate76inter12), .b(gate76inter1), .O(N393));
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );

  xor2  gate525(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate526(.a(gate173inter0), .b(s_46), .O(gate173inter1));
  and2  gate527(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate528(.a(s_46), .O(gate173inter3));
  inv1  gate529(.a(s_47), .O(gate173inter4));
  nand2 gate530(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate531(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate532(.a(N9), .O(gate173inter7));
  inv1  gate533(.a(N694), .O(gate173inter8));
  nand2 gate534(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate535(.a(s_47), .b(gate173inter3), .O(gate173inter10));
  nor2  gate536(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate537(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate538(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );

  xor2  gate553(.a(N696), .b(N17), .O(gate175inter0));
  nand2 gate554(.a(gate175inter0), .b(s_50), .O(gate175inter1));
  and2  gate555(.a(N696), .b(N17), .O(gate175inter2));
  inv1  gate556(.a(s_50), .O(gate175inter3));
  inv1  gate557(.a(s_51), .O(gate175inter4));
  nand2 gate558(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate559(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate560(.a(N17), .O(gate175inter7));
  inv1  gate561(.a(N696), .O(gate175inter8));
  nand2 gate562(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate563(.a(s_51), .b(gate175inter3), .O(gate175inter10));
  nor2  gate564(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate565(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate566(.a(gate175inter12), .b(gate175inter1), .O(N728));
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );
xor2 gate183( .a(N49), .b(N704), .O(N736) );

  xor2  gate343(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate344(.a(gate184inter0), .b(s_20), .O(gate184inter1));
  and2  gate345(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate346(.a(s_20), .O(gate184inter3));
  inv1  gate347(.a(s_21), .O(gate184inter4));
  nand2 gate348(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate349(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate350(.a(N53), .O(gate184inter7));
  inv1  gate351(.a(N705), .O(gate184inter8));
  nand2 gate352(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate353(.a(s_21), .b(gate184inter3), .O(gate184inter10));
  nor2  gate354(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate355(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate356(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate399(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate400(.a(gate186inter0), .b(s_28), .O(gate186inter1));
  and2  gate401(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate402(.a(s_28), .O(gate186inter3));
  inv1  gate403(.a(s_29), .O(gate186inter4));
  nand2 gate404(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate405(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate406(.a(N61), .O(gate186inter7));
  inv1  gate407(.a(N707), .O(gate186inter8));
  nand2 gate408(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate409(.a(s_29), .b(gate186inter3), .O(gate186inter10));
  nor2  gate410(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate411(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate412(.a(gate186inter12), .b(gate186inter1), .O(N739));
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );

  xor2  gate427(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate428(.a(gate199inter0), .b(s_32), .O(gate199inter1));
  and2  gate429(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate430(.a(s_32), .O(gate199inter3));
  inv1  gate431(.a(s_33), .O(gate199inter4));
  nand2 gate432(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate433(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate434(.a(N113), .O(gate199inter7));
  inv1  gate435(.a(N720), .O(gate199inter8));
  nand2 gate436(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate437(.a(s_33), .b(gate199inter3), .O(gate199inter10));
  nor2  gate438(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate439(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate440(.a(gate199inter12), .b(gate199inter1), .O(N752));

  xor2  gate357(.a(N721), .b(N117), .O(gate200inter0));
  nand2 gate358(.a(gate200inter0), .b(s_22), .O(gate200inter1));
  and2  gate359(.a(N721), .b(N117), .O(gate200inter2));
  inv1  gate360(.a(s_22), .O(gate200inter3));
  inv1  gate361(.a(s_23), .O(gate200inter4));
  nand2 gate362(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate363(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate364(.a(N117), .O(gate200inter7));
  inv1  gate365(.a(N721), .O(gate200inter8));
  nand2 gate366(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate367(.a(s_23), .b(gate200inter3), .O(gate200inter10));
  nor2  gate368(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate369(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate370(.a(gate200inter12), .b(gate200inter1), .O(N753));
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule