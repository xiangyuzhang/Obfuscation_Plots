module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1947(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1948(.a(gate12inter0), .b(s_200), .O(gate12inter1));
  and2  gate1949(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1950(.a(s_200), .O(gate12inter3));
  inv1  gate1951(.a(s_201), .O(gate12inter4));
  nand2 gate1952(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1953(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1954(.a(G7), .O(gate12inter7));
  inv1  gate1955(.a(G8), .O(gate12inter8));
  nand2 gate1956(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1957(.a(s_201), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1958(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1959(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1960(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate659(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate660(.a(gate14inter0), .b(s_16), .O(gate14inter1));
  and2  gate661(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate662(.a(s_16), .O(gate14inter3));
  inv1  gate663(.a(s_17), .O(gate14inter4));
  nand2 gate664(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate665(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate666(.a(G11), .O(gate14inter7));
  inv1  gate667(.a(G12), .O(gate14inter8));
  nand2 gate668(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate669(.a(s_17), .b(gate14inter3), .O(gate14inter10));
  nor2  gate670(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate671(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate672(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate981(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate982(.a(gate16inter0), .b(s_62), .O(gate16inter1));
  and2  gate983(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate984(.a(s_62), .O(gate16inter3));
  inv1  gate985(.a(s_63), .O(gate16inter4));
  nand2 gate986(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate987(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate988(.a(G15), .O(gate16inter7));
  inv1  gate989(.a(G16), .O(gate16inter8));
  nand2 gate990(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate991(.a(s_63), .b(gate16inter3), .O(gate16inter10));
  nor2  gate992(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate993(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate994(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate687(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate688(.a(gate21inter0), .b(s_20), .O(gate21inter1));
  and2  gate689(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate690(.a(s_20), .O(gate21inter3));
  inv1  gate691(.a(s_21), .O(gate21inter4));
  nand2 gate692(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate693(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate694(.a(G25), .O(gate21inter7));
  inv1  gate695(.a(G26), .O(gate21inter8));
  nand2 gate696(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate697(.a(s_21), .b(gate21inter3), .O(gate21inter10));
  nor2  gate698(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate699(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate700(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1261(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1262(.a(gate31inter0), .b(s_102), .O(gate31inter1));
  and2  gate1263(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1264(.a(s_102), .O(gate31inter3));
  inv1  gate1265(.a(s_103), .O(gate31inter4));
  nand2 gate1266(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1267(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1268(.a(G4), .O(gate31inter7));
  inv1  gate1269(.a(G8), .O(gate31inter8));
  nand2 gate1270(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1271(.a(s_103), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1272(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1273(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1274(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2017(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2018(.a(gate33inter0), .b(s_210), .O(gate33inter1));
  and2  gate2019(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2020(.a(s_210), .O(gate33inter3));
  inv1  gate2021(.a(s_211), .O(gate33inter4));
  nand2 gate2022(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2023(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2024(.a(G17), .O(gate33inter7));
  inv1  gate2025(.a(G21), .O(gate33inter8));
  nand2 gate2026(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2027(.a(s_211), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2028(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2029(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2030(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1905(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1906(.a(gate35inter0), .b(s_194), .O(gate35inter1));
  and2  gate1907(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1908(.a(s_194), .O(gate35inter3));
  inv1  gate1909(.a(s_195), .O(gate35inter4));
  nand2 gate1910(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1911(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1912(.a(G18), .O(gate35inter7));
  inv1  gate1913(.a(G22), .O(gate35inter8));
  nand2 gate1914(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1915(.a(s_195), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1916(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1917(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1918(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate1191(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1192(.a(gate36inter0), .b(s_92), .O(gate36inter1));
  and2  gate1193(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1194(.a(s_92), .O(gate36inter3));
  inv1  gate1195(.a(s_93), .O(gate36inter4));
  nand2 gate1196(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1197(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1198(.a(G26), .O(gate36inter7));
  inv1  gate1199(.a(G30), .O(gate36inter8));
  nand2 gate1200(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1201(.a(s_93), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1202(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1203(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1204(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate869(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate870(.a(gate39inter0), .b(s_46), .O(gate39inter1));
  and2  gate871(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate872(.a(s_46), .O(gate39inter3));
  inv1  gate873(.a(s_47), .O(gate39inter4));
  nand2 gate874(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate875(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate876(.a(G20), .O(gate39inter7));
  inv1  gate877(.a(G24), .O(gate39inter8));
  nand2 gate878(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate879(.a(s_47), .b(gate39inter3), .O(gate39inter10));
  nor2  gate880(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate881(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate882(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1233(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1234(.a(gate40inter0), .b(s_98), .O(gate40inter1));
  and2  gate1235(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1236(.a(s_98), .O(gate40inter3));
  inv1  gate1237(.a(s_99), .O(gate40inter4));
  nand2 gate1238(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1239(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1240(.a(G28), .O(gate40inter7));
  inv1  gate1241(.a(G32), .O(gate40inter8));
  nand2 gate1242(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1243(.a(s_99), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1244(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1245(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1246(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1975(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1976(.a(gate41inter0), .b(s_204), .O(gate41inter1));
  and2  gate1977(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1978(.a(s_204), .O(gate41inter3));
  inv1  gate1979(.a(s_205), .O(gate41inter4));
  nand2 gate1980(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1981(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1982(.a(G1), .O(gate41inter7));
  inv1  gate1983(.a(G266), .O(gate41inter8));
  nand2 gate1984(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1985(.a(s_205), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1986(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1987(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1988(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1625(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1626(.a(gate43inter0), .b(s_154), .O(gate43inter1));
  and2  gate1627(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1628(.a(s_154), .O(gate43inter3));
  inv1  gate1629(.a(s_155), .O(gate43inter4));
  nand2 gate1630(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1631(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1632(.a(G3), .O(gate43inter7));
  inv1  gate1633(.a(G269), .O(gate43inter8));
  nand2 gate1634(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1635(.a(s_155), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1636(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1637(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1638(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1891(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1892(.a(gate45inter0), .b(s_192), .O(gate45inter1));
  and2  gate1893(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1894(.a(s_192), .O(gate45inter3));
  inv1  gate1895(.a(s_193), .O(gate45inter4));
  nand2 gate1896(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1897(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1898(.a(G5), .O(gate45inter7));
  inv1  gate1899(.a(G272), .O(gate45inter8));
  nand2 gate1900(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1901(.a(s_193), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1902(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1903(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1904(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1345(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1346(.a(gate47inter0), .b(s_114), .O(gate47inter1));
  and2  gate1347(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1348(.a(s_114), .O(gate47inter3));
  inv1  gate1349(.a(s_115), .O(gate47inter4));
  nand2 gate1350(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1351(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1352(.a(G7), .O(gate47inter7));
  inv1  gate1353(.a(G275), .O(gate47inter8));
  nand2 gate1354(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1355(.a(s_115), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1356(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1357(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1358(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1863(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1864(.a(gate48inter0), .b(s_188), .O(gate48inter1));
  and2  gate1865(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1866(.a(s_188), .O(gate48inter3));
  inv1  gate1867(.a(s_189), .O(gate48inter4));
  nand2 gate1868(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1869(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1870(.a(G8), .O(gate48inter7));
  inv1  gate1871(.a(G275), .O(gate48inter8));
  nand2 gate1872(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1873(.a(s_189), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1874(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1875(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1876(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1639(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1640(.a(gate49inter0), .b(s_156), .O(gate49inter1));
  and2  gate1641(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1642(.a(s_156), .O(gate49inter3));
  inv1  gate1643(.a(s_157), .O(gate49inter4));
  nand2 gate1644(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1645(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1646(.a(G9), .O(gate49inter7));
  inv1  gate1647(.a(G278), .O(gate49inter8));
  nand2 gate1648(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1649(.a(s_157), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1650(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1651(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1652(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1037(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1038(.a(gate63inter0), .b(s_70), .O(gate63inter1));
  and2  gate1039(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1040(.a(s_70), .O(gate63inter3));
  inv1  gate1041(.a(s_71), .O(gate63inter4));
  nand2 gate1042(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1043(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1044(.a(G23), .O(gate63inter7));
  inv1  gate1045(.a(G299), .O(gate63inter8));
  nand2 gate1046(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1047(.a(s_71), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1048(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1049(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1050(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1009(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1010(.a(gate65inter0), .b(s_66), .O(gate65inter1));
  and2  gate1011(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1012(.a(s_66), .O(gate65inter3));
  inv1  gate1013(.a(s_67), .O(gate65inter4));
  nand2 gate1014(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1015(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1016(.a(G25), .O(gate65inter7));
  inv1  gate1017(.a(G302), .O(gate65inter8));
  nand2 gate1018(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1019(.a(s_67), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1020(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1021(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1022(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1709(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1710(.a(gate68inter0), .b(s_166), .O(gate68inter1));
  and2  gate1711(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1712(.a(s_166), .O(gate68inter3));
  inv1  gate1713(.a(s_167), .O(gate68inter4));
  nand2 gate1714(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1715(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1716(.a(G28), .O(gate68inter7));
  inv1  gate1717(.a(G305), .O(gate68inter8));
  nand2 gate1718(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1719(.a(s_167), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1720(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1721(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1722(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1513(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1514(.a(gate77inter0), .b(s_138), .O(gate77inter1));
  and2  gate1515(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1516(.a(s_138), .O(gate77inter3));
  inv1  gate1517(.a(s_139), .O(gate77inter4));
  nand2 gate1518(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1519(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1520(.a(G2), .O(gate77inter7));
  inv1  gate1521(.a(G320), .O(gate77inter8));
  nand2 gate1522(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1523(.a(s_139), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1524(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1525(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1526(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1737(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1738(.a(gate81inter0), .b(s_170), .O(gate81inter1));
  and2  gate1739(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1740(.a(s_170), .O(gate81inter3));
  inv1  gate1741(.a(s_171), .O(gate81inter4));
  nand2 gate1742(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1743(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1744(.a(G3), .O(gate81inter7));
  inv1  gate1745(.a(G326), .O(gate81inter8));
  nand2 gate1746(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1747(.a(s_171), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1748(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1749(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1750(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1373(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1374(.a(gate85inter0), .b(s_118), .O(gate85inter1));
  and2  gate1375(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1376(.a(s_118), .O(gate85inter3));
  inv1  gate1377(.a(s_119), .O(gate85inter4));
  nand2 gate1378(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1379(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1380(.a(G4), .O(gate85inter7));
  inv1  gate1381(.a(G332), .O(gate85inter8));
  nand2 gate1382(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1383(.a(s_119), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1384(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1385(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1386(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1023(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1024(.a(gate87inter0), .b(s_68), .O(gate87inter1));
  and2  gate1025(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1026(.a(s_68), .O(gate87inter3));
  inv1  gate1027(.a(s_69), .O(gate87inter4));
  nand2 gate1028(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1029(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1030(.a(G12), .O(gate87inter7));
  inv1  gate1031(.a(G335), .O(gate87inter8));
  nand2 gate1032(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1033(.a(s_69), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1034(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1035(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1036(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate785(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate786(.a(gate90inter0), .b(s_34), .O(gate90inter1));
  and2  gate787(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate788(.a(s_34), .O(gate90inter3));
  inv1  gate789(.a(s_35), .O(gate90inter4));
  nand2 gate790(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate791(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate792(.a(G21), .O(gate90inter7));
  inv1  gate793(.a(G338), .O(gate90inter8));
  nand2 gate794(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate795(.a(s_35), .b(gate90inter3), .O(gate90inter10));
  nor2  gate796(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate797(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate798(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate589(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate590(.a(gate95inter0), .b(s_6), .O(gate95inter1));
  and2  gate591(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate592(.a(s_6), .O(gate95inter3));
  inv1  gate593(.a(s_7), .O(gate95inter4));
  nand2 gate594(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate595(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate596(.a(G26), .O(gate95inter7));
  inv1  gate597(.a(G347), .O(gate95inter8));
  nand2 gate598(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate599(.a(s_7), .b(gate95inter3), .O(gate95inter10));
  nor2  gate600(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate601(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate602(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1849(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1850(.a(gate98inter0), .b(s_186), .O(gate98inter1));
  and2  gate1851(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1852(.a(s_186), .O(gate98inter3));
  inv1  gate1853(.a(s_187), .O(gate98inter4));
  nand2 gate1854(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1855(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1856(.a(G23), .O(gate98inter7));
  inv1  gate1857(.a(G350), .O(gate98inter8));
  nand2 gate1858(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1859(.a(s_187), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1860(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1861(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1862(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate883(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate884(.a(gate103inter0), .b(s_48), .O(gate103inter1));
  and2  gate885(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate886(.a(s_48), .O(gate103inter3));
  inv1  gate887(.a(s_49), .O(gate103inter4));
  nand2 gate888(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate889(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate890(.a(G28), .O(gate103inter7));
  inv1  gate891(.a(G359), .O(gate103inter8));
  nand2 gate892(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate893(.a(s_49), .b(gate103inter3), .O(gate103inter10));
  nor2  gate894(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate895(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate896(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1583(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1584(.a(gate106inter0), .b(s_148), .O(gate106inter1));
  and2  gate1585(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1586(.a(s_148), .O(gate106inter3));
  inv1  gate1587(.a(s_149), .O(gate106inter4));
  nand2 gate1588(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1589(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1590(.a(G364), .O(gate106inter7));
  inv1  gate1591(.a(G365), .O(gate106inter8));
  nand2 gate1592(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1593(.a(s_149), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1594(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1595(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1596(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1079(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1080(.a(gate115inter0), .b(s_76), .O(gate115inter1));
  and2  gate1081(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1082(.a(s_76), .O(gate115inter3));
  inv1  gate1083(.a(s_77), .O(gate115inter4));
  nand2 gate1084(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1085(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1086(.a(G382), .O(gate115inter7));
  inv1  gate1087(.a(G383), .O(gate115inter8));
  nand2 gate1088(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1089(.a(s_77), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1090(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1091(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1092(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate1051(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate1052(.a(gate118inter0), .b(s_72), .O(gate118inter1));
  and2  gate1053(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate1054(.a(s_72), .O(gate118inter3));
  inv1  gate1055(.a(s_73), .O(gate118inter4));
  nand2 gate1056(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1057(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1058(.a(G388), .O(gate118inter7));
  inv1  gate1059(.a(G389), .O(gate118inter8));
  nand2 gate1060(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1061(.a(s_73), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1062(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1063(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1064(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1205(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1206(.a(gate119inter0), .b(s_94), .O(gate119inter1));
  and2  gate1207(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1208(.a(s_94), .O(gate119inter3));
  inv1  gate1209(.a(s_95), .O(gate119inter4));
  nand2 gate1210(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1211(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1212(.a(G390), .O(gate119inter7));
  inv1  gate1213(.a(G391), .O(gate119inter8));
  nand2 gate1214(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1215(.a(s_95), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1216(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1217(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1218(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2045(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2046(.a(gate124inter0), .b(s_214), .O(gate124inter1));
  and2  gate2047(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2048(.a(s_214), .O(gate124inter3));
  inv1  gate2049(.a(s_215), .O(gate124inter4));
  nand2 gate2050(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2051(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2052(.a(G400), .O(gate124inter7));
  inv1  gate2053(.a(G401), .O(gate124inter8));
  nand2 gate2054(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2055(.a(s_215), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2056(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2057(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2058(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1457(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1458(.a(gate140inter0), .b(s_130), .O(gate140inter1));
  and2  gate1459(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1460(.a(s_130), .O(gate140inter3));
  inv1  gate1461(.a(s_131), .O(gate140inter4));
  nand2 gate1462(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1463(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1464(.a(G444), .O(gate140inter7));
  inv1  gate1465(.a(G447), .O(gate140inter8));
  nand2 gate1466(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1467(.a(s_131), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1468(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1469(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1470(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate561(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate562(.a(gate141inter0), .b(s_2), .O(gate141inter1));
  and2  gate563(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate564(.a(s_2), .O(gate141inter3));
  inv1  gate565(.a(s_3), .O(gate141inter4));
  nand2 gate566(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate567(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate568(.a(G450), .O(gate141inter7));
  inv1  gate569(.a(G453), .O(gate141inter8));
  nand2 gate570(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate571(.a(s_3), .b(gate141inter3), .O(gate141inter10));
  nor2  gate572(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate573(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate574(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate547(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate548(.a(gate145inter0), .b(s_0), .O(gate145inter1));
  and2  gate549(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate550(.a(s_0), .O(gate145inter3));
  inv1  gate551(.a(s_1), .O(gate145inter4));
  nand2 gate552(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate553(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate554(.a(G474), .O(gate145inter7));
  inv1  gate555(.a(G477), .O(gate145inter8));
  nand2 gate556(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate557(.a(s_1), .b(gate145inter3), .O(gate145inter10));
  nor2  gate558(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate559(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate560(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate2087(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2088(.a(gate149inter0), .b(s_220), .O(gate149inter1));
  and2  gate2089(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2090(.a(s_220), .O(gate149inter3));
  inv1  gate2091(.a(s_221), .O(gate149inter4));
  nand2 gate2092(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2093(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2094(.a(G498), .O(gate149inter7));
  inv1  gate2095(.a(G501), .O(gate149inter8));
  nand2 gate2096(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2097(.a(s_221), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2098(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2099(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2100(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate953(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate954(.a(gate154inter0), .b(s_58), .O(gate154inter1));
  and2  gate955(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate956(.a(s_58), .O(gate154inter3));
  inv1  gate957(.a(s_59), .O(gate154inter4));
  nand2 gate958(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate959(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate960(.a(G429), .O(gate154inter7));
  inv1  gate961(.a(G522), .O(gate154inter8));
  nand2 gate962(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate963(.a(s_59), .b(gate154inter3), .O(gate154inter10));
  nor2  gate964(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate965(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate966(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate911(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate912(.a(gate159inter0), .b(s_52), .O(gate159inter1));
  and2  gate913(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate914(.a(s_52), .O(gate159inter3));
  inv1  gate915(.a(s_53), .O(gate159inter4));
  nand2 gate916(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate917(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate918(.a(G444), .O(gate159inter7));
  inv1  gate919(.a(G531), .O(gate159inter8));
  nand2 gate920(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate921(.a(s_53), .b(gate159inter3), .O(gate159inter10));
  nor2  gate922(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate923(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate924(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1303(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1304(.a(gate161inter0), .b(s_108), .O(gate161inter1));
  and2  gate1305(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1306(.a(s_108), .O(gate161inter3));
  inv1  gate1307(.a(s_109), .O(gate161inter4));
  nand2 gate1308(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1309(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1310(.a(G450), .O(gate161inter7));
  inv1  gate1311(.a(G534), .O(gate161inter8));
  nand2 gate1312(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1313(.a(s_109), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1314(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1315(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1316(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1275(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1276(.a(gate163inter0), .b(s_104), .O(gate163inter1));
  and2  gate1277(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1278(.a(s_104), .O(gate163inter3));
  inv1  gate1279(.a(s_105), .O(gate163inter4));
  nand2 gate1280(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1281(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1282(.a(G456), .O(gate163inter7));
  inv1  gate1283(.a(G537), .O(gate163inter8));
  nand2 gate1284(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1285(.a(s_105), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1286(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1287(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1288(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate995(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate996(.a(gate164inter0), .b(s_64), .O(gate164inter1));
  and2  gate997(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate998(.a(s_64), .O(gate164inter3));
  inv1  gate999(.a(s_65), .O(gate164inter4));
  nand2 gate1000(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1001(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1002(.a(G459), .O(gate164inter7));
  inv1  gate1003(.a(G537), .O(gate164inter8));
  nand2 gate1004(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1005(.a(s_65), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1006(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1007(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1008(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1317(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1318(.a(gate168inter0), .b(s_110), .O(gate168inter1));
  and2  gate1319(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1320(.a(s_110), .O(gate168inter3));
  inv1  gate1321(.a(s_111), .O(gate168inter4));
  nand2 gate1322(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1323(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1324(.a(G471), .O(gate168inter7));
  inv1  gate1325(.a(G543), .O(gate168inter8));
  nand2 gate1326(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1327(.a(s_111), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1328(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1329(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1330(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2059(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2060(.a(gate173inter0), .b(s_216), .O(gate173inter1));
  and2  gate2061(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2062(.a(s_216), .O(gate173inter3));
  inv1  gate2063(.a(s_217), .O(gate173inter4));
  nand2 gate2064(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2065(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2066(.a(G486), .O(gate173inter7));
  inv1  gate2067(.a(G552), .O(gate173inter8));
  nand2 gate2068(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2069(.a(s_217), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2070(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2071(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2072(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1793(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1794(.a(gate174inter0), .b(s_178), .O(gate174inter1));
  and2  gate1795(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1796(.a(s_178), .O(gate174inter3));
  inv1  gate1797(.a(s_179), .O(gate174inter4));
  nand2 gate1798(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1799(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1800(.a(G489), .O(gate174inter7));
  inv1  gate1801(.a(G552), .O(gate174inter8));
  nand2 gate1802(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1803(.a(s_179), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1804(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1805(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1806(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1555(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1556(.a(gate176inter0), .b(s_144), .O(gate176inter1));
  and2  gate1557(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1558(.a(s_144), .O(gate176inter3));
  inv1  gate1559(.a(s_145), .O(gate176inter4));
  nand2 gate1560(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1561(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1562(.a(G495), .O(gate176inter7));
  inv1  gate1563(.a(G555), .O(gate176inter8));
  nand2 gate1564(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1565(.a(s_145), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1566(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1567(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1568(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1541(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1542(.a(gate178inter0), .b(s_142), .O(gate178inter1));
  and2  gate1543(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1544(.a(s_142), .O(gate178inter3));
  inv1  gate1545(.a(s_143), .O(gate178inter4));
  nand2 gate1546(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1547(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1548(.a(G501), .O(gate178inter7));
  inv1  gate1549(.a(G558), .O(gate178inter8));
  nand2 gate1550(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1551(.a(s_143), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1552(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1553(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1554(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1989(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1990(.a(gate182inter0), .b(s_206), .O(gate182inter1));
  and2  gate1991(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1992(.a(s_206), .O(gate182inter3));
  inv1  gate1993(.a(s_207), .O(gate182inter4));
  nand2 gate1994(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1995(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1996(.a(G513), .O(gate182inter7));
  inv1  gate1997(.a(G564), .O(gate182inter8));
  nand2 gate1998(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1999(.a(s_207), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2000(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2001(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2002(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate897(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate898(.a(gate187inter0), .b(s_50), .O(gate187inter1));
  and2  gate899(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate900(.a(s_50), .O(gate187inter3));
  inv1  gate901(.a(s_51), .O(gate187inter4));
  nand2 gate902(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate903(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate904(.a(G574), .O(gate187inter7));
  inv1  gate905(.a(G575), .O(gate187inter8));
  nand2 gate906(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate907(.a(s_51), .b(gate187inter3), .O(gate187inter10));
  nor2  gate908(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate909(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate910(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1765(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1766(.a(gate189inter0), .b(s_174), .O(gate189inter1));
  and2  gate1767(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1768(.a(s_174), .O(gate189inter3));
  inv1  gate1769(.a(s_175), .O(gate189inter4));
  nand2 gate1770(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1771(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1772(.a(G578), .O(gate189inter7));
  inv1  gate1773(.a(G579), .O(gate189inter8));
  nand2 gate1774(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1775(.a(s_175), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1776(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1777(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1778(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1835(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1836(.a(gate191inter0), .b(s_184), .O(gate191inter1));
  and2  gate1837(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1838(.a(s_184), .O(gate191inter3));
  inv1  gate1839(.a(s_185), .O(gate191inter4));
  nand2 gate1840(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1841(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1842(.a(G582), .O(gate191inter7));
  inv1  gate1843(.a(G583), .O(gate191inter8));
  nand2 gate1844(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1845(.a(s_185), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1846(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1847(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1848(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1499(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1500(.a(gate196inter0), .b(s_136), .O(gate196inter1));
  and2  gate1501(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1502(.a(s_136), .O(gate196inter3));
  inv1  gate1503(.a(s_137), .O(gate196inter4));
  nand2 gate1504(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1505(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1506(.a(G592), .O(gate196inter7));
  inv1  gate1507(.a(G593), .O(gate196inter8));
  nand2 gate1508(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1509(.a(s_137), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1510(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1511(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1512(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1471(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1472(.a(gate202inter0), .b(s_132), .O(gate202inter1));
  and2  gate1473(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1474(.a(s_132), .O(gate202inter3));
  inv1  gate1475(.a(s_133), .O(gate202inter4));
  nand2 gate1476(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1477(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1478(.a(G612), .O(gate202inter7));
  inv1  gate1479(.a(G617), .O(gate202inter8));
  nand2 gate1480(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1481(.a(s_133), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1482(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1483(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1484(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1093(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1094(.a(gate210inter0), .b(s_78), .O(gate210inter1));
  and2  gate1095(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1096(.a(s_78), .O(gate210inter3));
  inv1  gate1097(.a(s_79), .O(gate210inter4));
  nand2 gate1098(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1099(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1100(.a(G607), .O(gate210inter7));
  inv1  gate1101(.a(G666), .O(gate210inter8));
  nand2 gate1102(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1103(.a(s_79), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1104(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1105(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1106(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1779(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1780(.a(gate220inter0), .b(s_176), .O(gate220inter1));
  and2  gate1781(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1782(.a(s_176), .O(gate220inter3));
  inv1  gate1783(.a(s_177), .O(gate220inter4));
  nand2 gate1784(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1785(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1786(.a(G637), .O(gate220inter7));
  inv1  gate1787(.a(G681), .O(gate220inter8));
  nand2 gate1788(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1789(.a(s_177), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1790(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1791(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1792(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1961(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1962(.a(gate228inter0), .b(s_202), .O(gate228inter1));
  and2  gate1963(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1964(.a(s_202), .O(gate228inter3));
  inv1  gate1965(.a(s_203), .O(gate228inter4));
  nand2 gate1966(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1967(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1968(.a(G696), .O(gate228inter7));
  inv1  gate1969(.a(G697), .O(gate228inter8));
  nand2 gate1970(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1971(.a(s_203), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1972(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1973(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1974(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1723(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1724(.a(gate229inter0), .b(s_168), .O(gate229inter1));
  and2  gate1725(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1726(.a(s_168), .O(gate229inter3));
  inv1  gate1727(.a(s_169), .O(gate229inter4));
  nand2 gate1728(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1729(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1730(.a(G698), .O(gate229inter7));
  inv1  gate1731(.a(G699), .O(gate229inter8));
  nand2 gate1732(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1733(.a(s_169), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1734(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1735(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1736(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1681(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1682(.a(gate232inter0), .b(s_162), .O(gate232inter1));
  and2  gate1683(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1684(.a(s_162), .O(gate232inter3));
  inv1  gate1685(.a(s_163), .O(gate232inter4));
  nand2 gate1686(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1687(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1688(.a(G704), .O(gate232inter7));
  inv1  gate1689(.a(G705), .O(gate232inter8));
  nand2 gate1690(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1691(.a(s_163), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1692(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1693(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1694(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate939(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate940(.a(gate236inter0), .b(s_56), .O(gate236inter1));
  and2  gate941(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate942(.a(s_56), .O(gate236inter3));
  inv1  gate943(.a(s_57), .O(gate236inter4));
  nand2 gate944(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate945(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate946(.a(G251), .O(gate236inter7));
  inv1  gate947(.a(G727), .O(gate236inter8));
  nand2 gate948(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate949(.a(s_57), .b(gate236inter3), .O(gate236inter10));
  nor2  gate950(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate951(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate952(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1751(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1752(.a(gate242inter0), .b(s_172), .O(gate242inter1));
  and2  gate1753(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1754(.a(s_172), .O(gate242inter3));
  inv1  gate1755(.a(s_173), .O(gate242inter4));
  nand2 gate1756(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1757(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1758(.a(G718), .O(gate242inter7));
  inv1  gate1759(.a(G730), .O(gate242inter8));
  nand2 gate1760(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1761(.a(s_173), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1762(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1763(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1764(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate813(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate814(.a(gate244inter0), .b(s_38), .O(gate244inter1));
  and2  gate815(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate816(.a(s_38), .O(gate244inter3));
  inv1  gate817(.a(s_39), .O(gate244inter4));
  nand2 gate818(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate819(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate820(.a(G721), .O(gate244inter7));
  inv1  gate821(.a(G733), .O(gate244inter8));
  nand2 gate822(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate823(.a(s_39), .b(gate244inter3), .O(gate244inter10));
  nor2  gate824(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate825(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate826(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate827(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate828(.a(gate245inter0), .b(s_40), .O(gate245inter1));
  and2  gate829(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate830(.a(s_40), .O(gate245inter3));
  inv1  gate831(.a(s_41), .O(gate245inter4));
  nand2 gate832(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate833(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate834(.a(G248), .O(gate245inter7));
  inv1  gate835(.a(G736), .O(gate245inter8));
  nand2 gate836(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate837(.a(s_41), .b(gate245inter3), .O(gate245inter10));
  nor2  gate838(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate839(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate840(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1415(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1416(.a(gate246inter0), .b(s_124), .O(gate246inter1));
  and2  gate1417(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1418(.a(s_124), .O(gate246inter3));
  inv1  gate1419(.a(s_125), .O(gate246inter4));
  nand2 gate1420(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1421(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1422(.a(G724), .O(gate246inter7));
  inv1  gate1423(.a(G736), .O(gate246inter8));
  nand2 gate1424(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1425(.a(s_125), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1426(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1427(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1428(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate631(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate632(.a(gate248inter0), .b(s_12), .O(gate248inter1));
  and2  gate633(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate634(.a(s_12), .O(gate248inter3));
  inv1  gate635(.a(s_13), .O(gate248inter4));
  nand2 gate636(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate637(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate638(.a(G727), .O(gate248inter7));
  inv1  gate639(.a(G739), .O(gate248inter8));
  nand2 gate640(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate641(.a(s_13), .b(gate248inter3), .O(gate248inter10));
  nor2  gate642(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate643(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate644(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1695(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1696(.a(gate256inter0), .b(s_164), .O(gate256inter1));
  and2  gate1697(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1698(.a(s_164), .O(gate256inter3));
  inv1  gate1699(.a(s_165), .O(gate256inter4));
  nand2 gate1700(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1701(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1702(.a(G715), .O(gate256inter7));
  inv1  gate1703(.a(G751), .O(gate256inter8));
  nand2 gate1704(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1705(.a(s_165), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1706(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1707(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1708(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1667(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1668(.a(gate259inter0), .b(s_160), .O(gate259inter1));
  and2  gate1669(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1670(.a(s_160), .O(gate259inter3));
  inv1  gate1671(.a(s_161), .O(gate259inter4));
  nand2 gate1672(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1673(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1674(.a(G758), .O(gate259inter7));
  inv1  gate1675(.a(G759), .O(gate259inter8));
  nand2 gate1676(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1677(.a(s_161), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1678(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1679(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1680(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate799(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate800(.a(gate263inter0), .b(s_36), .O(gate263inter1));
  and2  gate801(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate802(.a(s_36), .O(gate263inter3));
  inv1  gate803(.a(s_37), .O(gate263inter4));
  nand2 gate804(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate805(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate806(.a(G766), .O(gate263inter7));
  inv1  gate807(.a(G767), .O(gate263inter8));
  nand2 gate808(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate809(.a(s_37), .b(gate263inter3), .O(gate263inter10));
  nor2  gate810(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate811(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate812(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1821(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1822(.a(gate266inter0), .b(s_182), .O(gate266inter1));
  and2  gate1823(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1824(.a(s_182), .O(gate266inter3));
  inv1  gate1825(.a(s_183), .O(gate266inter4));
  nand2 gate1826(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1827(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1828(.a(G645), .O(gate266inter7));
  inv1  gate1829(.a(G773), .O(gate266inter8));
  nand2 gate1830(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1831(.a(s_183), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1832(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1833(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1834(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate673(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate674(.a(gate271inter0), .b(s_18), .O(gate271inter1));
  and2  gate675(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate676(.a(s_18), .O(gate271inter3));
  inv1  gate677(.a(s_19), .O(gate271inter4));
  nand2 gate678(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate679(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate680(.a(G660), .O(gate271inter7));
  inv1  gate681(.a(G788), .O(gate271inter8));
  nand2 gate682(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate683(.a(s_19), .b(gate271inter3), .O(gate271inter10));
  nor2  gate684(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate685(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate686(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1401(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1402(.a(gate273inter0), .b(s_122), .O(gate273inter1));
  and2  gate1403(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1404(.a(s_122), .O(gate273inter3));
  inv1  gate1405(.a(s_123), .O(gate273inter4));
  nand2 gate1406(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1407(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1408(.a(G642), .O(gate273inter7));
  inv1  gate1409(.a(G794), .O(gate273inter8));
  nand2 gate1410(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1411(.a(s_123), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1412(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1413(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1414(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1933(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1934(.a(gate276inter0), .b(s_198), .O(gate276inter1));
  and2  gate1935(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1936(.a(s_198), .O(gate276inter3));
  inv1  gate1937(.a(s_199), .O(gate276inter4));
  nand2 gate1938(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1939(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1940(.a(G773), .O(gate276inter7));
  inv1  gate1941(.a(G797), .O(gate276inter8));
  nand2 gate1942(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1943(.a(s_199), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1944(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1945(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1946(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate771(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate772(.a(gate279inter0), .b(s_32), .O(gate279inter1));
  and2  gate773(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate774(.a(s_32), .O(gate279inter3));
  inv1  gate775(.a(s_33), .O(gate279inter4));
  nand2 gate776(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate777(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate778(.a(G651), .O(gate279inter7));
  inv1  gate779(.a(G803), .O(gate279inter8));
  nand2 gate780(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate781(.a(s_33), .b(gate279inter3), .O(gate279inter10));
  nor2  gate782(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate783(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate784(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1919(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1920(.a(gate285inter0), .b(s_196), .O(gate285inter1));
  and2  gate1921(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1922(.a(s_196), .O(gate285inter3));
  inv1  gate1923(.a(s_197), .O(gate285inter4));
  nand2 gate1924(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1925(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1926(.a(G660), .O(gate285inter7));
  inv1  gate1927(.a(G812), .O(gate285inter8));
  nand2 gate1928(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1929(.a(s_197), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1930(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1931(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1932(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1331(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1332(.a(gate290inter0), .b(s_112), .O(gate290inter1));
  and2  gate1333(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1334(.a(s_112), .O(gate290inter3));
  inv1  gate1335(.a(s_113), .O(gate290inter4));
  nand2 gate1336(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1337(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1338(.a(G820), .O(gate290inter7));
  inv1  gate1339(.a(G821), .O(gate290inter8));
  nand2 gate1340(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1341(.a(s_113), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1342(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1343(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1344(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1443(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1444(.a(gate387inter0), .b(s_128), .O(gate387inter1));
  and2  gate1445(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1446(.a(s_128), .O(gate387inter3));
  inv1  gate1447(.a(s_129), .O(gate387inter4));
  nand2 gate1448(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1449(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1450(.a(G1), .O(gate387inter7));
  inv1  gate1451(.a(G1036), .O(gate387inter8));
  nand2 gate1452(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1453(.a(s_129), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1454(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1455(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1456(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate2003(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2004(.a(gate390inter0), .b(s_208), .O(gate390inter1));
  and2  gate2005(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2006(.a(s_208), .O(gate390inter3));
  inv1  gate2007(.a(s_209), .O(gate390inter4));
  nand2 gate2008(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2009(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2010(.a(G4), .O(gate390inter7));
  inv1  gate2011(.a(G1045), .O(gate390inter8));
  nand2 gate2012(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2013(.a(s_209), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2014(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2015(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2016(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate645(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate646(.a(gate393inter0), .b(s_14), .O(gate393inter1));
  and2  gate647(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate648(.a(s_14), .O(gate393inter3));
  inv1  gate649(.a(s_15), .O(gate393inter4));
  nand2 gate650(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate651(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate652(.a(G7), .O(gate393inter7));
  inv1  gate653(.a(G1054), .O(gate393inter8));
  nand2 gate654(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate655(.a(s_15), .b(gate393inter3), .O(gate393inter10));
  nor2  gate656(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate657(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate658(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate575(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate576(.a(gate397inter0), .b(s_4), .O(gate397inter1));
  and2  gate577(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate578(.a(s_4), .O(gate397inter3));
  inv1  gate579(.a(s_5), .O(gate397inter4));
  nand2 gate580(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate581(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate582(.a(G11), .O(gate397inter7));
  inv1  gate583(.a(G1066), .O(gate397inter8));
  nand2 gate584(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate585(.a(s_5), .b(gate397inter3), .O(gate397inter10));
  nor2  gate586(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate587(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate588(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate701(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate702(.a(gate409inter0), .b(s_22), .O(gate409inter1));
  and2  gate703(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate704(.a(s_22), .O(gate409inter3));
  inv1  gate705(.a(s_23), .O(gate409inter4));
  nand2 gate706(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate707(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate708(.a(G23), .O(gate409inter7));
  inv1  gate709(.a(G1102), .O(gate409inter8));
  nand2 gate710(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate711(.a(s_23), .b(gate409inter3), .O(gate409inter10));
  nor2  gate712(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate713(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate714(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1121(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1122(.a(gate413inter0), .b(s_82), .O(gate413inter1));
  and2  gate1123(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1124(.a(s_82), .O(gate413inter3));
  inv1  gate1125(.a(s_83), .O(gate413inter4));
  nand2 gate1126(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1127(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1128(.a(G27), .O(gate413inter7));
  inv1  gate1129(.a(G1114), .O(gate413inter8));
  nand2 gate1130(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1131(.a(s_83), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1132(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1133(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1134(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1247(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1248(.a(gate419inter0), .b(s_100), .O(gate419inter1));
  and2  gate1249(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1250(.a(s_100), .O(gate419inter3));
  inv1  gate1251(.a(s_101), .O(gate419inter4));
  nand2 gate1252(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1253(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1254(.a(G1), .O(gate419inter7));
  inv1  gate1255(.a(G1132), .O(gate419inter8));
  nand2 gate1256(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1257(.a(s_101), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1258(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1259(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1260(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1177(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1178(.a(gate420inter0), .b(s_90), .O(gate420inter1));
  and2  gate1179(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1180(.a(s_90), .O(gate420inter3));
  inv1  gate1181(.a(s_91), .O(gate420inter4));
  nand2 gate1182(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1183(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1184(.a(G1036), .O(gate420inter7));
  inv1  gate1185(.a(G1132), .O(gate420inter8));
  nand2 gate1186(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1187(.a(s_91), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1188(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1189(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1190(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1065(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1066(.a(gate425inter0), .b(s_74), .O(gate425inter1));
  and2  gate1067(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1068(.a(s_74), .O(gate425inter3));
  inv1  gate1069(.a(s_75), .O(gate425inter4));
  nand2 gate1070(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1071(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1072(.a(G4), .O(gate425inter7));
  inv1  gate1073(.a(G1141), .O(gate425inter8));
  nand2 gate1074(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1075(.a(s_75), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1076(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1077(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1078(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1429(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1430(.a(gate426inter0), .b(s_126), .O(gate426inter1));
  and2  gate1431(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1432(.a(s_126), .O(gate426inter3));
  inv1  gate1433(.a(s_127), .O(gate426inter4));
  nand2 gate1434(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1435(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1436(.a(G1045), .O(gate426inter7));
  inv1  gate1437(.a(G1141), .O(gate426inter8));
  nand2 gate1438(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1439(.a(s_127), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1440(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1441(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1442(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1359(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1360(.a(gate427inter0), .b(s_116), .O(gate427inter1));
  and2  gate1361(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1362(.a(s_116), .O(gate427inter3));
  inv1  gate1363(.a(s_117), .O(gate427inter4));
  nand2 gate1364(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1365(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1366(.a(G5), .O(gate427inter7));
  inv1  gate1367(.a(G1144), .O(gate427inter8));
  nand2 gate1368(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1369(.a(s_117), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1370(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1371(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1372(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1807(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1808(.a(gate433inter0), .b(s_180), .O(gate433inter1));
  and2  gate1809(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1810(.a(s_180), .O(gate433inter3));
  inv1  gate1811(.a(s_181), .O(gate433inter4));
  nand2 gate1812(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1813(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1814(.a(G8), .O(gate433inter7));
  inv1  gate1815(.a(G1153), .O(gate433inter8));
  nand2 gate1816(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1817(.a(s_181), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1818(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1819(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1820(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate715(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate716(.a(gate435inter0), .b(s_24), .O(gate435inter1));
  and2  gate717(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate718(.a(s_24), .O(gate435inter3));
  inv1  gate719(.a(s_25), .O(gate435inter4));
  nand2 gate720(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate721(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate722(.a(G9), .O(gate435inter7));
  inv1  gate723(.a(G1156), .O(gate435inter8));
  nand2 gate724(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate725(.a(s_25), .b(gate435inter3), .O(gate435inter10));
  nor2  gate726(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate727(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate728(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1387(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1388(.a(gate438inter0), .b(s_120), .O(gate438inter1));
  and2  gate1389(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1390(.a(s_120), .O(gate438inter3));
  inv1  gate1391(.a(s_121), .O(gate438inter4));
  nand2 gate1392(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1393(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1394(.a(G1063), .O(gate438inter7));
  inv1  gate1395(.a(G1159), .O(gate438inter8));
  nand2 gate1396(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1397(.a(s_121), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1398(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1399(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1400(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate855(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate856(.a(gate439inter0), .b(s_44), .O(gate439inter1));
  and2  gate857(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate858(.a(s_44), .O(gate439inter3));
  inv1  gate859(.a(s_45), .O(gate439inter4));
  nand2 gate860(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate861(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate862(.a(G11), .O(gate439inter7));
  inv1  gate863(.a(G1162), .O(gate439inter8));
  nand2 gate864(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate865(.a(s_45), .b(gate439inter3), .O(gate439inter10));
  nor2  gate866(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate867(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate868(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2031(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2032(.a(gate441inter0), .b(s_212), .O(gate441inter1));
  and2  gate2033(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2034(.a(s_212), .O(gate441inter3));
  inv1  gate2035(.a(s_213), .O(gate441inter4));
  nand2 gate2036(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2037(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2038(.a(G12), .O(gate441inter7));
  inv1  gate2039(.a(G1165), .O(gate441inter8));
  nand2 gate2040(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2041(.a(s_213), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2042(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2043(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2044(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1653(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1654(.a(gate443inter0), .b(s_158), .O(gate443inter1));
  and2  gate1655(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1656(.a(s_158), .O(gate443inter3));
  inv1  gate1657(.a(s_159), .O(gate443inter4));
  nand2 gate1658(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1659(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1660(.a(G13), .O(gate443inter7));
  inv1  gate1661(.a(G1168), .O(gate443inter8));
  nand2 gate1662(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1663(.a(s_159), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1664(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1665(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1666(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1135(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1136(.a(gate447inter0), .b(s_84), .O(gate447inter1));
  and2  gate1137(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1138(.a(s_84), .O(gate447inter3));
  inv1  gate1139(.a(s_85), .O(gate447inter4));
  nand2 gate1140(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1141(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1142(.a(G15), .O(gate447inter7));
  inv1  gate1143(.a(G1174), .O(gate447inter8));
  nand2 gate1144(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1145(.a(s_85), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1146(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1147(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1148(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1877(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1878(.a(gate451inter0), .b(s_190), .O(gate451inter1));
  and2  gate1879(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1880(.a(s_190), .O(gate451inter3));
  inv1  gate1881(.a(s_191), .O(gate451inter4));
  nand2 gate1882(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1883(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1884(.a(G17), .O(gate451inter7));
  inv1  gate1885(.a(G1180), .O(gate451inter8));
  nand2 gate1886(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1887(.a(s_191), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1888(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1889(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1890(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate925(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate926(.a(gate455inter0), .b(s_54), .O(gate455inter1));
  and2  gate927(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate928(.a(s_54), .O(gate455inter3));
  inv1  gate929(.a(s_55), .O(gate455inter4));
  nand2 gate930(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate931(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate932(.a(G19), .O(gate455inter7));
  inv1  gate933(.a(G1186), .O(gate455inter8));
  nand2 gate934(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate935(.a(s_55), .b(gate455inter3), .O(gate455inter10));
  nor2  gate936(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate937(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate938(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate841(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate842(.a(gate456inter0), .b(s_42), .O(gate456inter1));
  and2  gate843(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate844(.a(s_42), .O(gate456inter3));
  inv1  gate845(.a(s_43), .O(gate456inter4));
  nand2 gate846(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate847(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate848(.a(G1090), .O(gate456inter7));
  inv1  gate849(.a(G1186), .O(gate456inter8));
  nand2 gate850(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate851(.a(s_43), .b(gate456inter3), .O(gate456inter10));
  nor2  gate852(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate853(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate854(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate617(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate618(.a(gate459inter0), .b(s_10), .O(gate459inter1));
  and2  gate619(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate620(.a(s_10), .O(gate459inter3));
  inv1  gate621(.a(s_11), .O(gate459inter4));
  nand2 gate622(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate623(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate624(.a(G21), .O(gate459inter7));
  inv1  gate625(.a(G1192), .O(gate459inter8));
  nand2 gate626(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate627(.a(s_11), .b(gate459inter3), .O(gate459inter10));
  nor2  gate628(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate629(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate630(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate967(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate968(.a(gate462inter0), .b(s_60), .O(gate462inter1));
  and2  gate969(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate970(.a(s_60), .O(gate462inter3));
  inv1  gate971(.a(s_61), .O(gate462inter4));
  nand2 gate972(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate973(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate974(.a(G1099), .O(gate462inter7));
  inv1  gate975(.a(G1195), .O(gate462inter8));
  nand2 gate976(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate977(.a(s_61), .b(gate462inter3), .O(gate462inter10));
  nor2  gate978(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate979(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate980(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1289(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1290(.a(gate463inter0), .b(s_106), .O(gate463inter1));
  and2  gate1291(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1292(.a(s_106), .O(gate463inter3));
  inv1  gate1293(.a(s_107), .O(gate463inter4));
  nand2 gate1294(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1295(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1296(.a(G23), .O(gate463inter7));
  inv1  gate1297(.a(G1198), .O(gate463inter8));
  nand2 gate1298(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1299(.a(s_107), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1300(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1301(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1302(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1107(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1108(.a(gate464inter0), .b(s_80), .O(gate464inter1));
  and2  gate1109(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1110(.a(s_80), .O(gate464inter3));
  inv1  gate1111(.a(s_81), .O(gate464inter4));
  nand2 gate1112(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1113(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1114(.a(G1102), .O(gate464inter7));
  inv1  gate1115(.a(G1198), .O(gate464inter8));
  nand2 gate1116(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1117(.a(s_81), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1118(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1119(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1120(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate743(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate744(.a(gate465inter0), .b(s_28), .O(gate465inter1));
  and2  gate745(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate746(.a(s_28), .O(gate465inter3));
  inv1  gate747(.a(s_29), .O(gate465inter4));
  nand2 gate748(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate749(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate750(.a(G24), .O(gate465inter7));
  inv1  gate751(.a(G1201), .O(gate465inter8));
  nand2 gate752(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate753(.a(s_29), .b(gate465inter3), .O(gate465inter10));
  nor2  gate754(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate755(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate756(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1569(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1570(.a(gate466inter0), .b(s_146), .O(gate466inter1));
  and2  gate1571(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1572(.a(s_146), .O(gate466inter3));
  inv1  gate1573(.a(s_147), .O(gate466inter4));
  nand2 gate1574(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1575(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1576(.a(G1105), .O(gate466inter7));
  inv1  gate1577(.a(G1201), .O(gate466inter8));
  nand2 gate1578(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1579(.a(s_147), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1580(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1581(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1582(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate729(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate730(.a(gate478inter0), .b(s_26), .O(gate478inter1));
  and2  gate731(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate732(.a(s_26), .O(gate478inter3));
  inv1  gate733(.a(s_27), .O(gate478inter4));
  nand2 gate734(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate735(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate736(.a(G1123), .O(gate478inter7));
  inv1  gate737(.a(G1219), .O(gate478inter8));
  nand2 gate738(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate739(.a(s_27), .b(gate478inter3), .O(gate478inter10));
  nor2  gate740(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate741(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate742(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1219(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1220(.a(gate486inter0), .b(s_96), .O(gate486inter1));
  and2  gate1221(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1222(.a(s_96), .O(gate486inter3));
  inv1  gate1223(.a(s_97), .O(gate486inter4));
  nand2 gate1224(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1225(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1226(.a(G1234), .O(gate486inter7));
  inv1  gate1227(.a(G1235), .O(gate486inter8));
  nand2 gate1228(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1229(.a(s_97), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1230(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1231(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1232(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1527(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1528(.a(gate489inter0), .b(s_140), .O(gate489inter1));
  and2  gate1529(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1530(.a(s_140), .O(gate489inter3));
  inv1  gate1531(.a(s_141), .O(gate489inter4));
  nand2 gate1532(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1533(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1534(.a(G1240), .O(gate489inter7));
  inv1  gate1535(.a(G1241), .O(gate489inter8));
  nand2 gate1536(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1537(.a(s_141), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1538(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1539(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1540(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1611(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1612(.a(gate496inter0), .b(s_152), .O(gate496inter1));
  and2  gate1613(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1614(.a(s_152), .O(gate496inter3));
  inv1  gate1615(.a(s_153), .O(gate496inter4));
  nand2 gate1616(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1617(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1618(.a(G1254), .O(gate496inter7));
  inv1  gate1619(.a(G1255), .O(gate496inter8));
  nand2 gate1620(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1621(.a(s_153), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1622(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1623(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1624(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1597(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1598(.a(gate501inter0), .b(s_150), .O(gate501inter1));
  and2  gate1599(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1600(.a(s_150), .O(gate501inter3));
  inv1  gate1601(.a(s_151), .O(gate501inter4));
  nand2 gate1602(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1603(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1604(.a(G1264), .O(gate501inter7));
  inv1  gate1605(.a(G1265), .O(gate501inter8));
  nand2 gate1606(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1607(.a(s_151), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1608(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1609(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1610(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate757(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate758(.a(gate503inter0), .b(s_30), .O(gate503inter1));
  and2  gate759(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate760(.a(s_30), .O(gate503inter3));
  inv1  gate761(.a(s_31), .O(gate503inter4));
  nand2 gate762(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate763(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate764(.a(G1268), .O(gate503inter7));
  inv1  gate765(.a(G1269), .O(gate503inter8));
  nand2 gate766(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate767(.a(s_31), .b(gate503inter3), .O(gate503inter10));
  nor2  gate768(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate769(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate770(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1485(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1486(.a(gate506inter0), .b(s_134), .O(gate506inter1));
  and2  gate1487(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1488(.a(s_134), .O(gate506inter3));
  inv1  gate1489(.a(s_135), .O(gate506inter4));
  nand2 gate1490(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1491(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1492(.a(G1274), .O(gate506inter7));
  inv1  gate1493(.a(G1275), .O(gate506inter8));
  nand2 gate1494(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1495(.a(s_135), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1496(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1497(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1498(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate1149(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1150(.a(gate508inter0), .b(s_86), .O(gate508inter1));
  and2  gate1151(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1152(.a(s_86), .O(gate508inter3));
  inv1  gate1153(.a(s_87), .O(gate508inter4));
  nand2 gate1154(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1155(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1156(.a(G1278), .O(gate508inter7));
  inv1  gate1157(.a(G1279), .O(gate508inter8));
  nand2 gate1158(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1159(.a(s_87), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1160(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1161(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1162(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2073(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2074(.a(gate509inter0), .b(s_218), .O(gate509inter1));
  and2  gate2075(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2076(.a(s_218), .O(gate509inter3));
  inv1  gate2077(.a(s_219), .O(gate509inter4));
  nand2 gate2078(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2079(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2080(.a(G1280), .O(gate509inter7));
  inv1  gate2081(.a(G1281), .O(gate509inter8));
  nand2 gate2082(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2083(.a(s_219), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2084(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2085(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2086(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1163(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1164(.a(gate510inter0), .b(s_88), .O(gate510inter1));
  and2  gate1165(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1166(.a(s_88), .O(gate510inter3));
  inv1  gate1167(.a(s_89), .O(gate510inter4));
  nand2 gate1168(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1169(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1170(.a(G1282), .O(gate510inter7));
  inv1  gate1171(.a(G1283), .O(gate510inter8));
  nand2 gate1172(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1173(.a(s_89), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1174(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1175(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1176(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate603(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate604(.a(gate511inter0), .b(s_8), .O(gate511inter1));
  and2  gate605(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate606(.a(s_8), .O(gate511inter3));
  inv1  gate607(.a(s_9), .O(gate511inter4));
  nand2 gate608(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate609(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate610(.a(G1284), .O(gate511inter7));
  inv1  gate611(.a(G1285), .O(gate511inter8));
  nand2 gate612(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate613(.a(s_9), .b(gate511inter3), .O(gate511inter10));
  nor2  gate614(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate615(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate616(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule