module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );

  xor2  gate469(.a(N85), .b(N81), .O(gate11inter0));
  nand2 gate470(.a(gate11inter0), .b(s_38), .O(gate11inter1));
  and2  gate471(.a(N85), .b(N81), .O(gate11inter2));
  inv1  gate472(.a(s_38), .O(gate11inter3));
  inv1  gate473(.a(s_39), .O(gate11inter4));
  nand2 gate474(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate475(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate476(.a(N81), .O(gate11inter7));
  inv1  gate477(.a(N85), .O(gate11inter8));
  nand2 gate478(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate479(.a(s_39), .b(gate11inter3), .O(gate11inter10));
  nor2  gate480(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate481(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate482(.a(gate11inter12), .b(gate11inter1), .O(N260));

  xor2  gate427(.a(N93), .b(N89), .O(gate12inter0));
  nand2 gate428(.a(gate12inter0), .b(s_32), .O(gate12inter1));
  and2  gate429(.a(N93), .b(N89), .O(gate12inter2));
  inv1  gate430(.a(s_32), .O(gate12inter3));
  inv1  gate431(.a(s_33), .O(gate12inter4));
  nand2 gate432(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate433(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate434(.a(N89), .O(gate12inter7));
  inv1  gate435(.a(N93), .O(gate12inter8));
  nand2 gate436(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate437(.a(s_33), .b(gate12inter3), .O(gate12inter10));
  nor2  gate438(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate439(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate440(.a(gate12inter12), .b(gate12inter1), .O(N261));
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate399(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate400(.a(gate25inter0), .b(s_28), .O(gate25inter1));
  and2  gate401(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate402(.a(s_28), .O(gate25inter3));
  inv1  gate403(.a(s_29), .O(gate25inter4));
  nand2 gate404(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate405(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate406(.a(N1), .O(gate25inter7));
  inv1  gate407(.a(N17), .O(gate25inter8));
  nand2 gate408(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate409(.a(s_29), .b(gate25inter3), .O(gate25inter10));
  nor2  gate410(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate411(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate412(.a(gate25inter12), .b(gate25inter1), .O(N274));

  xor2  gate357(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate358(.a(gate26inter0), .b(s_22), .O(gate26inter1));
  and2  gate359(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate360(.a(s_22), .O(gate26inter3));
  inv1  gate361(.a(s_23), .O(gate26inter4));
  nand2 gate362(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate363(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate364(.a(N33), .O(gate26inter7));
  inv1  gate365(.a(N49), .O(gate26inter8));
  nand2 gate366(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate367(.a(s_23), .b(gate26inter3), .O(gate26inter10));
  nor2  gate368(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate369(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate370(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );

  xor2  gate371(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate372(.a(gate28inter0), .b(s_24), .O(gate28inter1));
  and2  gate373(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate374(.a(s_24), .O(gate28inter3));
  inv1  gate375(.a(s_25), .O(gate28inter4));
  nand2 gate376(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate377(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate378(.a(N37), .O(gate28inter7));
  inv1  gate379(.a(N53), .O(gate28inter8));
  nand2 gate380(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate381(.a(s_25), .b(gate28inter3), .O(gate28inter10));
  nor2  gate382(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate383(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate384(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate343(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate344(.a(gate30inter0), .b(s_20), .O(gate30inter1));
  and2  gate345(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate346(.a(s_20), .O(gate30inter3));
  inv1  gate347(.a(s_21), .O(gate30inter4));
  nand2 gate348(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate349(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate350(.a(N41), .O(gate30inter7));
  inv1  gate351(.a(N57), .O(gate30inter8));
  nand2 gate352(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate353(.a(s_21), .b(gate30inter3), .O(gate30inter10));
  nor2  gate354(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate355(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate356(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );

  xor2  gate217(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate218(.a(gate40inter0), .b(s_2), .O(gate40inter1));
  and2  gate219(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate220(.a(s_2), .O(gate40inter3));
  inv1  gate221(.a(s_3), .O(gate40inter4));
  nand2 gate222(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate223(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate224(.a(N109), .O(gate40inter7));
  inv1  gate225(.a(N125), .O(gate40inter8));
  nand2 gate226(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate227(.a(s_3), .b(gate40inter3), .O(gate40inter10));
  nor2  gate228(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate229(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate230(.a(gate40inter12), .b(gate40inter1), .O(N289));
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );

  xor2  gate301(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate302(.a(gate43inter0), .b(s_14), .O(gate43inter1));
  and2  gate303(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate304(.a(s_14), .O(gate43inter3));
  inv1  gate305(.a(s_15), .O(gate43inter4));
  nand2 gate306(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate307(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate308(.a(N254), .O(gate43inter7));
  inv1  gate309(.a(N255), .O(gate43inter8));
  nand2 gate310(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate311(.a(s_15), .b(gate43inter3), .O(gate43inter10));
  nor2  gate312(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate313(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate314(.a(gate43inter12), .b(gate43inter1), .O(N296));

  xor2  gate329(.a(N257), .b(N256), .O(gate44inter0));
  nand2 gate330(.a(gate44inter0), .b(s_18), .O(gate44inter1));
  and2  gate331(.a(N257), .b(N256), .O(gate44inter2));
  inv1  gate332(.a(s_18), .O(gate44inter3));
  inv1  gate333(.a(s_19), .O(gate44inter4));
  nand2 gate334(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate335(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate336(.a(N256), .O(gate44inter7));
  inv1  gate337(.a(N257), .O(gate44inter8));
  nand2 gate338(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate339(.a(s_19), .b(gate44inter3), .O(gate44inter10));
  nor2  gate340(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate341(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate342(.a(gate44inter12), .b(gate44inter1), .O(N299));
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate553(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate554(.a(gate47inter0), .b(s_50), .O(gate47inter1));
  and2  gate555(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate556(.a(s_50), .O(gate47inter3));
  inv1  gate557(.a(s_51), .O(gate47inter4));
  nand2 gate558(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate559(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate560(.a(N262), .O(gate47inter7));
  inv1  gate561(.a(N263), .O(gate47inter8));
  nand2 gate562(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate563(.a(s_51), .b(gate47inter3), .O(gate47inter10));
  nor2  gate564(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate565(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate566(.a(gate47inter12), .b(gate47inter1), .O(N308));
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );

  xor2  gate273(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate274(.a(gate57inter0), .b(s_10), .O(gate57inter1));
  and2  gate275(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate276(.a(s_10), .O(gate57inter3));
  inv1  gate277(.a(s_11), .O(gate57inter4));
  nand2 gate278(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate279(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate280(.a(N290), .O(gate57inter7));
  inv1  gate281(.a(N293), .O(gate57inter8));
  nand2 gate282(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate283(.a(s_11), .b(gate57inter3), .O(gate57inter10));
  nor2  gate284(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate285(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate286(.a(gate57inter12), .b(gate57inter1), .O(N338));

  xor2  gate231(.a(N299), .b(N296), .O(gate58inter0));
  nand2 gate232(.a(gate58inter0), .b(s_4), .O(gate58inter1));
  and2  gate233(.a(N299), .b(N296), .O(gate58inter2));
  inv1  gate234(.a(s_4), .O(gate58inter3));
  inv1  gate235(.a(s_5), .O(gate58inter4));
  nand2 gate236(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate237(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate238(.a(N296), .O(gate58inter7));
  inv1  gate239(.a(N299), .O(gate58inter8));
  nand2 gate240(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate241(.a(s_5), .b(gate58inter3), .O(gate58inter10));
  nor2  gate242(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate243(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate244(.a(gate58inter12), .b(gate58inter1), .O(N339));
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );

  xor2  gate441(.a(N305), .b(N302), .O(gate61inter0));
  nand2 gate442(.a(gate61inter0), .b(s_34), .O(gate61inter1));
  and2  gate443(.a(N305), .b(N302), .O(gate61inter2));
  inv1  gate444(.a(s_34), .O(gate61inter3));
  inv1  gate445(.a(s_35), .O(gate61inter4));
  nand2 gate446(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate447(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate448(.a(N302), .O(gate61inter7));
  inv1  gate449(.a(N305), .O(gate61inter8));
  nand2 gate450(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate451(.a(s_35), .b(gate61inter3), .O(gate61inter10));
  nor2  gate452(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate453(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate454(.a(gate61inter12), .b(gate61inter1), .O(N342));
xor2 gate62( .a(N308), .b(N311), .O(N343) );

  xor2  gate385(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate386(.a(gate63inter0), .b(s_26), .O(gate63inter1));
  and2  gate387(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate388(.a(s_26), .O(gate63inter3));
  inv1  gate389(.a(s_27), .O(gate63inter4));
  nand2 gate390(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate391(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate392(.a(N302), .O(gate63inter7));
  inv1  gate393(.a(N308), .O(gate63inter8));
  nand2 gate394(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate395(.a(s_27), .b(gate63inter3), .O(gate63inter10));
  nor2  gate396(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate397(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate398(.a(gate63inter12), .b(gate63inter1), .O(N344));
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );

  xor2  gate455(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate456(.a(gate67inter0), .b(s_36), .O(gate67inter1));
  and2  gate457(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate458(.a(s_36), .O(gate67inter3));
  inv1  gate459(.a(s_37), .O(gate67inter4));
  nand2 gate460(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate461(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate462(.a(N268), .O(gate67inter7));
  inv1  gate463(.a(N344), .O(gate67inter8));
  nand2 gate464(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate465(.a(s_37), .b(gate67inter3), .O(gate67inter10));
  nor2  gate466(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate467(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate468(.a(gate67inter12), .b(gate67inter1), .O(N348));
xor2 gate68( .a(N269), .b(N345), .O(N349) );

  xor2  gate315(.a(N338), .b(N270), .O(gate69inter0));
  nand2 gate316(.a(gate69inter0), .b(s_16), .O(gate69inter1));
  and2  gate317(.a(N338), .b(N270), .O(gate69inter2));
  inv1  gate318(.a(s_16), .O(gate69inter3));
  inv1  gate319(.a(s_17), .O(gate69inter4));
  nand2 gate320(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate321(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate322(.a(N270), .O(gate69inter7));
  inv1  gate323(.a(N338), .O(gate69inter8));
  nand2 gate324(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate325(.a(s_17), .b(gate69inter3), .O(gate69inter10));
  nor2  gate326(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate327(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate328(.a(gate69inter12), .b(gate69inter1), .O(N350));
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );

  xor2  gate287(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate288(.a(gate77inter0), .b(s_12), .O(gate77inter1));
  and2  gate289(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate290(.a(s_12), .O(gate77inter3));
  inv1  gate291(.a(s_13), .O(gate77inter4));
  nand2 gate292(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate293(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate294(.a(N318), .O(gate77inter7));
  inv1  gate295(.a(N350), .O(gate77inter8));
  nand2 gate296(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate297(.a(s_13), .b(gate77inter3), .O(gate77inter10));
  nor2  gate298(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate299(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate300(.a(gate77inter12), .b(gate77inter1), .O(N406));
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate539(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate540(.a(gate177inter0), .b(s_48), .O(gate177inter1));
  and2  gate541(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate542(.a(s_48), .O(gate177inter3));
  inv1  gate543(.a(s_49), .O(gate177inter4));
  nand2 gate544(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate545(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate546(.a(N25), .O(gate177inter7));
  inv1  gate547(.a(N698), .O(gate177inter8));
  nand2 gate548(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate549(.a(s_49), .b(gate177inter3), .O(gate177inter10));
  nor2  gate550(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate551(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate552(.a(gate177inter12), .b(gate177inter1), .O(N730));
xor2 gate178( .a(N29), .b(N699), .O(N731) );

  xor2  gate413(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate414(.a(gate179inter0), .b(s_30), .O(gate179inter1));
  and2  gate415(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate416(.a(s_30), .O(gate179inter3));
  inv1  gate417(.a(s_31), .O(gate179inter4));
  nand2 gate418(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate419(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate420(.a(N33), .O(gate179inter7));
  inv1  gate421(.a(N700), .O(gate179inter8));
  nand2 gate422(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate423(.a(s_31), .b(gate179inter3), .O(gate179inter10));
  nor2  gate424(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate425(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate426(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );

  xor2  gate245(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate246(.a(gate182inter0), .b(s_6), .O(gate182inter1));
  and2  gate247(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate248(.a(s_6), .O(gate182inter3));
  inv1  gate249(.a(s_7), .O(gate182inter4));
  nand2 gate250(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate251(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate252(.a(N45), .O(gate182inter7));
  inv1  gate253(.a(N703), .O(gate182inter8));
  nand2 gate254(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate255(.a(s_7), .b(gate182inter3), .O(gate182inter10));
  nor2  gate256(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate257(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate258(.a(gate182inter12), .b(gate182inter1), .O(N735));

  xor2  gate525(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate526(.a(gate183inter0), .b(s_46), .O(gate183inter1));
  and2  gate527(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate528(.a(s_46), .O(gate183inter3));
  inv1  gate529(.a(s_47), .O(gate183inter4));
  nand2 gate530(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate531(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate532(.a(N49), .O(gate183inter7));
  inv1  gate533(.a(N704), .O(gate183inter8));
  nand2 gate534(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate535(.a(s_47), .b(gate183inter3), .O(gate183inter10));
  nor2  gate536(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate537(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate538(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );

  xor2  gate203(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate204(.a(gate186inter0), .b(s_0), .O(gate186inter1));
  and2  gate205(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate206(.a(s_0), .O(gate186inter3));
  inv1  gate207(.a(s_1), .O(gate186inter4));
  nand2 gate208(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate209(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate210(.a(N61), .O(gate186inter7));
  inv1  gate211(.a(N707), .O(gate186inter8));
  nand2 gate212(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate213(.a(s_1), .b(gate186inter3), .O(gate186inter10));
  nor2  gate214(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate215(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate216(.a(gate186inter12), .b(gate186inter1), .O(N739));
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );

  xor2  gate497(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate498(.a(gate192inter0), .b(s_42), .O(gate192inter1));
  and2  gate499(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate500(.a(s_42), .O(gate192inter3));
  inv1  gate501(.a(s_43), .O(gate192inter4));
  nand2 gate502(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate503(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate504(.a(N85), .O(gate192inter7));
  inv1  gate505(.a(N713), .O(gate192inter8));
  nand2 gate506(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate507(.a(s_43), .b(gate192inter3), .O(gate192inter10));
  nor2  gate508(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate509(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate510(.a(gate192inter12), .b(gate192inter1), .O(N745));

  xor2  gate259(.a(N714), .b(N89), .O(gate193inter0));
  nand2 gate260(.a(gate193inter0), .b(s_8), .O(gate193inter1));
  and2  gate261(.a(N714), .b(N89), .O(gate193inter2));
  inv1  gate262(.a(s_8), .O(gate193inter3));
  inv1  gate263(.a(s_9), .O(gate193inter4));
  nand2 gate264(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate265(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate266(.a(N89), .O(gate193inter7));
  inv1  gate267(.a(N714), .O(gate193inter8));
  nand2 gate268(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate269(.a(s_9), .b(gate193inter3), .O(gate193inter10));
  nor2  gate270(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate271(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate272(.a(gate193inter12), .b(gate193inter1), .O(N746));
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );

  xor2  gate511(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate512(.a(gate196inter0), .b(s_44), .O(gate196inter1));
  and2  gate513(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate514(.a(s_44), .O(gate196inter3));
  inv1  gate515(.a(s_45), .O(gate196inter4));
  nand2 gate516(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate517(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate518(.a(N101), .O(gate196inter7));
  inv1  gate519(.a(N717), .O(gate196inter8));
  nand2 gate520(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate521(.a(s_45), .b(gate196inter3), .O(gate196inter10));
  nor2  gate522(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate523(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate524(.a(gate196inter12), .b(gate196inter1), .O(N749));
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );

  xor2  gate483(.a(N720), .b(N113), .O(gate199inter0));
  nand2 gate484(.a(gate199inter0), .b(s_40), .O(gate199inter1));
  and2  gate485(.a(N720), .b(N113), .O(gate199inter2));
  inv1  gate486(.a(s_40), .O(gate199inter3));
  inv1  gate487(.a(s_41), .O(gate199inter4));
  nand2 gate488(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate489(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate490(.a(N113), .O(gate199inter7));
  inv1  gate491(.a(N720), .O(gate199inter8));
  nand2 gate492(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate493(.a(s_41), .b(gate199inter3), .O(gate199inter10));
  nor2  gate494(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate495(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate496(.a(gate199inter12), .b(gate199inter1), .O(N752));
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule