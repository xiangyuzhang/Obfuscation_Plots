module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate743(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate744(.a(gate19inter0), .b(s_28), .O(gate19inter1));
  and2  gate745(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate746(.a(s_28), .O(gate19inter3));
  inv1  gate747(.a(s_29), .O(gate19inter4));
  nand2 gate748(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate749(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate750(.a(G21), .O(gate19inter7));
  inv1  gate751(.a(G22), .O(gate19inter8));
  nand2 gate752(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate753(.a(s_29), .b(gate19inter3), .O(gate19inter10));
  nor2  gate754(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate755(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate756(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1457(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1458(.a(gate33inter0), .b(s_130), .O(gate33inter1));
  and2  gate1459(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1460(.a(s_130), .O(gate33inter3));
  inv1  gate1461(.a(s_131), .O(gate33inter4));
  nand2 gate1462(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1463(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1464(.a(G17), .O(gate33inter7));
  inv1  gate1465(.a(G21), .O(gate33inter8));
  nand2 gate1466(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1467(.a(s_131), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1468(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1469(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1470(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1639(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1640(.a(gate36inter0), .b(s_156), .O(gate36inter1));
  and2  gate1641(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1642(.a(s_156), .O(gate36inter3));
  inv1  gate1643(.a(s_157), .O(gate36inter4));
  nand2 gate1644(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1645(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1646(.a(G26), .O(gate36inter7));
  inv1  gate1647(.a(G30), .O(gate36inter8));
  nand2 gate1648(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1649(.a(s_157), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1650(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1651(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1652(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1303(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1304(.a(gate40inter0), .b(s_108), .O(gate40inter1));
  and2  gate1305(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1306(.a(s_108), .O(gate40inter3));
  inv1  gate1307(.a(s_109), .O(gate40inter4));
  nand2 gate1308(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1309(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1310(.a(G28), .O(gate40inter7));
  inv1  gate1311(.a(G32), .O(gate40inter8));
  nand2 gate1312(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1313(.a(s_109), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1314(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1315(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1316(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1555(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1556(.a(gate45inter0), .b(s_144), .O(gate45inter1));
  and2  gate1557(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1558(.a(s_144), .O(gate45inter3));
  inv1  gate1559(.a(s_145), .O(gate45inter4));
  nand2 gate1560(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1561(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1562(.a(G5), .O(gate45inter7));
  inv1  gate1563(.a(G272), .O(gate45inter8));
  nand2 gate1564(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1565(.a(s_145), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1566(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1567(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1568(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1009(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1010(.a(gate54inter0), .b(s_66), .O(gate54inter1));
  and2  gate1011(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1012(.a(s_66), .O(gate54inter3));
  inv1  gate1013(.a(s_67), .O(gate54inter4));
  nand2 gate1014(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1015(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1016(.a(G14), .O(gate54inter7));
  inv1  gate1017(.a(G284), .O(gate54inter8));
  nand2 gate1018(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1019(.a(s_67), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1020(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1021(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1022(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate911(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate912(.a(gate57inter0), .b(s_52), .O(gate57inter1));
  and2  gate913(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate914(.a(s_52), .O(gate57inter3));
  inv1  gate915(.a(s_53), .O(gate57inter4));
  nand2 gate916(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate917(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate918(.a(G17), .O(gate57inter7));
  inv1  gate919(.a(G290), .O(gate57inter8));
  nand2 gate920(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate921(.a(s_53), .b(gate57inter3), .O(gate57inter10));
  nor2  gate922(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate923(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate924(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1233(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1234(.a(gate62inter0), .b(s_98), .O(gate62inter1));
  and2  gate1235(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1236(.a(s_98), .O(gate62inter3));
  inv1  gate1237(.a(s_99), .O(gate62inter4));
  nand2 gate1238(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1239(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1240(.a(G22), .O(gate62inter7));
  inv1  gate1241(.a(G296), .O(gate62inter8));
  nand2 gate1242(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1243(.a(s_99), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1244(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1245(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1246(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1317(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1318(.a(gate63inter0), .b(s_110), .O(gate63inter1));
  and2  gate1319(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1320(.a(s_110), .O(gate63inter3));
  inv1  gate1321(.a(s_111), .O(gate63inter4));
  nand2 gate1322(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1323(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1324(.a(G23), .O(gate63inter7));
  inv1  gate1325(.a(G299), .O(gate63inter8));
  nand2 gate1326(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1327(.a(s_111), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1328(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1329(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1330(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate995(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate996(.a(gate66inter0), .b(s_64), .O(gate66inter1));
  and2  gate997(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate998(.a(s_64), .O(gate66inter3));
  inv1  gate999(.a(s_65), .O(gate66inter4));
  nand2 gate1000(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1001(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1002(.a(G26), .O(gate66inter7));
  inv1  gate1003(.a(G302), .O(gate66inter8));
  nand2 gate1004(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1005(.a(s_65), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1006(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1007(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1008(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1135(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1136(.a(gate68inter0), .b(s_84), .O(gate68inter1));
  and2  gate1137(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1138(.a(s_84), .O(gate68inter3));
  inv1  gate1139(.a(s_85), .O(gate68inter4));
  nand2 gate1140(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1141(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1142(.a(G28), .O(gate68inter7));
  inv1  gate1143(.a(G305), .O(gate68inter8));
  nand2 gate1144(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1145(.a(s_85), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1146(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1147(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1148(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1597(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1598(.a(gate70inter0), .b(s_150), .O(gate70inter1));
  and2  gate1599(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1600(.a(s_150), .O(gate70inter3));
  inv1  gate1601(.a(s_151), .O(gate70inter4));
  nand2 gate1602(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1603(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1604(.a(G30), .O(gate70inter7));
  inv1  gate1605(.a(G308), .O(gate70inter8));
  nand2 gate1606(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1607(.a(s_151), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1608(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1609(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1610(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1485(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1486(.a(gate74inter0), .b(s_134), .O(gate74inter1));
  and2  gate1487(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1488(.a(s_134), .O(gate74inter3));
  inv1  gate1489(.a(s_135), .O(gate74inter4));
  nand2 gate1490(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1491(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1492(.a(G5), .O(gate74inter7));
  inv1  gate1493(.a(G314), .O(gate74inter8));
  nand2 gate1494(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1495(.a(s_135), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1496(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1497(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1498(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate883(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate884(.a(gate82inter0), .b(s_48), .O(gate82inter1));
  and2  gate885(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate886(.a(s_48), .O(gate82inter3));
  inv1  gate887(.a(s_49), .O(gate82inter4));
  nand2 gate888(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate889(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate890(.a(G7), .O(gate82inter7));
  inv1  gate891(.a(G326), .O(gate82inter8));
  nand2 gate892(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate893(.a(s_49), .b(gate82inter3), .O(gate82inter10));
  nor2  gate894(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate895(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate896(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate645(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate646(.a(gate83inter0), .b(s_14), .O(gate83inter1));
  and2  gate647(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate648(.a(s_14), .O(gate83inter3));
  inv1  gate649(.a(s_15), .O(gate83inter4));
  nand2 gate650(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate651(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate652(.a(G11), .O(gate83inter7));
  inv1  gate653(.a(G329), .O(gate83inter8));
  nand2 gate654(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate655(.a(s_15), .b(gate83inter3), .O(gate83inter10));
  nor2  gate656(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate657(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate658(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate561(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate562(.a(gate93inter0), .b(s_2), .O(gate93inter1));
  and2  gate563(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate564(.a(s_2), .O(gate93inter3));
  inv1  gate565(.a(s_3), .O(gate93inter4));
  nand2 gate566(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate567(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate568(.a(G18), .O(gate93inter7));
  inv1  gate569(.a(G344), .O(gate93inter8));
  nand2 gate570(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate571(.a(s_3), .b(gate93inter3), .O(gate93inter10));
  nor2  gate572(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate573(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate574(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1051(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1052(.a(gate96inter0), .b(s_72), .O(gate96inter1));
  and2  gate1053(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1054(.a(s_72), .O(gate96inter3));
  inv1  gate1055(.a(s_73), .O(gate96inter4));
  nand2 gate1056(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1057(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1058(.a(G30), .O(gate96inter7));
  inv1  gate1059(.a(G347), .O(gate96inter8));
  nand2 gate1060(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1061(.a(s_73), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1062(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1063(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1064(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1611(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1612(.a(gate110inter0), .b(s_152), .O(gate110inter1));
  and2  gate1613(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1614(.a(s_152), .O(gate110inter3));
  inv1  gate1615(.a(s_153), .O(gate110inter4));
  nand2 gate1616(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1617(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1618(.a(G372), .O(gate110inter7));
  inv1  gate1619(.a(G373), .O(gate110inter8));
  nand2 gate1620(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1621(.a(s_153), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1622(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1623(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1624(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1471(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1472(.a(gate111inter0), .b(s_132), .O(gate111inter1));
  and2  gate1473(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1474(.a(s_132), .O(gate111inter3));
  inv1  gate1475(.a(s_133), .O(gate111inter4));
  nand2 gate1476(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1477(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1478(.a(G374), .O(gate111inter7));
  inv1  gate1479(.a(G375), .O(gate111inter8));
  nand2 gate1480(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1481(.a(s_133), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1482(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1483(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1484(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1247(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1248(.a(gate117inter0), .b(s_100), .O(gate117inter1));
  and2  gate1249(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1250(.a(s_100), .O(gate117inter3));
  inv1  gate1251(.a(s_101), .O(gate117inter4));
  nand2 gate1252(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1253(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1254(.a(G386), .O(gate117inter7));
  inv1  gate1255(.a(G387), .O(gate117inter8));
  nand2 gate1256(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1257(.a(s_101), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1258(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1259(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1260(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate673(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate674(.a(gate122inter0), .b(s_18), .O(gate122inter1));
  and2  gate675(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate676(.a(s_18), .O(gate122inter3));
  inv1  gate677(.a(s_19), .O(gate122inter4));
  nand2 gate678(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate679(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate680(.a(G396), .O(gate122inter7));
  inv1  gate681(.a(G397), .O(gate122inter8));
  nand2 gate682(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate683(.a(s_19), .b(gate122inter3), .O(gate122inter10));
  nor2  gate684(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate685(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate686(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate575(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate576(.a(gate123inter0), .b(s_4), .O(gate123inter1));
  and2  gate577(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate578(.a(s_4), .O(gate123inter3));
  inv1  gate579(.a(s_5), .O(gate123inter4));
  nand2 gate580(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate581(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate582(.a(G398), .O(gate123inter7));
  inv1  gate583(.a(G399), .O(gate123inter8));
  nand2 gate584(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate585(.a(s_5), .b(gate123inter3), .O(gate123inter10));
  nor2  gate586(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate587(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate588(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate827(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate828(.a(gate127inter0), .b(s_40), .O(gate127inter1));
  and2  gate829(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate830(.a(s_40), .O(gate127inter3));
  inv1  gate831(.a(s_41), .O(gate127inter4));
  nand2 gate832(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate833(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate834(.a(G406), .O(gate127inter7));
  inv1  gate835(.a(G407), .O(gate127inter8));
  nand2 gate836(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate837(.a(s_41), .b(gate127inter3), .O(gate127inter10));
  nor2  gate838(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate839(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate840(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate841(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate842(.a(gate128inter0), .b(s_42), .O(gate128inter1));
  and2  gate843(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate844(.a(s_42), .O(gate128inter3));
  inv1  gate845(.a(s_43), .O(gate128inter4));
  nand2 gate846(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate847(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate848(.a(G408), .O(gate128inter7));
  inv1  gate849(.a(G409), .O(gate128inter8));
  nand2 gate850(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate851(.a(s_43), .b(gate128inter3), .O(gate128inter10));
  nor2  gate852(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate853(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate854(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1415(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1416(.a(gate129inter0), .b(s_124), .O(gate129inter1));
  and2  gate1417(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1418(.a(s_124), .O(gate129inter3));
  inv1  gate1419(.a(s_125), .O(gate129inter4));
  nand2 gate1420(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1421(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1422(.a(G410), .O(gate129inter7));
  inv1  gate1423(.a(G411), .O(gate129inter8));
  nand2 gate1424(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1425(.a(s_125), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1426(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1427(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1428(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1107(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1108(.a(gate140inter0), .b(s_80), .O(gate140inter1));
  and2  gate1109(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1110(.a(s_80), .O(gate140inter3));
  inv1  gate1111(.a(s_81), .O(gate140inter4));
  nand2 gate1112(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1113(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1114(.a(G444), .O(gate140inter7));
  inv1  gate1115(.a(G447), .O(gate140inter8));
  nand2 gate1116(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1117(.a(s_81), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1118(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1119(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1120(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1163(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1164(.a(gate144inter0), .b(s_88), .O(gate144inter1));
  and2  gate1165(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1166(.a(s_88), .O(gate144inter3));
  inv1  gate1167(.a(s_89), .O(gate144inter4));
  nand2 gate1168(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1169(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1170(.a(G468), .O(gate144inter7));
  inv1  gate1171(.a(G471), .O(gate144inter8));
  nand2 gate1172(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1173(.a(s_89), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1174(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1175(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1176(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1177(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1178(.a(gate147inter0), .b(s_90), .O(gate147inter1));
  and2  gate1179(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1180(.a(s_90), .O(gate147inter3));
  inv1  gate1181(.a(s_91), .O(gate147inter4));
  nand2 gate1182(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1183(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1184(.a(G486), .O(gate147inter7));
  inv1  gate1185(.a(G489), .O(gate147inter8));
  nand2 gate1186(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1187(.a(s_91), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1188(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1189(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1190(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate631(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate632(.a(gate148inter0), .b(s_12), .O(gate148inter1));
  and2  gate633(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate634(.a(s_12), .O(gate148inter3));
  inv1  gate635(.a(s_13), .O(gate148inter4));
  nand2 gate636(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate637(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate638(.a(G492), .O(gate148inter7));
  inv1  gate639(.a(G495), .O(gate148inter8));
  nand2 gate640(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate641(.a(s_13), .b(gate148inter3), .O(gate148inter10));
  nor2  gate642(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate643(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate644(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1191(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1192(.a(gate150inter0), .b(s_92), .O(gate150inter1));
  and2  gate1193(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1194(.a(s_92), .O(gate150inter3));
  inv1  gate1195(.a(s_93), .O(gate150inter4));
  nand2 gate1196(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1197(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1198(.a(G504), .O(gate150inter7));
  inv1  gate1199(.a(G507), .O(gate150inter8));
  nand2 gate1200(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1201(.a(s_93), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1202(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1203(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1204(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate1429(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1430(.a(gate151inter0), .b(s_126), .O(gate151inter1));
  and2  gate1431(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1432(.a(s_126), .O(gate151inter3));
  inv1  gate1433(.a(s_127), .O(gate151inter4));
  nand2 gate1434(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1435(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1436(.a(G510), .O(gate151inter7));
  inv1  gate1437(.a(G513), .O(gate151inter8));
  nand2 gate1438(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1439(.a(s_127), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1440(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1441(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1442(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1569(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1570(.a(gate156inter0), .b(s_146), .O(gate156inter1));
  and2  gate1571(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1572(.a(s_146), .O(gate156inter3));
  inv1  gate1573(.a(s_147), .O(gate156inter4));
  nand2 gate1574(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1575(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1576(.a(G435), .O(gate156inter7));
  inv1  gate1577(.a(G525), .O(gate156inter8));
  nand2 gate1578(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1579(.a(s_147), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1580(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1581(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1582(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1275(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1276(.a(gate160inter0), .b(s_104), .O(gate160inter1));
  and2  gate1277(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1278(.a(s_104), .O(gate160inter3));
  inv1  gate1279(.a(s_105), .O(gate160inter4));
  nand2 gate1280(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1281(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1282(.a(G447), .O(gate160inter7));
  inv1  gate1283(.a(G531), .O(gate160inter8));
  nand2 gate1284(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1285(.a(s_105), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1286(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1287(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1288(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate981(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate982(.a(gate174inter0), .b(s_62), .O(gate174inter1));
  and2  gate983(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate984(.a(s_62), .O(gate174inter3));
  inv1  gate985(.a(s_63), .O(gate174inter4));
  nand2 gate986(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate987(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate988(.a(G489), .O(gate174inter7));
  inv1  gate989(.a(G552), .O(gate174inter8));
  nand2 gate990(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate991(.a(s_63), .b(gate174inter3), .O(gate174inter10));
  nor2  gate992(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate993(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate994(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1513(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1514(.a(gate181inter0), .b(s_138), .O(gate181inter1));
  and2  gate1515(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1516(.a(s_138), .O(gate181inter3));
  inv1  gate1517(.a(s_139), .O(gate181inter4));
  nand2 gate1518(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1519(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1520(.a(G510), .O(gate181inter7));
  inv1  gate1521(.a(G564), .O(gate181inter8));
  nand2 gate1522(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1523(.a(s_139), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1524(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1525(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1526(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate967(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate968(.a(gate183inter0), .b(s_60), .O(gate183inter1));
  and2  gate969(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate970(.a(s_60), .O(gate183inter3));
  inv1  gate971(.a(s_61), .O(gate183inter4));
  nand2 gate972(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate973(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate974(.a(G516), .O(gate183inter7));
  inv1  gate975(.a(G567), .O(gate183inter8));
  nand2 gate976(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate977(.a(s_61), .b(gate183inter3), .O(gate183inter10));
  nor2  gate978(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate979(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate980(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1499(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1500(.a(gate184inter0), .b(s_136), .O(gate184inter1));
  and2  gate1501(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1502(.a(s_136), .O(gate184inter3));
  inv1  gate1503(.a(s_137), .O(gate184inter4));
  nand2 gate1504(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1505(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1506(.a(G519), .O(gate184inter7));
  inv1  gate1507(.a(G567), .O(gate184inter8));
  nand2 gate1508(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1509(.a(s_137), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1510(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1511(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1512(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1093(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1094(.a(gate186inter0), .b(s_78), .O(gate186inter1));
  and2  gate1095(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1096(.a(s_78), .O(gate186inter3));
  inv1  gate1097(.a(s_79), .O(gate186inter4));
  nand2 gate1098(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1099(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1100(.a(G572), .O(gate186inter7));
  inv1  gate1101(.a(G573), .O(gate186inter8));
  nand2 gate1102(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1103(.a(s_79), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1104(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1105(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1106(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1079(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1080(.a(gate190inter0), .b(s_76), .O(gate190inter1));
  and2  gate1081(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1082(.a(s_76), .O(gate190inter3));
  inv1  gate1083(.a(s_77), .O(gate190inter4));
  nand2 gate1084(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1085(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1086(.a(G580), .O(gate190inter7));
  inv1  gate1087(.a(G581), .O(gate190inter8));
  nand2 gate1088(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1089(.a(s_77), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1090(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1091(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1092(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1037(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1038(.a(gate197inter0), .b(s_70), .O(gate197inter1));
  and2  gate1039(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1040(.a(s_70), .O(gate197inter3));
  inv1  gate1041(.a(s_71), .O(gate197inter4));
  nand2 gate1042(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1043(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1044(.a(G594), .O(gate197inter7));
  inv1  gate1045(.a(G595), .O(gate197inter8));
  nand2 gate1046(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1047(.a(s_71), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1048(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1049(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1050(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate729(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate730(.a(gate201inter0), .b(s_26), .O(gate201inter1));
  and2  gate731(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate732(.a(s_26), .O(gate201inter3));
  inv1  gate733(.a(s_27), .O(gate201inter4));
  nand2 gate734(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate735(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate736(.a(G602), .O(gate201inter7));
  inv1  gate737(.a(G607), .O(gate201inter8));
  nand2 gate738(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate739(.a(s_27), .b(gate201inter3), .O(gate201inter10));
  nor2  gate740(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate741(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate742(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate589(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate590(.a(gate202inter0), .b(s_6), .O(gate202inter1));
  and2  gate591(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate592(.a(s_6), .O(gate202inter3));
  inv1  gate593(.a(s_7), .O(gate202inter4));
  nand2 gate594(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate595(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate596(.a(G612), .O(gate202inter7));
  inv1  gate597(.a(G617), .O(gate202inter8));
  nand2 gate598(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate599(.a(s_7), .b(gate202inter3), .O(gate202inter10));
  nor2  gate600(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate601(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate602(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1121(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1122(.a(gate213inter0), .b(s_82), .O(gate213inter1));
  and2  gate1123(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1124(.a(s_82), .O(gate213inter3));
  inv1  gate1125(.a(s_83), .O(gate213inter4));
  nand2 gate1126(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1127(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1128(.a(G602), .O(gate213inter7));
  inv1  gate1129(.a(G672), .O(gate213inter8));
  nand2 gate1130(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1131(.a(s_83), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1132(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1133(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1134(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate659(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate660(.a(gate216inter0), .b(s_16), .O(gate216inter1));
  and2  gate661(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate662(.a(s_16), .O(gate216inter3));
  inv1  gate663(.a(s_17), .O(gate216inter4));
  nand2 gate664(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate665(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate666(.a(G617), .O(gate216inter7));
  inv1  gate667(.a(G675), .O(gate216inter8));
  nand2 gate668(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate669(.a(s_17), .b(gate216inter3), .O(gate216inter10));
  nor2  gate670(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate671(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate672(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1541(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1542(.a(gate219inter0), .b(s_142), .O(gate219inter1));
  and2  gate1543(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1544(.a(s_142), .O(gate219inter3));
  inv1  gate1545(.a(s_143), .O(gate219inter4));
  nand2 gate1546(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1547(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1548(.a(G632), .O(gate219inter7));
  inv1  gate1549(.a(G681), .O(gate219inter8));
  nand2 gate1550(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1551(.a(s_143), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1552(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1553(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1554(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1373(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1374(.a(gate220inter0), .b(s_118), .O(gate220inter1));
  and2  gate1375(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1376(.a(s_118), .O(gate220inter3));
  inv1  gate1377(.a(s_119), .O(gate220inter4));
  nand2 gate1378(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1379(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1380(.a(G637), .O(gate220inter7));
  inv1  gate1381(.a(G681), .O(gate220inter8));
  nand2 gate1382(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1383(.a(s_119), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1384(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1385(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1386(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate799(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate800(.a(gate226inter0), .b(s_36), .O(gate226inter1));
  and2  gate801(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate802(.a(s_36), .O(gate226inter3));
  inv1  gate803(.a(s_37), .O(gate226inter4));
  nand2 gate804(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate805(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate806(.a(G692), .O(gate226inter7));
  inv1  gate807(.a(G693), .O(gate226inter8));
  nand2 gate808(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate809(.a(s_37), .b(gate226inter3), .O(gate226inter10));
  nor2  gate810(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate811(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate812(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate785(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate786(.a(gate231inter0), .b(s_34), .O(gate231inter1));
  and2  gate787(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate788(.a(s_34), .O(gate231inter3));
  inv1  gate789(.a(s_35), .O(gate231inter4));
  nand2 gate790(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate791(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate792(.a(G702), .O(gate231inter7));
  inv1  gate793(.a(G703), .O(gate231inter8));
  nand2 gate794(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate795(.a(s_35), .b(gate231inter3), .O(gate231inter10));
  nor2  gate796(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate797(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate798(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate701(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate702(.a(gate240inter0), .b(s_22), .O(gate240inter1));
  and2  gate703(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate704(.a(s_22), .O(gate240inter3));
  inv1  gate705(.a(s_23), .O(gate240inter4));
  nand2 gate706(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate707(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate708(.a(G263), .O(gate240inter7));
  inv1  gate709(.a(G715), .O(gate240inter8));
  nand2 gate710(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate711(.a(s_23), .b(gate240inter3), .O(gate240inter10));
  nor2  gate712(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate713(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate714(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate953(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate954(.a(gate249inter0), .b(s_58), .O(gate249inter1));
  and2  gate955(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate956(.a(s_58), .O(gate249inter3));
  inv1  gate957(.a(s_59), .O(gate249inter4));
  nand2 gate958(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate959(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate960(.a(G254), .O(gate249inter7));
  inv1  gate961(.a(G742), .O(gate249inter8));
  nand2 gate962(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate963(.a(s_59), .b(gate249inter3), .O(gate249inter10));
  nor2  gate964(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate965(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate966(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1205(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1206(.a(gate261inter0), .b(s_94), .O(gate261inter1));
  and2  gate1207(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1208(.a(s_94), .O(gate261inter3));
  inv1  gate1209(.a(s_95), .O(gate261inter4));
  nand2 gate1210(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1211(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1212(.a(G762), .O(gate261inter7));
  inv1  gate1213(.a(G763), .O(gate261inter8));
  nand2 gate1214(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1215(.a(s_95), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1216(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1217(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1218(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1345(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1346(.a(gate264inter0), .b(s_114), .O(gate264inter1));
  and2  gate1347(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1348(.a(s_114), .O(gate264inter3));
  inv1  gate1349(.a(s_115), .O(gate264inter4));
  nand2 gate1350(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1351(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1352(.a(G768), .O(gate264inter7));
  inv1  gate1353(.a(G769), .O(gate264inter8));
  nand2 gate1354(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1355(.a(s_115), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1356(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1357(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1358(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate687(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate688(.a(gate265inter0), .b(s_20), .O(gate265inter1));
  and2  gate689(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate690(.a(s_20), .O(gate265inter3));
  inv1  gate691(.a(s_21), .O(gate265inter4));
  nand2 gate692(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate693(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate694(.a(G642), .O(gate265inter7));
  inv1  gate695(.a(G770), .O(gate265inter8));
  nand2 gate696(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate697(.a(s_21), .b(gate265inter3), .O(gate265inter10));
  nor2  gate698(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate699(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate700(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1219(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1220(.a(gate269inter0), .b(s_96), .O(gate269inter1));
  and2  gate1221(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1222(.a(s_96), .O(gate269inter3));
  inv1  gate1223(.a(s_97), .O(gate269inter4));
  nand2 gate1224(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1225(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1226(.a(G654), .O(gate269inter7));
  inv1  gate1227(.a(G782), .O(gate269inter8));
  nand2 gate1228(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1229(.a(s_97), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1230(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1231(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1232(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1667(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1668(.a(gate276inter0), .b(s_160), .O(gate276inter1));
  and2  gate1669(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1670(.a(s_160), .O(gate276inter3));
  inv1  gate1671(.a(s_161), .O(gate276inter4));
  nand2 gate1672(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1673(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1674(.a(G773), .O(gate276inter7));
  inv1  gate1675(.a(G797), .O(gate276inter8));
  nand2 gate1676(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1677(.a(s_161), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1678(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1679(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1680(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1387(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1388(.a(gate281inter0), .b(s_120), .O(gate281inter1));
  and2  gate1389(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1390(.a(s_120), .O(gate281inter3));
  inv1  gate1391(.a(s_121), .O(gate281inter4));
  nand2 gate1392(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1393(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1394(.a(G654), .O(gate281inter7));
  inv1  gate1395(.a(G806), .O(gate281inter8));
  nand2 gate1396(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1397(.a(s_121), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1398(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1399(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1400(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1527(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1528(.a(gate289inter0), .b(s_140), .O(gate289inter1));
  and2  gate1529(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1530(.a(s_140), .O(gate289inter3));
  inv1  gate1531(.a(s_141), .O(gate289inter4));
  nand2 gate1532(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1533(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1534(.a(G818), .O(gate289inter7));
  inv1  gate1535(.a(G819), .O(gate289inter8));
  nand2 gate1536(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1537(.a(s_141), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1538(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1539(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1540(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate855(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate856(.a(gate292inter0), .b(s_44), .O(gate292inter1));
  and2  gate857(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate858(.a(s_44), .O(gate292inter3));
  inv1  gate859(.a(s_45), .O(gate292inter4));
  nand2 gate860(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate861(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate862(.a(G824), .O(gate292inter7));
  inv1  gate863(.a(G825), .O(gate292inter8));
  nand2 gate864(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate865(.a(s_45), .b(gate292inter3), .O(gate292inter10));
  nor2  gate866(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate867(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate868(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1149(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1150(.a(gate293inter0), .b(s_86), .O(gate293inter1));
  and2  gate1151(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1152(.a(s_86), .O(gate293inter3));
  inv1  gate1153(.a(s_87), .O(gate293inter4));
  nand2 gate1154(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1155(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1156(.a(G828), .O(gate293inter7));
  inv1  gate1157(.a(G829), .O(gate293inter8));
  nand2 gate1158(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1159(.a(s_87), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1160(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1161(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1162(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1401(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1402(.a(gate387inter0), .b(s_122), .O(gate387inter1));
  and2  gate1403(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1404(.a(s_122), .O(gate387inter3));
  inv1  gate1405(.a(s_123), .O(gate387inter4));
  nand2 gate1406(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1407(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1408(.a(G1), .O(gate387inter7));
  inv1  gate1409(.a(G1036), .O(gate387inter8));
  nand2 gate1410(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1411(.a(s_123), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1412(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1413(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1414(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate897(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate898(.a(gate390inter0), .b(s_50), .O(gate390inter1));
  and2  gate899(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate900(.a(s_50), .O(gate390inter3));
  inv1  gate901(.a(s_51), .O(gate390inter4));
  nand2 gate902(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate903(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate904(.a(G4), .O(gate390inter7));
  inv1  gate905(.a(G1045), .O(gate390inter8));
  nand2 gate906(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate907(.a(s_51), .b(gate390inter3), .O(gate390inter10));
  nor2  gate908(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate909(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate910(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1023(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1024(.a(gate392inter0), .b(s_68), .O(gate392inter1));
  and2  gate1025(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1026(.a(s_68), .O(gate392inter3));
  inv1  gate1027(.a(s_69), .O(gate392inter4));
  nand2 gate1028(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1029(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1030(.a(G6), .O(gate392inter7));
  inv1  gate1031(.a(G1051), .O(gate392inter8));
  nand2 gate1032(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1033(.a(s_69), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1034(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1035(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1036(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1261(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1262(.a(gate403inter0), .b(s_102), .O(gate403inter1));
  and2  gate1263(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1264(.a(s_102), .O(gate403inter3));
  inv1  gate1265(.a(s_103), .O(gate403inter4));
  nand2 gate1266(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1267(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1268(.a(G17), .O(gate403inter7));
  inv1  gate1269(.a(G1084), .O(gate403inter8));
  nand2 gate1270(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1271(.a(s_103), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1272(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1273(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1274(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1583(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1584(.a(gate407inter0), .b(s_148), .O(gate407inter1));
  and2  gate1585(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1586(.a(s_148), .O(gate407inter3));
  inv1  gate1587(.a(s_149), .O(gate407inter4));
  nand2 gate1588(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1589(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1590(.a(G21), .O(gate407inter7));
  inv1  gate1591(.a(G1096), .O(gate407inter8));
  nand2 gate1592(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1593(.a(s_149), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1594(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1595(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1596(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate715(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate716(.a(gate408inter0), .b(s_24), .O(gate408inter1));
  and2  gate717(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate718(.a(s_24), .O(gate408inter3));
  inv1  gate719(.a(s_25), .O(gate408inter4));
  nand2 gate720(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate721(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate722(.a(G22), .O(gate408inter7));
  inv1  gate723(.a(G1099), .O(gate408inter8));
  nand2 gate724(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate725(.a(s_25), .b(gate408inter3), .O(gate408inter10));
  nor2  gate726(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate727(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate728(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate547(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate548(.a(gate413inter0), .b(s_0), .O(gate413inter1));
  and2  gate549(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate550(.a(s_0), .O(gate413inter3));
  inv1  gate551(.a(s_1), .O(gate413inter4));
  nand2 gate552(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate553(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate554(.a(G27), .O(gate413inter7));
  inv1  gate555(.a(G1114), .O(gate413inter8));
  nand2 gate556(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate557(.a(s_1), .b(gate413inter3), .O(gate413inter10));
  nor2  gate558(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate559(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate560(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1359(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1360(.a(gate416inter0), .b(s_116), .O(gate416inter1));
  and2  gate1361(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1362(.a(s_116), .O(gate416inter3));
  inv1  gate1363(.a(s_117), .O(gate416inter4));
  nand2 gate1364(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1365(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1366(.a(G30), .O(gate416inter7));
  inv1  gate1367(.a(G1123), .O(gate416inter8));
  nand2 gate1368(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1369(.a(s_117), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1370(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1371(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1372(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate617(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate618(.a(gate418inter0), .b(s_10), .O(gate418inter1));
  and2  gate619(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate620(.a(s_10), .O(gate418inter3));
  inv1  gate621(.a(s_11), .O(gate418inter4));
  nand2 gate622(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate623(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate624(.a(G32), .O(gate418inter7));
  inv1  gate625(.a(G1129), .O(gate418inter8));
  nand2 gate626(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate627(.a(s_11), .b(gate418inter3), .O(gate418inter10));
  nor2  gate628(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate629(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate630(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate757(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate758(.a(gate430inter0), .b(s_30), .O(gate430inter1));
  and2  gate759(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate760(.a(s_30), .O(gate430inter3));
  inv1  gate761(.a(s_31), .O(gate430inter4));
  nand2 gate762(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate763(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate764(.a(G1051), .O(gate430inter7));
  inv1  gate765(.a(G1147), .O(gate430inter8));
  nand2 gate766(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate767(.a(s_31), .b(gate430inter3), .O(gate430inter10));
  nor2  gate768(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate769(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate770(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate925(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate926(.a(gate436inter0), .b(s_54), .O(gate436inter1));
  and2  gate927(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate928(.a(s_54), .O(gate436inter3));
  inv1  gate929(.a(s_55), .O(gate436inter4));
  nand2 gate930(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate931(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate932(.a(G1060), .O(gate436inter7));
  inv1  gate933(.a(G1156), .O(gate436inter8));
  nand2 gate934(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate935(.a(s_55), .b(gate436inter3), .O(gate436inter10));
  nor2  gate936(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate937(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate938(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1065(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1066(.a(gate439inter0), .b(s_74), .O(gate439inter1));
  and2  gate1067(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1068(.a(s_74), .O(gate439inter3));
  inv1  gate1069(.a(s_75), .O(gate439inter4));
  nand2 gate1070(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1071(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1072(.a(G11), .O(gate439inter7));
  inv1  gate1073(.a(G1162), .O(gate439inter8));
  nand2 gate1074(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1075(.a(s_75), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1076(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1077(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1078(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1443(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1444(.a(gate441inter0), .b(s_128), .O(gate441inter1));
  and2  gate1445(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1446(.a(s_128), .O(gate441inter3));
  inv1  gate1447(.a(s_129), .O(gate441inter4));
  nand2 gate1448(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1449(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1450(.a(G12), .O(gate441inter7));
  inv1  gate1451(.a(G1165), .O(gate441inter8));
  nand2 gate1452(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1453(.a(s_129), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1454(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1455(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1456(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate813(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate814(.a(gate447inter0), .b(s_38), .O(gate447inter1));
  and2  gate815(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate816(.a(s_38), .O(gate447inter3));
  inv1  gate817(.a(s_39), .O(gate447inter4));
  nand2 gate818(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate819(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate820(.a(G15), .O(gate447inter7));
  inv1  gate821(.a(G1174), .O(gate447inter8));
  nand2 gate822(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate823(.a(s_39), .b(gate447inter3), .O(gate447inter10));
  nor2  gate824(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate825(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate826(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate939(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate940(.a(gate456inter0), .b(s_56), .O(gate456inter1));
  and2  gate941(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate942(.a(s_56), .O(gate456inter3));
  inv1  gate943(.a(s_57), .O(gate456inter4));
  nand2 gate944(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate945(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate946(.a(G1090), .O(gate456inter7));
  inv1  gate947(.a(G1186), .O(gate456inter8));
  nand2 gate948(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate949(.a(s_57), .b(gate456inter3), .O(gate456inter10));
  nor2  gate950(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate951(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate952(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate869(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate870(.a(gate459inter0), .b(s_46), .O(gate459inter1));
  and2  gate871(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate872(.a(s_46), .O(gate459inter3));
  inv1  gate873(.a(s_47), .O(gate459inter4));
  nand2 gate874(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate875(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate876(.a(G21), .O(gate459inter7));
  inv1  gate877(.a(G1192), .O(gate459inter8));
  nand2 gate878(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate879(.a(s_47), .b(gate459inter3), .O(gate459inter10));
  nor2  gate880(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate881(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate882(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1289(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1290(.a(gate474inter0), .b(s_106), .O(gate474inter1));
  and2  gate1291(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1292(.a(s_106), .O(gate474inter3));
  inv1  gate1293(.a(s_107), .O(gate474inter4));
  nand2 gate1294(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1295(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1296(.a(G1117), .O(gate474inter7));
  inv1  gate1297(.a(G1213), .O(gate474inter8));
  nand2 gate1298(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1299(.a(s_107), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1300(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1301(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1302(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1331(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1332(.a(gate490inter0), .b(s_112), .O(gate490inter1));
  and2  gate1333(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1334(.a(s_112), .O(gate490inter3));
  inv1  gate1335(.a(s_113), .O(gate490inter4));
  nand2 gate1336(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1337(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1338(.a(G1242), .O(gate490inter7));
  inv1  gate1339(.a(G1243), .O(gate490inter8));
  nand2 gate1340(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1341(.a(s_113), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1342(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1343(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1344(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1653(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1654(.a(gate501inter0), .b(s_158), .O(gate501inter1));
  and2  gate1655(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1656(.a(s_158), .O(gate501inter3));
  inv1  gate1657(.a(s_159), .O(gate501inter4));
  nand2 gate1658(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1659(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1660(.a(G1264), .O(gate501inter7));
  inv1  gate1661(.a(G1265), .O(gate501inter8));
  nand2 gate1662(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1663(.a(s_159), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1664(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1665(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1666(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate771(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate772(.a(gate503inter0), .b(s_32), .O(gate503inter1));
  and2  gate773(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate774(.a(s_32), .O(gate503inter3));
  inv1  gate775(.a(s_33), .O(gate503inter4));
  nand2 gate776(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate777(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate778(.a(G1268), .O(gate503inter7));
  inv1  gate779(.a(G1269), .O(gate503inter8));
  nand2 gate780(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate781(.a(s_33), .b(gate503inter3), .O(gate503inter10));
  nor2  gate782(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate783(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate784(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1625(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1626(.a(gate509inter0), .b(s_154), .O(gate509inter1));
  and2  gate1627(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1628(.a(s_154), .O(gate509inter3));
  inv1  gate1629(.a(s_155), .O(gate509inter4));
  nand2 gate1630(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1631(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1632(.a(G1280), .O(gate509inter7));
  inv1  gate1633(.a(G1281), .O(gate509inter8));
  nand2 gate1634(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1635(.a(s_155), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1636(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1637(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1638(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate603(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate604(.a(gate513inter0), .b(s_8), .O(gate513inter1));
  and2  gate605(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate606(.a(s_8), .O(gate513inter3));
  inv1  gate607(.a(s_9), .O(gate513inter4));
  nand2 gate608(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate609(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate610(.a(G1288), .O(gate513inter7));
  inv1  gate611(.a(G1289), .O(gate513inter8));
  nand2 gate612(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate613(.a(s_9), .b(gate513inter3), .O(gate513inter10));
  nor2  gate614(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate615(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate616(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule