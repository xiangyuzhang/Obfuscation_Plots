module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1359(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1360(.a(gate17inter0), .b(s_116), .O(gate17inter1));
  and2  gate1361(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1362(.a(s_116), .O(gate17inter3));
  inv1  gate1363(.a(s_117), .O(gate17inter4));
  nand2 gate1364(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1365(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1366(.a(G17), .O(gate17inter7));
  inv1  gate1367(.a(G18), .O(gate17inter8));
  nand2 gate1368(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1369(.a(s_117), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1370(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1371(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1372(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1009(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1010(.a(gate21inter0), .b(s_66), .O(gate21inter1));
  and2  gate1011(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1012(.a(s_66), .O(gate21inter3));
  inv1  gate1013(.a(s_67), .O(gate21inter4));
  nand2 gate1014(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1015(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1016(.a(G25), .O(gate21inter7));
  inv1  gate1017(.a(G26), .O(gate21inter8));
  nand2 gate1018(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1019(.a(s_67), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1020(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1021(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1022(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1219(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1220(.a(gate23inter0), .b(s_96), .O(gate23inter1));
  and2  gate1221(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1222(.a(s_96), .O(gate23inter3));
  inv1  gate1223(.a(s_97), .O(gate23inter4));
  nand2 gate1224(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1225(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1226(.a(G29), .O(gate23inter7));
  inv1  gate1227(.a(G30), .O(gate23inter8));
  nand2 gate1228(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1229(.a(s_97), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1230(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1231(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1232(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate757(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate758(.a(gate28inter0), .b(s_30), .O(gate28inter1));
  and2  gate759(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate760(.a(s_30), .O(gate28inter3));
  inv1  gate761(.a(s_31), .O(gate28inter4));
  nand2 gate762(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate763(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate764(.a(G10), .O(gate28inter7));
  inv1  gate765(.a(G14), .O(gate28inter8));
  nand2 gate766(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate767(.a(s_31), .b(gate28inter3), .O(gate28inter10));
  nor2  gate768(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate769(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate770(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate869(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate870(.a(gate31inter0), .b(s_46), .O(gate31inter1));
  and2  gate871(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate872(.a(s_46), .O(gate31inter3));
  inv1  gate873(.a(s_47), .O(gate31inter4));
  nand2 gate874(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate875(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate876(.a(G4), .O(gate31inter7));
  inv1  gate877(.a(G8), .O(gate31inter8));
  nand2 gate878(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate879(.a(s_47), .b(gate31inter3), .O(gate31inter10));
  nor2  gate880(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate881(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate882(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate841(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate842(.a(gate44inter0), .b(s_42), .O(gate44inter1));
  and2  gate843(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate844(.a(s_42), .O(gate44inter3));
  inv1  gate845(.a(s_43), .O(gate44inter4));
  nand2 gate846(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate847(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate848(.a(G4), .O(gate44inter7));
  inv1  gate849(.a(G269), .O(gate44inter8));
  nand2 gate850(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate851(.a(s_43), .b(gate44inter3), .O(gate44inter10));
  nor2  gate852(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate853(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate854(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate687(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate688(.a(gate59inter0), .b(s_20), .O(gate59inter1));
  and2  gate689(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate690(.a(s_20), .O(gate59inter3));
  inv1  gate691(.a(s_21), .O(gate59inter4));
  nand2 gate692(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate693(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate694(.a(G19), .O(gate59inter7));
  inv1  gate695(.a(G293), .O(gate59inter8));
  nand2 gate696(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate697(.a(s_21), .b(gate59inter3), .O(gate59inter10));
  nor2  gate698(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate699(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate700(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1135(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1136(.a(gate66inter0), .b(s_84), .O(gate66inter1));
  and2  gate1137(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1138(.a(s_84), .O(gate66inter3));
  inv1  gate1139(.a(s_85), .O(gate66inter4));
  nand2 gate1140(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1141(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1142(.a(G26), .O(gate66inter7));
  inv1  gate1143(.a(G302), .O(gate66inter8));
  nand2 gate1144(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1145(.a(s_85), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1146(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1147(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1148(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1401(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1402(.a(gate71inter0), .b(s_122), .O(gate71inter1));
  and2  gate1403(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1404(.a(s_122), .O(gate71inter3));
  inv1  gate1405(.a(s_123), .O(gate71inter4));
  nand2 gate1406(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1407(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1408(.a(G31), .O(gate71inter7));
  inv1  gate1409(.a(G311), .O(gate71inter8));
  nand2 gate1410(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1411(.a(s_123), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1412(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1413(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1414(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate855(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate856(.a(gate82inter0), .b(s_44), .O(gate82inter1));
  and2  gate857(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate858(.a(s_44), .O(gate82inter3));
  inv1  gate859(.a(s_45), .O(gate82inter4));
  nand2 gate860(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate861(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate862(.a(G7), .O(gate82inter7));
  inv1  gate863(.a(G326), .O(gate82inter8));
  nand2 gate864(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate865(.a(s_45), .b(gate82inter3), .O(gate82inter10));
  nor2  gate866(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate867(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate868(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate729(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate730(.a(gate95inter0), .b(s_26), .O(gate95inter1));
  and2  gate731(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate732(.a(s_26), .O(gate95inter3));
  inv1  gate733(.a(s_27), .O(gate95inter4));
  nand2 gate734(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate735(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate736(.a(G26), .O(gate95inter7));
  inv1  gate737(.a(G347), .O(gate95inter8));
  nand2 gate738(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate739(.a(s_27), .b(gate95inter3), .O(gate95inter10));
  nor2  gate740(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate741(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate742(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate645(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate646(.a(gate100inter0), .b(s_14), .O(gate100inter1));
  and2  gate647(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate648(.a(s_14), .O(gate100inter3));
  inv1  gate649(.a(s_15), .O(gate100inter4));
  nand2 gate650(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate651(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate652(.a(G31), .O(gate100inter7));
  inv1  gate653(.a(G353), .O(gate100inter8));
  nand2 gate654(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate655(.a(s_15), .b(gate100inter3), .O(gate100inter10));
  nor2  gate656(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate657(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate658(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1317(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1318(.a(gate105inter0), .b(s_110), .O(gate105inter1));
  and2  gate1319(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1320(.a(s_110), .O(gate105inter3));
  inv1  gate1321(.a(s_111), .O(gate105inter4));
  nand2 gate1322(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1323(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1324(.a(G362), .O(gate105inter7));
  inv1  gate1325(.a(G363), .O(gate105inter8));
  nand2 gate1326(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1327(.a(s_111), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1328(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1329(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1330(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1429(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1430(.a(gate107inter0), .b(s_126), .O(gate107inter1));
  and2  gate1431(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1432(.a(s_126), .O(gate107inter3));
  inv1  gate1433(.a(s_127), .O(gate107inter4));
  nand2 gate1434(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1435(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1436(.a(G366), .O(gate107inter7));
  inv1  gate1437(.a(G367), .O(gate107inter8));
  nand2 gate1438(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1439(.a(s_127), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1440(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1441(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1442(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate659(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate660(.a(gate112inter0), .b(s_16), .O(gate112inter1));
  and2  gate661(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate662(.a(s_16), .O(gate112inter3));
  inv1  gate663(.a(s_17), .O(gate112inter4));
  nand2 gate664(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate665(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate666(.a(G376), .O(gate112inter7));
  inv1  gate667(.a(G377), .O(gate112inter8));
  nand2 gate668(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate669(.a(s_17), .b(gate112inter3), .O(gate112inter10));
  nor2  gate670(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate671(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate672(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1233(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1234(.a(gate127inter0), .b(s_98), .O(gate127inter1));
  and2  gate1235(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1236(.a(s_98), .O(gate127inter3));
  inv1  gate1237(.a(s_99), .O(gate127inter4));
  nand2 gate1238(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1239(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1240(.a(G406), .O(gate127inter7));
  inv1  gate1241(.a(G407), .O(gate127inter8));
  nand2 gate1242(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1243(.a(s_99), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1244(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1245(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1246(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate561(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate562(.a(gate130inter0), .b(s_2), .O(gate130inter1));
  and2  gate563(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate564(.a(s_2), .O(gate130inter3));
  inv1  gate565(.a(s_3), .O(gate130inter4));
  nand2 gate566(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate567(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate568(.a(G412), .O(gate130inter7));
  inv1  gate569(.a(G413), .O(gate130inter8));
  nand2 gate570(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate571(.a(s_3), .b(gate130inter3), .O(gate130inter10));
  nor2  gate572(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate573(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate574(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1261(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1262(.a(gate138inter0), .b(s_102), .O(gate138inter1));
  and2  gate1263(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1264(.a(s_102), .O(gate138inter3));
  inv1  gate1265(.a(s_103), .O(gate138inter4));
  nand2 gate1266(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1267(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1268(.a(G432), .O(gate138inter7));
  inv1  gate1269(.a(G435), .O(gate138inter8));
  nand2 gate1270(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1271(.a(s_103), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1272(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1273(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1274(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1177(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1178(.a(gate148inter0), .b(s_90), .O(gate148inter1));
  and2  gate1179(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1180(.a(s_90), .O(gate148inter3));
  inv1  gate1181(.a(s_91), .O(gate148inter4));
  nand2 gate1182(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1183(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1184(.a(G492), .O(gate148inter7));
  inv1  gate1185(.a(G495), .O(gate148inter8));
  nand2 gate1186(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1187(.a(s_91), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1188(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1189(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1190(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1275(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1276(.a(gate151inter0), .b(s_104), .O(gate151inter1));
  and2  gate1277(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1278(.a(s_104), .O(gate151inter3));
  inv1  gate1279(.a(s_105), .O(gate151inter4));
  nand2 gate1280(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1281(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1282(.a(G510), .O(gate151inter7));
  inv1  gate1283(.a(G513), .O(gate151inter8));
  nand2 gate1284(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1285(.a(s_105), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1286(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1287(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1288(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate771(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate772(.a(gate160inter0), .b(s_32), .O(gate160inter1));
  and2  gate773(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate774(.a(s_32), .O(gate160inter3));
  inv1  gate775(.a(s_33), .O(gate160inter4));
  nand2 gate776(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate777(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate778(.a(G447), .O(gate160inter7));
  inv1  gate779(.a(G531), .O(gate160inter8));
  nand2 gate780(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate781(.a(s_33), .b(gate160inter3), .O(gate160inter10));
  nor2  gate782(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate783(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate784(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate995(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate996(.a(gate167inter0), .b(s_64), .O(gate167inter1));
  and2  gate997(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate998(.a(s_64), .O(gate167inter3));
  inv1  gate999(.a(s_65), .O(gate167inter4));
  nand2 gate1000(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1001(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1002(.a(G468), .O(gate167inter7));
  inv1  gate1003(.a(G543), .O(gate167inter8));
  nand2 gate1004(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1005(.a(s_65), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1006(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1007(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1008(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1023(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1024(.a(gate175inter0), .b(s_68), .O(gate175inter1));
  and2  gate1025(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1026(.a(s_68), .O(gate175inter3));
  inv1  gate1027(.a(s_69), .O(gate175inter4));
  nand2 gate1028(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1029(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1030(.a(G492), .O(gate175inter7));
  inv1  gate1031(.a(G555), .O(gate175inter8));
  nand2 gate1032(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1033(.a(s_69), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1034(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1035(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1036(.a(gate175inter12), .b(gate175inter1), .O(G592));

  xor2  gate1331(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1332(.a(gate176inter0), .b(s_112), .O(gate176inter1));
  and2  gate1333(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1334(.a(s_112), .O(gate176inter3));
  inv1  gate1335(.a(s_113), .O(gate176inter4));
  nand2 gate1336(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1337(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1338(.a(G495), .O(gate176inter7));
  inv1  gate1339(.a(G555), .O(gate176inter8));
  nand2 gate1340(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1341(.a(s_113), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1342(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1343(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1344(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate883(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate884(.a(gate181inter0), .b(s_48), .O(gate181inter1));
  and2  gate885(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate886(.a(s_48), .O(gate181inter3));
  inv1  gate887(.a(s_49), .O(gate181inter4));
  nand2 gate888(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate889(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate890(.a(G510), .O(gate181inter7));
  inv1  gate891(.a(G564), .O(gate181inter8));
  nand2 gate892(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate893(.a(s_49), .b(gate181inter3), .O(gate181inter10));
  nor2  gate894(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate895(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate896(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate953(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate954(.a(gate188inter0), .b(s_58), .O(gate188inter1));
  and2  gate955(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate956(.a(s_58), .O(gate188inter3));
  inv1  gate957(.a(s_59), .O(gate188inter4));
  nand2 gate958(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate959(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate960(.a(G576), .O(gate188inter7));
  inv1  gate961(.a(G577), .O(gate188inter8));
  nand2 gate962(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate963(.a(s_59), .b(gate188inter3), .O(gate188inter10));
  nor2  gate964(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate965(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate966(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate673(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate674(.a(gate190inter0), .b(s_18), .O(gate190inter1));
  and2  gate675(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate676(.a(s_18), .O(gate190inter3));
  inv1  gate677(.a(s_19), .O(gate190inter4));
  nand2 gate678(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate679(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate680(.a(G580), .O(gate190inter7));
  inv1  gate681(.a(G581), .O(gate190inter8));
  nand2 gate682(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate683(.a(s_19), .b(gate190inter3), .O(gate190inter10));
  nor2  gate684(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate685(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate686(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate547(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate548(.a(gate195inter0), .b(s_0), .O(gate195inter1));
  and2  gate549(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate550(.a(s_0), .O(gate195inter3));
  inv1  gate551(.a(s_1), .O(gate195inter4));
  nand2 gate552(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate553(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate554(.a(G590), .O(gate195inter7));
  inv1  gate555(.a(G591), .O(gate195inter8));
  nand2 gate556(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate557(.a(s_1), .b(gate195inter3), .O(gate195inter10));
  nor2  gate558(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate559(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate560(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1289(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1290(.a(gate196inter0), .b(s_106), .O(gate196inter1));
  and2  gate1291(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1292(.a(s_106), .O(gate196inter3));
  inv1  gate1293(.a(s_107), .O(gate196inter4));
  nand2 gate1294(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1295(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1296(.a(G592), .O(gate196inter7));
  inv1  gate1297(.a(G593), .O(gate196inter8));
  nand2 gate1298(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1299(.a(s_107), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1300(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1301(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1302(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate631(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate632(.a(gate212inter0), .b(s_12), .O(gate212inter1));
  and2  gate633(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate634(.a(s_12), .O(gate212inter3));
  inv1  gate635(.a(s_13), .O(gate212inter4));
  nand2 gate636(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate637(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate638(.a(G617), .O(gate212inter7));
  inv1  gate639(.a(G669), .O(gate212inter8));
  nand2 gate640(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate641(.a(s_13), .b(gate212inter3), .O(gate212inter10));
  nor2  gate642(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate643(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate644(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate981(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate982(.a(gate213inter0), .b(s_62), .O(gate213inter1));
  and2  gate983(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate984(.a(s_62), .O(gate213inter3));
  inv1  gate985(.a(s_63), .O(gate213inter4));
  nand2 gate986(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate987(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate988(.a(G602), .O(gate213inter7));
  inv1  gate989(.a(G672), .O(gate213inter8));
  nand2 gate990(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate991(.a(s_63), .b(gate213inter3), .O(gate213inter10));
  nor2  gate992(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate993(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate994(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1037(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1038(.a(gate218inter0), .b(s_70), .O(gate218inter1));
  and2  gate1039(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1040(.a(s_70), .O(gate218inter3));
  inv1  gate1041(.a(s_71), .O(gate218inter4));
  nand2 gate1042(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1043(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1044(.a(G627), .O(gate218inter7));
  inv1  gate1045(.a(G678), .O(gate218inter8));
  nand2 gate1046(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1047(.a(s_71), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1048(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1049(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1050(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1345(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1346(.a(gate233inter0), .b(s_114), .O(gate233inter1));
  and2  gate1347(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1348(.a(s_114), .O(gate233inter3));
  inv1  gate1349(.a(s_115), .O(gate233inter4));
  nand2 gate1350(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1351(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1352(.a(G242), .O(gate233inter7));
  inv1  gate1353(.a(G718), .O(gate233inter8));
  nand2 gate1354(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1355(.a(s_115), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1356(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1357(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1358(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1093(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1094(.a(gate234inter0), .b(s_78), .O(gate234inter1));
  and2  gate1095(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1096(.a(s_78), .O(gate234inter3));
  inv1  gate1097(.a(s_79), .O(gate234inter4));
  nand2 gate1098(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1099(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1100(.a(G245), .O(gate234inter7));
  inv1  gate1101(.a(G721), .O(gate234inter8));
  nand2 gate1102(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1103(.a(s_79), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1104(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1105(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1106(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate939(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate940(.a(gate251inter0), .b(s_56), .O(gate251inter1));
  and2  gate941(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate942(.a(s_56), .O(gate251inter3));
  inv1  gate943(.a(s_57), .O(gate251inter4));
  nand2 gate944(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate945(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate946(.a(G257), .O(gate251inter7));
  inv1  gate947(.a(G745), .O(gate251inter8));
  nand2 gate948(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate949(.a(s_57), .b(gate251inter3), .O(gate251inter10));
  nor2  gate950(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate951(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate952(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1065(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1066(.a(gate254inter0), .b(s_74), .O(gate254inter1));
  and2  gate1067(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1068(.a(s_74), .O(gate254inter3));
  inv1  gate1069(.a(s_75), .O(gate254inter4));
  nand2 gate1070(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1071(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1072(.a(G712), .O(gate254inter7));
  inv1  gate1073(.a(G748), .O(gate254inter8));
  nand2 gate1074(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1075(.a(s_75), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1076(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1077(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1078(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate911(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate912(.a(gate256inter0), .b(s_52), .O(gate256inter1));
  and2  gate913(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate914(.a(s_52), .O(gate256inter3));
  inv1  gate915(.a(s_53), .O(gate256inter4));
  nand2 gate916(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate917(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate918(.a(G715), .O(gate256inter7));
  inv1  gate919(.a(G751), .O(gate256inter8));
  nand2 gate920(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate921(.a(s_53), .b(gate256inter3), .O(gate256inter10));
  nor2  gate922(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate923(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate924(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate617(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate618(.a(gate266inter0), .b(s_10), .O(gate266inter1));
  and2  gate619(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate620(.a(s_10), .O(gate266inter3));
  inv1  gate621(.a(s_11), .O(gate266inter4));
  nand2 gate622(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate623(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate624(.a(G645), .O(gate266inter7));
  inv1  gate625(.a(G773), .O(gate266inter8));
  nand2 gate626(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate627(.a(s_11), .b(gate266inter3), .O(gate266inter10));
  nor2  gate628(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate629(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate630(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1051(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1052(.a(gate269inter0), .b(s_72), .O(gate269inter1));
  and2  gate1053(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1054(.a(s_72), .O(gate269inter3));
  inv1  gate1055(.a(s_73), .O(gate269inter4));
  nand2 gate1056(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1057(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1058(.a(G654), .O(gate269inter7));
  inv1  gate1059(.a(G782), .O(gate269inter8));
  nand2 gate1060(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1061(.a(s_73), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1062(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1063(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1064(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate925(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate926(.a(gate272inter0), .b(s_54), .O(gate272inter1));
  and2  gate927(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate928(.a(s_54), .O(gate272inter3));
  inv1  gate929(.a(s_55), .O(gate272inter4));
  nand2 gate930(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate931(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate932(.a(G663), .O(gate272inter7));
  inv1  gate933(.a(G791), .O(gate272inter8));
  nand2 gate934(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate935(.a(s_55), .b(gate272inter3), .O(gate272inter10));
  nor2  gate936(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate937(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate938(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate897(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate898(.a(gate387inter0), .b(s_50), .O(gate387inter1));
  and2  gate899(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate900(.a(s_50), .O(gate387inter3));
  inv1  gate901(.a(s_51), .O(gate387inter4));
  nand2 gate902(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate903(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate904(.a(G1), .O(gate387inter7));
  inv1  gate905(.a(G1036), .O(gate387inter8));
  nand2 gate906(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate907(.a(s_51), .b(gate387inter3), .O(gate387inter10));
  nor2  gate908(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate909(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate910(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate799(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate800(.a(gate390inter0), .b(s_36), .O(gate390inter1));
  and2  gate801(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate802(.a(s_36), .O(gate390inter3));
  inv1  gate803(.a(s_37), .O(gate390inter4));
  nand2 gate804(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate805(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate806(.a(G4), .O(gate390inter7));
  inv1  gate807(.a(G1045), .O(gate390inter8));
  nand2 gate808(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate809(.a(s_37), .b(gate390inter3), .O(gate390inter10));
  nor2  gate810(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate811(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate812(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate967(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate968(.a(gate392inter0), .b(s_60), .O(gate392inter1));
  and2  gate969(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate970(.a(s_60), .O(gate392inter3));
  inv1  gate971(.a(s_61), .O(gate392inter4));
  nand2 gate972(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate973(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate974(.a(G6), .O(gate392inter7));
  inv1  gate975(.a(G1051), .O(gate392inter8));
  nand2 gate976(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate977(.a(s_61), .b(gate392inter3), .O(gate392inter10));
  nor2  gate978(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate979(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate980(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate701(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate702(.a(gate405inter0), .b(s_22), .O(gate405inter1));
  and2  gate703(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate704(.a(s_22), .O(gate405inter3));
  inv1  gate705(.a(s_23), .O(gate405inter4));
  nand2 gate706(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate707(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate708(.a(G19), .O(gate405inter7));
  inv1  gate709(.a(G1090), .O(gate405inter8));
  nand2 gate710(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate711(.a(s_23), .b(gate405inter3), .O(gate405inter10));
  nor2  gate712(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate713(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate714(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate715(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate716(.a(gate409inter0), .b(s_24), .O(gate409inter1));
  and2  gate717(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate718(.a(s_24), .O(gate409inter3));
  inv1  gate719(.a(s_25), .O(gate409inter4));
  nand2 gate720(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate721(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate722(.a(G23), .O(gate409inter7));
  inv1  gate723(.a(G1102), .O(gate409inter8));
  nand2 gate724(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate725(.a(s_25), .b(gate409inter3), .O(gate409inter10));
  nor2  gate726(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate727(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate728(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1121(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1122(.a(gate411inter0), .b(s_82), .O(gate411inter1));
  and2  gate1123(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1124(.a(s_82), .O(gate411inter3));
  inv1  gate1125(.a(s_83), .O(gate411inter4));
  nand2 gate1126(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1127(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1128(.a(G25), .O(gate411inter7));
  inv1  gate1129(.a(G1108), .O(gate411inter8));
  nand2 gate1130(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1131(.a(s_83), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1132(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1133(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1134(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate603(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate604(.a(gate413inter0), .b(s_8), .O(gate413inter1));
  and2  gate605(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate606(.a(s_8), .O(gate413inter3));
  inv1  gate607(.a(s_9), .O(gate413inter4));
  nand2 gate608(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate609(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate610(.a(G27), .O(gate413inter7));
  inv1  gate611(.a(G1114), .O(gate413inter8));
  nand2 gate612(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate613(.a(s_9), .b(gate413inter3), .O(gate413inter10));
  nor2  gate614(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate615(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate616(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1247(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1248(.a(gate415inter0), .b(s_100), .O(gate415inter1));
  and2  gate1249(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1250(.a(s_100), .O(gate415inter3));
  inv1  gate1251(.a(s_101), .O(gate415inter4));
  nand2 gate1252(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1253(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1254(.a(G29), .O(gate415inter7));
  inv1  gate1255(.a(G1120), .O(gate415inter8));
  nand2 gate1256(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1257(.a(s_101), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1258(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1259(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1260(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate575(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate576(.a(gate416inter0), .b(s_4), .O(gate416inter1));
  and2  gate577(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate578(.a(s_4), .O(gate416inter3));
  inv1  gate579(.a(s_5), .O(gate416inter4));
  nand2 gate580(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate581(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate582(.a(G30), .O(gate416inter7));
  inv1  gate583(.a(G1123), .O(gate416inter8));
  nand2 gate584(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate585(.a(s_5), .b(gate416inter3), .O(gate416inter10));
  nor2  gate586(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate587(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate588(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1079(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1080(.a(gate425inter0), .b(s_76), .O(gate425inter1));
  and2  gate1081(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1082(.a(s_76), .O(gate425inter3));
  inv1  gate1083(.a(s_77), .O(gate425inter4));
  nand2 gate1084(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1085(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1086(.a(G4), .O(gate425inter7));
  inv1  gate1087(.a(G1141), .O(gate425inter8));
  nand2 gate1088(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1089(.a(s_77), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1090(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1091(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1092(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate813(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate814(.a(gate433inter0), .b(s_38), .O(gate433inter1));
  and2  gate815(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate816(.a(s_38), .O(gate433inter3));
  inv1  gate817(.a(s_39), .O(gate433inter4));
  nand2 gate818(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate819(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate820(.a(G8), .O(gate433inter7));
  inv1  gate821(.a(G1153), .O(gate433inter8));
  nand2 gate822(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate823(.a(s_39), .b(gate433inter3), .O(gate433inter10));
  nor2  gate824(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate825(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate826(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate785(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate786(.a(gate445inter0), .b(s_34), .O(gate445inter1));
  and2  gate787(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate788(.a(s_34), .O(gate445inter3));
  inv1  gate789(.a(s_35), .O(gate445inter4));
  nand2 gate790(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate791(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate792(.a(G14), .O(gate445inter7));
  inv1  gate793(.a(G1171), .O(gate445inter8));
  nand2 gate794(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate795(.a(s_35), .b(gate445inter3), .O(gate445inter10));
  nor2  gate796(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate797(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate798(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1443(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1444(.a(gate452inter0), .b(s_128), .O(gate452inter1));
  and2  gate1445(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1446(.a(s_128), .O(gate452inter3));
  inv1  gate1447(.a(s_129), .O(gate452inter4));
  nand2 gate1448(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1449(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1450(.a(G1084), .O(gate452inter7));
  inv1  gate1451(.a(G1180), .O(gate452inter8));
  nand2 gate1452(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1453(.a(s_129), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1454(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1455(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1456(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1415(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1416(.a(gate466inter0), .b(s_124), .O(gate466inter1));
  and2  gate1417(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1418(.a(s_124), .O(gate466inter3));
  inv1  gate1419(.a(s_125), .O(gate466inter4));
  nand2 gate1420(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1421(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1422(.a(G1105), .O(gate466inter7));
  inv1  gate1423(.a(G1201), .O(gate466inter8));
  nand2 gate1424(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1425(.a(s_125), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1426(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1427(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1428(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1457(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1458(.a(gate468inter0), .b(s_130), .O(gate468inter1));
  and2  gate1459(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1460(.a(s_130), .O(gate468inter3));
  inv1  gate1461(.a(s_131), .O(gate468inter4));
  nand2 gate1462(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1463(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1464(.a(G1108), .O(gate468inter7));
  inv1  gate1465(.a(G1204), .O(gate468inter8));
  nand2 gate1466(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1467(.a(s_131), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1468(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1469(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1470(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1205(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1206(.a(gate476inter0), .b(s_94), .O(gate476inter1));
  and2  gate1207(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1208(.a(s_94), .O(gate476inter3));
  inv1  gate1209(.a(s_95), .O(gate476inter4));
  nand2 gate1210(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1211(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1212(.a(G1120), .O(gate476inter7));
  inv1  gate1213(.a(G1216), .O(gate476inter8));
  nand2 gate1214(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1215(.a(s_95), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1216(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1217(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1218(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1303(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1304(.a(gate480inter0), .b(s_108), .O(gate480inter1));
  and2  gate1305(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1306(.a(s_108), .O(gate480inter3));
  inv1  gate1307(.a(s_109), .O(gate480inter4));
  nand2 gate1308(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1309(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1310(.a(G1126), .O(gate480inter7));
  inv1  gate1311(.a(G1222), .O(gate480inter8));
  nand2 gate1312(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1313(.a(s_109), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1314(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1315(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1316(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1191(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1192(.a(gate481inter0), .b(s_92), .O(gate481inter1));
  and2  gate1193(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1194(.a(s_92), .O(gate481inter3));
  inv1  gate1195(.a(s_93), .O(gate481inter4));
  nand2 gate1196(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1197(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1198(.a(G32), .O(gate481inter7));
  inv1  gate1199(.a(G1225), .O(gate481inter8));
  nand2 gate1200(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1201(.a(s_93), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1202(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1203(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1204(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate827(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate828(.a(gate484inter0), .b(s_40), .O(gate484inter1));
  and2  gate829(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate830(.a(s_40), .O(gate484inter3));
  inv1  gate831(.a(s_41), .O(gate484inter4));
  nand2 gate832(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate833(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate834(.a(G1230), .O(gate484inter7));
  inv1  gate835(.a(G1231), .O(gate484inter8));
  nand2 gate836(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate837(.a(s_41), .b(gate484inter3), .O(gate484inter10));
  nor2  gate838(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate839(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate840(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1373(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1374(.a(gate490inter0), .b(s_118), .O(gate490inter1));
  and2  gate1375(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1376(.a(s_118), .O(gate490inter3));
  inv1  gate1377(.a(s_119), .O(gate490inter4));
  nand2 gate1378(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1379(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1380(.a(G1242), .O(gate490inter7));
  inv1  gate1381(.a(G1243), .O(gate490inter8));
  nand2 gate1382(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1383(.a(s_119), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1384(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1385(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1386(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1149(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1150(.a(gate491inter0), .b(s_86), .O(gate491inter1));
  and2  gate1151(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1152(.a(s_86), .O(gate491inter3));
  inv1  gate1153(.a(s_87), .O(gate491inter4));
  nand2 gate1154(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1155(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1156(.a(G1244), .O(gate491inter7));
  inv1  gate1157(.a(G1245), .O(gate491inter8));
  nand2 gate1158(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1159(.a(s_87), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1160(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1161(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1162(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1163(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1164(.a(gate496inter0), .b(s_88), .O(gate496inter1));
  and2  gate1165(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1166(.a(s_88), .O(gate496inter3));
  inv1  gate1167(.a(s_89), .O(gate496inter4));
  nand2 gate1168(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1169(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1170(.a(G1254), .O(gate496inter7));
  inv1  gate1171(.a(G1255), .O(gate496inter8));
  nand2 gate1172(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1173(.a(s_89), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1174(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1175(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1176(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate589(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate590(.a(gate497inter0), .b(s_6), .O(gate497inter1));
  and2  gate591(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate592(.a(s_6), .O(gate497inter3));
  inv1  gate593(.a(s_7), .O(gate497inter4));
  nand2 gate594(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate595(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate596(.a(G1256), .O(gate497inter7));
  inv1  gate597(.a(G1257), .O(gate497inter8));
  nand2 gate598(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate599(.a(s_7), .b(gate497inter3), .O(gate497inter10));
  nor2  gate600(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate601(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate602(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1387(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1388(.a(gate498inter0), .b(s_120), .O(gate498inter1));
  and2  gate1389(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1390(.a(s_120), .O(gate498inter3));
  inv1  gate1391(.a(s_121), .O(gate498inter4));
  nand2 gate1392(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1393(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1394(.a(G1258), .O(gate498inter7));
  inv1  gate1395(.a(G1259), .O(gate498inter8));
  nand2 gate1396(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1397(.a(s_121), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1398(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1399(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1400(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1107(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1108(.a(gate499inter0), .b(s_80), .O(gate499inter1));
  and2  gate1109(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1110(.a(s_80), .O(gate499inter3));
  inv1  gate1111(.a(s_81), .O(gate499inter4));
  nand2 gate1112(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1113(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1114(.a(G1260), .O(gate499inter7));
  inv1  gate1115(.a(G1261), .O(gate499inter8));
  nand2 gate1116(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1117(.a(s_81), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1118(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1119(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1120(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate743(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate744(.a(gate505inter0), .b(s_28), .O(gate505inter1));
  and2  gate745(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate746(.a(s_28), .O(gate505inter3));
  inv1  gate747(.a(s_29), .O(gate505inter4));
  nand2 gate748(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate749(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate750(.a(G1272), .O(gate505inter7));
  inv1  gate751(.a(G1273), .O(gate505inter8));
  nand2 gate752(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate753(.a(s_29), .b(gate505inter3), .O(gate505inter10));
  nor2  gate754(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate755(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate756(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule