module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate939(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate940(.a(gate9inter0), .b(s_56), .O(gate9inter1));
  and2  gate941(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate942(.a(s_56), .O(gate9inter3));
  inv1  gate943(.a(s_57), .O(gate9inter4));
  nand2 gate944(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate945(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate946(.a(G1), .O(gate9inter7));
  inv1  gate947(.a(G2), .O(gate9inter8));
  nand2 gate948(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate949(.a(s_57), .b(gate9inter3), .O(gate9inter10));
  nor2  gate950(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate951(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate952(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2395(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2396(.a(gate13inter0), .b(s_264), .O(gate13inter1));
  and2  gate2397(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2398(.a(s_264), .O(gate13inter3));
  inv1  gate2399(.a(s_265), .O(gate13inter4));
  nand2 gate2400(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2401(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2402(.a(G9), .O(gate13inter7));
  inv1  gate2403(.a(G10), .O(gate13inter8));
  nand2 gate2404(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2405(.a(s_265), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2406(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2407(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2408(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1107(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1108(.a(gate18inter0), .b(s_80), .O(gate18inter1));
  and2  gate1109(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1110(.a(s_80), .O(gate18inter3));
  inv1  gate1111(.a(s_81), .O(gate18inter4));
  nand2 gate1112(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1113(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1114(.a(G19), .O(gate18inter7));
  inv1  gate1115(.a(G20), .O(gate18inter8));
  nand2 gate1116(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1117(.a(s_81), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1118(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1119(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1120(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate561(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate562(.a(gate24inter0), .b(s_2), .O(gate24inter1));
  and2  gate563(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate564(.a(s_2), .O(gate24inter3));
  inv1  gate565(.a(s_3), .O(gate24inter4));
  nand2 gate566(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate567(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate568(.a(G31), .O(gate24inter7));
  inv1  gate569(.a(G32), .O(gate24inter8));
  nand2 gate570(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate571(.a(s_3), .b(gate24inter3), .O(gate24inter10));
  nor2  gate572(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate573(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate574(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate659(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate660(.a(gate28inter0), .b(s_16), .O(gate28inter1));
  and2  gate661(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate662(.a(s_16), .O(gate28inter3));
  inv1  gate663(.a(s_17), .O(gate28inter4));
  nand2 gate664(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate665(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate666(.a(G10), .O(gate28inter7));
  inv1  gate667(.a(G14), .O(gate28inter8));
  nand2 gate668(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate669(.a(s_17), .b(gate28inter3), .O(gate28inter10));
  nor2  gate670(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate671(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate672(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1961(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1962(.a(gate29inter0), .b(s_202), .O(gate29inter1));
  and2  gate1963(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1964(.a(s_202), .O(gate29inter3));
  inv1  gate1965(.a(s_203), .O(gate29inter4));
  nand2 gate1966(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1967(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1968(.a(G3), .O(gate29inter7));
  inv1  gate1969(.a(G7), .O(gate29inter8));
  nand2 gate1970(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1971(.a(s_203), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1972(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1973(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1974(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1555(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1556(.a(gate37inter0), .b(s_144), .O(gate37inter1));
  and2  gate1557(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1558(.a(s_144), .O(gate37inter3));
  inv1  gate1559(.a(s_145), .O(gate37inter4));
  nand2 gate1560(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1561(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1562(.a(G19), .O(gate37inter7));
  inv1  gate1563(.a(G23), .O(gate37inter8));
  nand2 gate1564(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1565(.a(s_145), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1566(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1567(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1568(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1513(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1514(.a(gate39inter0), .b(s_138), .O(gate39inter1));
  and2  gate1515(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1516(.a(s_138), .O(gate39inter3));
  inv1  gate1517(.a(s_139), .O(gate39inter4));
  nand2 gate1518(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1519(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1520(.a(G20), .O(gate39inter7));
  inv1  gate1521(.a(G24), .O(gate39inter8));
  nand2 gate1522(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1523(.a(s_139), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1524(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1525(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1526(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1205(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1206(.a(gate40inter0), .b(s_94), .O(gate40inter1));
  and2  gate1207(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1208(.a(s_94), .O(gate40inter3));
  inv1  gate1209(.a(s_95), .O(gate40inter4));
  nand2 gate1210(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1211(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1212(.a(G28), .O(gate40inter7));
  inv1  gate1213(.a(G32), .O(gate40inter8));
  nand2 gate1214(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1215(.a(s_95), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1216(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1217(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1218(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate743(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate744(.a(gate46inter0), .b(s_28), .O(gate46inter1));
  and2  gate745(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate746(.a(s_28), .O(gate46inter3));
  inv1  gate747(.a(s_29), .O(gate46inter4));
  nand2 gate748(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate749(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate750(.a(G6), .O(gate46inter7));
  inv1  gate751(.a(G272), .O(gate46inter8));
  nand2 gate752(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate753(.a(s_29), .b(gate46inter3), .O(gate46inter10));
  nor2  gate754(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate755(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate756(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate2339(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2340(.a(gate47inter0), .b(s_256), .O(gate47inter1));
  and2  gate2341(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2342(.a(s_256), .O(gate47inter3));
  inv1  gate2343(.a(s_257), .O(gate47inter4));
  nand2 gate2344(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2345(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2346(.a(G7), .O(gate47inter7));
  inv1  gate2347(.a(G275), .O(gate47inter8));
  nand2 gate2348(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2349(.a(s_257), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2350(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2351(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2352(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1163(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1164(.a(gate48inter0), .b(s_88), .O(gate48inter1));
  and2  gate1165(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1166(.a(s_88), .O(gate48inter3));
  inv1  gate1167(.a(s_89), .O(gate48inter4));
  nand2 gate1168(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1169(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1170(.a(G8), .O(gate48inter7));
  inv1  gate1171(.a(G275), .O(gate48inter8));
  nand2 gate1172(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1173(.a(s_89), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1174(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1175(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1176(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate2297(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2298(.a(gate53inter0), .b(s_250), .O(gate53inter1));
  and2  gate2299(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2300(.a(s_250), .O(gate53inter3));
  inv1  gate2301(.a(s_251), .O(gate53inter4));
  nand2 gate2302(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2303(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2304(.a(G13), .O(gate53inter7));
  inv1  gate2305(.a(G284), .O(gate53inter8));
  nand2 gate2306(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2307(.a(s_251), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2308(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2309(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2310(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate2115(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2116(.a(gate60inter0), .b(s_224), .O(gate60inter1));
  and2  gate2117(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2118(.a(s_224), .O(gate60inter3));
  inv1  gate2119(.a(s_225), .O(gate60inter4));
  nand2 gate2120(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2121(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2122(.a(G20), .O(gate60inter7));
  inv1  gate2123(.a(G293), .O(gate60inter8));
  nand2 gate2124(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2125(.a(s_225), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2126(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2127(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2128(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1135(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1136(.a(gate64inter0), .b(s_84), .O(gate64inter1));
  and2  gate1137(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1138(.a(s_84), .O(gate64inter3));
  inv1  gate1139(.a(s_85), .O(gate64inter4));
  nand2 gate1140(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1141(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1142(.a(G24), .O(gate64inter7));
  inv1  gate1143(.a(G299), .O(gate64inter8));
  nand2 gate1144(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1145(.a(s_85), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1146(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1147(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1148(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate575(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate576(.a(gate67inter0), .b(s_4), .O(gate67inter1));
  and2  gate577(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate578(.a(s_4), .O(gate67inter3));
  inv1  gate579(.a(s_5), .O(gate67inter4));
  nand2 gate580(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate581(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate582(.a(G27), .O(gate67inter7));
  inv1  gate583(.a(G305), .O(gate67inter8));
  nand2 gate584(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate585(.a(s_5), .b(gate67inter3), .O(gate67inter10));
  nor2  gate586(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate587(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate588(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2255(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2256(.a(gate70inter0), .b(s_244), .O(gate70inter1));
  and2  gate2257(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2258(.a(s_244), .O(gate70inter3));
  inv1  gate2259(.a(s_245), .O(gate70inter4));
  nand2 gate2260(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2261(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2262(.a(G30), .O(gate70inter7));
  inv1  gate2263(.a(G308), .O(gate70inter8));
  nand2 gate2264(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2265(.a(s_245), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2266(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2267(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2268(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate631(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate632(.a(gate75inter0), .b(s_12), .O(gate75inter1));
  and2  gate633(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate634(.a(s_12), .O(gate75inter3));
  inv1  gate635(.a(s_13), .O(gate75inter4));
  nand2 gate636(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate637(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate638(.a(G9), .O(gate75inter7));
  inv1  gate639(.a(G317), .O(gate75inter8));
  nand2 gate640(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate641(.a(s_13), .b(gate75inter3), .O(gate75inter10));
  nor2  gate642(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate643(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate644(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1401(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1402(.a(gate80inter0), .b(s_122), .O(gate80inter1));
  and2  gate1403(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1404(.a(s_122), .O(gate80inter3));
  inv1  gate1405(.a(s_123), .O(gate80inter4));
  nand2 gate1406(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1407(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1408(.a(G14), .O(gate80inter7));
  inv1  gate1409(.a(G323), .O(gate80inter8));
  nand2 gate1410(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1411(.a(s_123), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1412(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1413(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1414(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2213(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2214(.a(gate81inter0), .b(s_238), .O(gate81inter1));
  and2  gate2215(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2216(.a(s_238), .O(gate81inter3));
  inv1  gate2217(.a(s_239), .O(gate81inter4));
  nand2 gate2218(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2219(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2220(.a(G3), .O(gate81inter7));
  inv1  gate2221(.a(G326), .O(gate81inter8));
  nand2 gate2222(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2223(.a(s_239), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2224(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2225(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2226(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate2367(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2368(.a(gate83inter0), .b(s_260), .O(gate83inter1));
  and2  gate2369(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2370(.a(s_260), .O(gate83inter3));
  inv1  gate2371(.a(s_261), .O(gate83inter4));
  nand2 gate2372(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2373(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2374(.a(G11), .O(gate83inter7));
  inv1  gate2375(.a(G329), .O(gate83inter8));
  nand2 gate2376(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2377(.a(s_261), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2378(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2379(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2380(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1219(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1220(.a(gate85inter0), .b(s_96), .O(gate85inter1));
  and2  gate1221(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1222(.a(s_96), .O(gate85inter3));
  inv1  gate1223(.a(s_97), .O(gate85inter4));
  nand2 gate1224(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1225(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1226(.a(G4), .O(gate85inter7));
  inv1  gate1227(.a(G332), .O(gate85inter8));
  nand2 gate1228(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1229(.a(s_97), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1230(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1231(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1232(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1835(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1836(.a(gate88inter0), .b(s_184), .O(gate88inter1));
  and2  gate1837(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1838(.a(s_184), .O(gate88inter3));
  inv1  gate1839(.a(s_185), .O(gate88inter4));
  nand2 gate1840(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1841(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1842(.a(G16), .O(gate88inter7));
  inv1  gate1843(.a(G335), .O(gate88inter8));
  nand2 gate1844(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1845(.a(s_185), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1846(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1847(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1848(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1681(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1682(.a(gate91inter0), .b(s_162), .O(gate91inter1));
  and2  gate1683(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1684(.a(s_162), .O(gate91inter3));
  inv1  gate1685(.a(s_163), .O(gate91inter4));
  nand2 gate1686(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1687(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1688(.a(G25), .O(gate91inter7));
  inv1  gate1689(.a(G341), .O(gate91inter8));
  nand2 gate1690(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1691(.a(s_163), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1692(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1693(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1694(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate715(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate716(.a(gate100inter0), .b(s_24), .O(gate100inter1));
  and2  gate717(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate718(.a(s_24), .O(gate100inter3));
  inv1  gate719(.a(s_25), .O(gate100inter4));
  nand2 gate720(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate721(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate722(.a(G31), .O(gate100inter7));
  inv1  gate723(.a(G353), .O(gate100inter8));
  nand2 gate724(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate725(.a(s_25), .b(gate100inter3), .O(gate100inter10));
  nor2  gate726(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate727(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate728(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate701(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate702(.a(gate101inter0), .b(s_22), .O(gate101inter1));
  and2  gate703(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate704(.a(s_22), .O(gate101inter3));
  inv1  gate705(.a(s_23), .O(gate101inter4));
  nand2 gate706(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate707(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate708(.a(G20), .O(gate101inter7));
  inv1  gate709(.a(G356), .O(gate101inter8));
  nand2 gate710(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate711(.a(s_23), .b(gate101inter3), .O(gate101inter10));
  nor2  gate712(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate713(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate714(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1919(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1920(.a(gate104inter0), .b(s_196), .O(gate104inter1));
  and2  gate1921(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1922(.a(s_196), .O(gate104inter3));
  inv1  gate1923(.a(s_197), .O(gate104inter4));
  nand2 gate1924(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1925(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1926(.a(G32), .O(gate104inter7));
  inv1  gate1927(.a(G359), .O(gate104inter8));
  nand2 gate1928(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1929(.a(s_197), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1930(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1931(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1932(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate883(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate884(.a(gate105inter0), .b(s_48), .O(gate105inter1));
  and2  gate885(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate886(.a(s_48), .O(gate105inter3));
  inv1  gate887(.a(s_49), .O(gate105inter4));
  nand2 gate888(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate889(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate890(.a(G362), .O(gate105inter7));
  inv1  gate891(.a(G363), .O(gate105inter8));
  nand2 gate892(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate893(.a(s_49), .b(gate105inter3), .O(gate105inter10));
  nor2  gate894(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate895(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate896(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1191(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1192(.a(gate111inter0), .b(s_92), .O(gate111inter1));
  and2  gate1193(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1194(.a(s_92), .O(gate111inter3));
  inv1  gate1195(.a(s_93), .O(gate111inter4));
  nand2 gate1196(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1197(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1198(.a(G374), .O(gate111inter7));
  inv1  gate1199(.a(G375), .O(gate111inter8));
  nand2 gate1200(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1201(.a(s_93), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1202(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1203(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1204(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate617(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate618(.a(gate112inter0), .b(s_10), .O(gate112inter1));
  and2  gate619(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate620(.a(s_10), .O(gate112inter3));
  inv1  gate621(.a(s_11), .O(gate112inter4));
  nand2 gate622(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate623(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate624(.a(G376), .O(gate112inter7));
  inv1  gate625(.a(G377), .O(gate112inter8));
  nand2 gate626(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate627(.a(s_11), .b(gate112inter3), .O(gate112inter10));
  nor2  gate628(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate629(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate630(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate1779(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1780(.a(gate113inter0), .b(s_176), .O(gate113inter1));
  and2  gate1781(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1782(.a(s_176), .O(gate113inter3));
  inv1  gate1783(.a(s_177), .O(gate113inter4));
  nand2 gate1784(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1785(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1786(.a(G378), .O(gate113inter7));
  inv1  gate1787(.a(G379), .O(gate113inter8));
  nand2 gate1788(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1789(.a(s_177), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1790(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1791(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1792(.a(gate113inter12), .b(gate113inter1), .O(G450));

  xor2  gate799(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate800(.a(gate114inter0), .b(s_36), .O(gate114inter1));
  and2  gate801(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate802(.a(s_36), .O(gate114inter3));
  inv1  gate803(.a(s_37), .O(gate114inter4));
  nand2 gate804(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate805(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate806(.a(G380), .O(gate114inter7));
  inv1  gate807(.a(G381), .O(gate114inter8));
  nand2 gate808(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate809(.a(s_37), .b(gate114inter3), .O(gate114inter10));
  nor2  gate810(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate811(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate812(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2423(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2424(.a(gate119inter0), .b(s_268), .O(gate119inter1));
  and2  gate2425(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2426(.a(s_268), .O(gate119inter3));
  inv1  gate2427(.a(s_269), .O(gate119inter4));
  nand2 gate2428(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2429(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2430(.a(G390), .O(gate119inter7));
  inv1  gate2431(.a(G391), .O(gate119inter8));
  nand2 gate2432(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2433(.a(s_269), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2434(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2435(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2436(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1023(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1024(.a(gate126inter0), .b(s_68), .O(gate126inter1));
  and2  gate1025(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1026(.a(s_68), .O(gate126inter3));
  inv1  gate1027(.a(s_69), .O(gate126inter4));
  nand2 gate1028(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1029(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1030(.a(G404), .O(gate126inter7));
  inv1  gate1031(.a(G405), .O(gate126inter8));
  nand2 gate1032(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1033(.a(s_69), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1034(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1035(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1036(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1289(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1290(.a(gate130inter0), .b(s_106), .O(gate130inter1));
  and2  gate1291(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1292(.a(s_106), .O(gate130inter3));
  inv1  gate1293(.a(s_107), .O(gate130inter4));
  nand2 gate1294(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1295(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1296(.a(G412), .O(gate130inter7));
  inv1  gate1297(.a(G413), .O(gate130inter8));
  nand2 gate1298(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1299(.a(s_107), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1300(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1301(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1302(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate687(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate688(.a(gate135inter0), .b(s_20), .O(gate135inter1));
  and2  gate689(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate690(.a(s_20), .O(gate135inter3));
  inv1  gate691(.a(s_21), .O(gate135inter4));
  nand2 gate692(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate693(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate694(.a(G422), .O(gate135inter7));
  inv1  gate695(.a(G423), .O(gate135inter8));
  nand2 gate696(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate697(.a(s_21), .b(gate135inter3), .O(gate135inter10));
  nor2  gate698(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate699(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate700(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1471(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1472(.a(gate137inter0), .b(s_132), .O(gate137inter1));
  and2  gate1473(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1474(.a(s_132), .O(gate137inter3));
  inv1  gate1475(.a(s_133), .O(gate137inter4));
  nand2 gate1476(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1477(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1478(.a(G426), .O(gate137inter7));
  inv1  gate1479(.a(G429), .O(gate137inter8));
  nand2 gate1480(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1481(.a(s_133), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1482(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1483(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1484(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2059(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2060(.a(gate144inter0), .b(s_216), .O(gate144inter1));
  and2  gate2061(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2062(.a(s_216), .O(gate144inter3));
  inv1  gate2063(.a(s_217), .O(gate144inter4));
  nand2 gate2064(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2065(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2066(.a(G468), .O(gate144inter7));
  inv1  gate2067(.a(G471), .O(gate144inter8));
  nand2 gate2068(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2069(.a(s_217), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2070(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2071(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2072(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2241(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2242(.a(gate146inter0), .b(s_242), .O(gate146inter1));
  and2  gate2243(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2244(.a(s_242), .O(gate146inter3));
  inv1  gate2245(.a(s_243), .O(gate146inter4));
  nand2 gate2246(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2247(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2248(.a(G480), .O(gate146inter7));
  inv1  gate2249(.a(G483), .O(gate146inter8));
  nand2 gate2250(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2251(.a(s_243), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2252(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2253(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2254(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1009(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1010(.a(gate148inter0), .b(s_66), .O(gate148inter1));
  and2  gate1011(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1012(.a(s_66), .O(gate148inter3));
  inv1  gate1013(.a(s_67), .O(gate148inter4));
  nand2 gate1014(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1015(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1016(.a(G492), .O(gate148inter7));
  inv1  gate1017(.a(G495), .O(gate148inter8));
  nand2 gate1018(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1019(.a(s_67), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1020(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1021(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1022(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate2381(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate2382(.a(gate149inter0), .b(s_262), .O(gate149inter1));
  and2  gate2383(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate2384(.a(s_262), .O(gate149inter3));
  inv1  gate2385(.a(s_263), .O(gate149inter4));
  nand2 gate2386(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate2387(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate2388(.a(G498), .O(gate149inter7));
  inv1  gate2389(.a(G501), .O(gate149inter8));
  nand2 gate2390(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate2391(.a(s_263), .b(gate149inter3), .O(gate149inter10));
  nor2  gate2392(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate2393(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate2394(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1261(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1262(.a(gate153inter0), .b(s_102), .O(gate153inter1));
  and2  gate1263(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1264(.a(s_102), .O(gate153inter3));
  inv1  gate1265(.a(s_103), .O(gate153inter4));
  nand2 gate1266(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1267(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1268(.a(G426), .O(gate153inter7));
  inv1  gate1269(.a(G522), .O(gate153inter8));
  nand2 gate1270(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1271(.a(s_103), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1272(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1273(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1274(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1905(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1906(.a(gate154inter0), .b(s_194), .O(gate154inter1));
  and2  gate1907(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1908(.a(s_194), .O(gate154inter3));
  inv1  gate1909(.a(s_195), .O(gate154inter4));
  nand2 gate1910(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1911(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1912(.a(G429), .O(gate154inter7));
  inv1  gate1913(.a(G522), .O(gate154inter8));
  nand2 gate1914(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1915(.a(s_195), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1916(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1917(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1918(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1625(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1626(.a(gate155inter0), .b(s_154), .O(gate155inter1));
  and2  gate1627(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1628(.a(s_154), .O(gate155inter3));
  inv1  gate1629(.a(s_155), .O(gate155inter4));
  nand2 gate1630(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1631(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1632(.a(G432), .O(gate155inter7));
  inv1  gate1633(.a(G525), .O(gate155inter8));
  nand2 gate1634(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1635(.a(s_155), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1636(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1637(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1638(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1331(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1332(.a(gate156inter0), .b(s_112), .O(gate156inter1));
  and2  gate1333(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1334(.a(s_112), .O(gate156inter3));
  inv1  gate1335(.a(s_113), .O(gate156inter4));
  nand2 gate1336(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1337(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1338(.a(G435), .O(gate156inter7));
  inv1  gate1339(.a(G525), .O(gate156inter8));
  nand2 gate1340(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1341(.a(s_113), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1342(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1343(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1344(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1849(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1850(.a(gate159inter0), .b(s_186), .O(gate159inter1));
  and2  gate1851(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1852(.a(s_186), .O(gate159inter3));
  inv1  gate1853(.a(s_187), .O(gate159inter4));
  nand2 gate1854(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1855(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1856(.a(G444), .O(gate159inter7));
  inv1  gate1857(.a(G531), .O(gate159inter8));
  nand2 gate1858(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1859(.a(s_187), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1860(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1861(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1862(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1751(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1752(.a(gate162inter0), .b(s_172), .O(gate162inter1));
  and2  gate1753(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1754(.a(s_172), .O(gate162inter3));
  inv1  gate1755(.a(s_173), .O(gate162inter4));
  nand2 gate1756(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1757(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1758(.a(G453), .O(gate162inter7));
  inv1  gate1759(.a(G534), .O(gate162inter8));
  nand2 gate1760(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1761(.a(s_173), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1762(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1763(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1764(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1359(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1360(.a(gate164inter0), .b(s_116), .O(gate164inter1));
  and2  gate1361(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1362(.a(s_116), .O(gate164inter3));
  inv1  gate1363(.a(s_117), .O(gate164inter4));
  nand2 gate1364(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1365(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1366(.a(G459), .O(gate164inter7));
  inv1  gate1367(.a(G537), .O(gate164inter8));
  nand2 gate1368(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1369(.a(s_117), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1370(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1371(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1372(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2031(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2032(.a(gate166inter0), .b(s_212), .O(gate166inter1));
  and2  gate2033(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2034(.a(s_212), .O(gate166inter3));
  inv1  gate2035(.a(s_213), .O(gate166inter4));
  nand2 gate2036(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2037(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2038(.a(G465), .O(gate166inter7));
  inv1  gate2039(.a(G540), .O(gate166inter8));
  nand2 gate2040(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2041(.a(s_213), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2042(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2043(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2044(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1667(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1668(.a(gate168inter0), .b(s_160), .O(gate168inter1));
  and2  gate1669(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1670(.a(s_160), .O(gate168inter3));
  inv1  gate1671(.a(s_161), .O(gate168inter4));
  nand2 gate1672(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1673(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1674(.a(G471), .O(gate168inter7));
  inv1  gate1675(.a(G543), .O(gate168inter8));
  nand2 gate1676(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1677(.a(s_161), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1678(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1679(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1680(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2003(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2004(.a(gate169inter0), .b(s_208), .O(gate169inter1));
  and2  gate2005(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2006(.a(s_208), .O(gate169inter3));
  inv1  gate2007(.a(s_209), .O(gate169inter4));
  nand2 gate2008(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2009(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2010(.a(G474), .O(gate169inter7));
  inv1  gate2011(.a(G546), .O(gate169inter8));
  nand2 gate2012(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2013(.a(s_209), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2014(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2015(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2016(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate967(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate968(.a(gate172inter0), .b(s_60), .O(gate172inter1));
  and2  gate969(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate970(.a(s_60), .O(gate172inter3));
  inv1  gate971(.a(s_61), .O(gate172inter4));
  nand2 gate972(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate973(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate974(.a(G483), .O(gate172inter7));
  inv1  gate975(.a(G549), .O(gate172inter8));
  nand2 gate976(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate977(.a(s_61), .b(gate172inter3), .O(gate172inter10));
  nor2  gate978(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate979(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate980(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1723(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1724(.a(gate174inter0), .b(s_168), .O(gate174inter1));
  and2  gate1725(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1726(.a(s_168), .O(gate174inter3));
  inv1  gate1727(.a(s_169), .O(gate174inter4));
  nand2 gate1728(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1729(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1730(.a(G489), .O(gate174inter7));
  inv1  gate1731(.a(G552), .O(gate174inter8));
  nand2 gate1732(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1733(.a(s_169), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1734(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1735(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1736(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1121(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1122(.a(gate183inter0), .b(s_82), .O(gate183inter1));
  and2  gate1123(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1124(.a(s_82), .O(gate183inter3));
  inv1  gate1125(.a(s_83), .O(gate183inter4));
  nand2 gate1126(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1127(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1128(.a(G516), .O(gate183inter7));
  inv1  gate1129(.a(G567), .O(gate183inter8));
  nand2 gate1130(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1131(.a(s_83), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1132(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1133(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1134(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate995(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate996(.a(gate186inter0), .b(s_64), .O(gate186inter1));
  and2  gate997(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate998(.a(s_64), .O(gate186inter3));
  inv1  gate999(.a(s_65), .O(gate186inter4));
  nand2 gate1000(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1001(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1002(.a(G572), .O(gate186inter7));
  inv1  gate1003(.a(G573), .O(gate186inter8));
  nand2 gate1004(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1005(.a(s_65), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1006(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1007(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1008(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1807(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1808(.a(gate188inter0), .b(s_180), .O(gate188inter1));
  and2  gate1809(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1810(.a(s_180), .O(gate188inter3));
  inv1  gate1811(.a(s_181), .O(gate188inter4));
  nand2 gate1812(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1813(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1814(.a(G576), .O(gate188inter7));
  inv1  gate1815(.a(G577), .O(gate188inter8));
  nand2 gate1816(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1817(.a(s_181), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1818(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1819(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1820(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1821(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1822(.a(gate195inter0), .b(s_182), .O(gate195inter1));
  and2  gate1823(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1824(.a(s_182), .O(gate195inter3));
  inv1  gate1825(.a(s_183), .O(gate195inter4));
  nand2 gate1826(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1827(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1828(.a(G590), .O(gate195inter7));
  inv1  gate1829(.a(G591), .O(gate195inter8));
  nand2 gate1830(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1831(.a(s_183), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1832(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1833(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1834(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2437(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2438(.a(gate196inter0), .b(s_270), .O(gate196inter1));
  and2  gate2439(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2440(.a(s_270), .O(gate196inter3));
  inv1  gate2441(.a(s_271), .O(gate196inter4));
  nand2 gate2442(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2443(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2444(.a(G592), .O(gate196inter7));
  inv1  gate2445(.a(G593), .O(gate196inter8));
  nand2 gate2446(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2447(.a(s_271), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2448(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2449(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2450(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1303(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1304(.a(gate197inter0), .b(s_108), .O(gate197inter1));
  and2  gate1305(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1306(.a(s_108), .O(gate197inter3));
  inv1  gate1307(.a(s_109), .O(gate197inter4));
  nand2 gate1308(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1309(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1310(.a(G594), .O(gate197inter7));
  inv1  gate1311(.a(G595), .O(gate197inter8));
  nand2 gate1312(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1313(.a(s_109), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1314(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1315(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1316(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1737(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1738(.a(gate199inter0), .b(s_170), .O(gate199inter1));
  and2  gate1739(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1740(.a(s_170), .O(gate199inter3));
  inv1  gate1741(.a(s_171), .O(gate199inter4));
  nand2 gate1742(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1743(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1744(.a(G598), .O(gate199inter7));
  inv1  gate1745(.a(G599), .O(gate199inter8));
  nand2 gate1746(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1747(.a(s_171), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1748(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1749(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1750(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1233(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1234(.a(gate200inter0), .b(s_98), .O(gate200inter1));
  and2  gate1235(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1236(.a(s_98), .O(gate200inter3));
  inv1  gate1237(.a(s_99), .O(gate200inter4));
  nand2 gate1238(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1239(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1240(.a(G600), .O(gate200inter7));
  inv1  gate1241(.a(G601), .O(gate200inter8));
  nand2 gate1242(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1243(.a(s_99), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1244(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1245(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1246(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2311(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2312(.a(gate203inter0), .b(s_252), .O(gate203inter1));
  and2  gate2313(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2314(.a(s_252), .O(gate203inter3));
  inv1  gate2315(.a(s_253), .O(gate203inter4));
  nand2 gate2316(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2317(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2318(.a(G602), .O(gate203inter7));
  inv1  gate2319(.a(G612), .O(gate203inter8));
  nand2 gate2320(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2321(.a(s_253), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2322(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2323(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2324(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate2269(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2270(.a(gate204inter0), .b(s_246), .O(gate204inter1));
  and2  gate2271(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2272(.a(s_246), .O(gate204inter3));
  inv1  gate2273(.a(s_247), .O(gate204inter4));
  nand2 gate2274(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2275(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2276(.a(G607), .O(gate204inter7));
  inv1  gate2277(.a(G617), .O(gate204inter8));
  nand2 gate2278(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2279(.a(s_247), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2280(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2281(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2282(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1429(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1430(.a(gate205inter0), .b(s_126), .O(gate205inter1));
  and2  gate1431(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1432(.a(s_126), .O(gate205inter3));
  inv1  gate1433(.a(s_127), .O(gate205inter4));
  nand2 gate1434(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1435(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1436(.a(G622), .O(gate205inter7));
  inv1  gate1437(.a(G627), .O(gate205inter8));
  nand2 gate1438(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1439(.a(s_127), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1440(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1441(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1442(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1275(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1276(.a(gate207inter0), .b(s_104), .O(gate207inter1));
  and2  gate1277(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1278(.a(s_104), .O(gate207inter3));
  inv1  gate1279(.a(s_105), .O(gate207inter4));
  nand2 gate1280(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1281(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1282(.a(G622), .O(gate207inter7));
  inv1  gate1283(.a(G632), .O(gate207inter8));
  nand2 gate1284(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1285(.a(s_105), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1286(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1287(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1288(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate2283(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate2284(.a(gate209inter0), .b(s_248), .O(gate209inter1));
  and2  gate2285(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate2286(.a(s_248), .O(gate209inter3));
  inv1  gate2287(.a(s_249), .O(gate209inter4));
  nand2 gate2288(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate2289(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate2290(.a(G602), .O(gate209inter7));
  inv1  gate2291(.a(G666), .O(gate209inter8));
  nand2 gate2292(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate2293(.a(s_249), .b(gate209inter3), .O(gate209inter10));
  nor2  gate2294(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate2295(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate2296(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate911(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate912(.a(gate213inter0), .b(s_52), .O(gate213inter1));
  and2  gate913(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate914(.a(s_52), .O(gate213inter3));
  inv1  gate915(.a(s_53), .O(gate213inter4));
  nand2 gate916(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate917(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate918(.a(G602), .O(gate213inter7));
  inv1  gate919(.a(G672), .O(gate213inter8));
  nand2 gate920(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate921(.a(s_53), .b(gate213inter3), .O(gate213inter10));
  nor2  gate922(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate923(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate924(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2409(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2410(.a(gate215inter0), .b(s_266), .O(gate215inter1));
  and2  gate2411(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2412(.a(s_266), .O(gate215inter3));
  inv1  gate2413(.a(s_267), .O(gate215inter4));
  nand2 gate2414(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2415(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2416(.a(G607), .O(gate215inter7));
  inv1  gate2417(.a(G675), .O(gate215inter8));
  nand2 gate2418(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2419(.a(s_267), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2420(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2421(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2422(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1877(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1878(.a(gate217inter0), .b(s_190), .O(gate217inter1));
  and2  gate1879(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1880(.a(s_190), .O(gate217inter3));
  inv1  gate1881(.a(s_191), .O(gate217inter4));
  nand2 gate1882(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1883(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1884(.a(G622), .O(gate217inter7));
  inv1  gate1885(.a(G678), .O(gate217inter8));
  nand2 gate1886(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1887(.a(s_191), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1888(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1889(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1890(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate841(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate842(.a(gate222inter0), .b(s_42), .O(gate222inter1));
  and2  gate843(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate844(.a(s_42), .O(gate222inter3));
  inv1  gate845(.a(s_43), .O(gate222inter4));
  nand2 gate846(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate847(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate848(.a(G632), .O(gate222inter7));
  inv1  gate849(.a(G684), .O(gate222inter8));
  nand2 gate850(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate851(.a(s_43), .b(gate222inter3), .O(gate222inter10));
  nor2  gate852(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate853(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate854(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2199(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2200(.a(gate223inter0), .b(s_236), .O(gate223inter1));
  and2  gate2201(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2202(.a(s_236), .O(gate223inter3));
  inv1  gate2203(.a(s_237), .O(gate223inter4));
  nand2 gate2204(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2205(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2206(.a(G627), .O(gate223inter7));
  inv1  gate2207(.a(G687), .O(gate223inter8));
  nand2 gate2208(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2209(.a(s_237), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2210(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2211(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2212(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1037(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1038(.a(gate232inter0), .b(s_70), .O(gate232inter1));
  and2  gate1039(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1040(.a(s_70), .O(gate232inter3));
  inv1  gate1041(.a(s_71), .O(gate232inter4));
  nand2 gate1042(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1043(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1044(.a(G704), .O(gate232inter7));
  inv1  gate1045(.a(G705), .O(gate232inter8));
  nand2 gate1046(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1047(.a(s_71), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1048(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1049(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1050(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1317(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1318(.a(gate236inter0), .b(s_110), .O(gate236inter1));
  and2  gate1319(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1320(.a(s_110), .O(gate236inter3));
  inv1  gate1321(.a(s_111), .O(gate236inter4));
  nand2 gate1322(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1323(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1324(.a(G251), .O(gate236inter7));
  inv1  gate1325(.a(G727), .O(gate236inter8));
  nand2 gate1326(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1327(.a(s_111), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1328(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1329(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1330(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1653(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1654(.a(gate238inter0), .b(s_158), .O(gate238inter1));
  and2  gate1655(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1656(.a(s_158), .O(gate238inter3));
  inv1  gate1657(.a(s_159), .O(gate238inter4));
  nand2 gate1658(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1659(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1660(.a(G257), .O(gate238inter7));
  inv1  gate1661(.a(G709), .O(gate238inter8));
  nand2 gate1662(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1663(.a(s_159), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1664(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1665(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1666(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1345(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1346(.a(gate241inter0), .b(s_114), .O(gate241inter1));
  and2  gate1347(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1348(.a(s_114), .O(gate241inter3));
  inv1  gate1349(.a(s_115), .O(gate241inter4));
  nand2 gate1350(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1351(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1352(.a(G242), .O(gate241inter7));
  inv1  gate1353(.a(G730), .O(gate241inter8));
  nand2 gate1354(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1355(.a(s_115), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1356(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1357(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1358(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1611(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1612(.a(gate242inter0), .b(s_152), .O(gate242inter1));
  and2  gate1613(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1614(.a(s_152), .O(gate242inter3));
  inv1  gate1615(.a(s_153), .O(gate242inter4));
  nand2 gate1616(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1617(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1618(.a(G718), .O(gate242inter7));
  inv1  gate1619(.a(G730), .O(gate242inter8));
  nand2 gate1620(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1621(.a(s_153), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1622(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1623(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1624(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1597(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1598(.a(gate250inter0), .b(s_150), .O(gate250inter1));
  and2  gate1599(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1600(.a(s_150), .O(gate250inter3));
  inv1  gate1601(.a(s_151), .O(gate250inter4));
  nand2 gate1602(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1603(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1604(.a(G706), .O(gate250inter7));
  inv1  gate1605(.a(G742), .O(gate250inter8));
  nand2 gate1606(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1607(.a(s_151), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1608(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1609(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1610(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1387(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1388(.a(gate253inter0), .b(s_120), .O(gate253inter1));
  and2  gate1389(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1390(.a(s_120), .O(gate253inter3));
  inv1  gate1391(.a(s_121), .O(gate253inter4));
  nand2 gate1392(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1393(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1394(.a(G260), .O(gate253inter7));
  inv1  gate1395(.a(G748), .O(gate253inter8));
  nand2 gate1396(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1397(.a(s_121), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1398(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1399(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1400(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1485(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1486(.a(gate256inter0), .b(s_134), .O(gate256inter1));
  and2  gate1487(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1488(.a(s_134), .O(gate256inter3));
  inv1  gate1489(.a(s_135), .O(gate256inter4));
  nand2 gate1490(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1491(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1492(.a(G715), .O(gate256inter7));
  inv1  gate1493(.a(G751), .O(gate256inter8));
  nand2 gate1494(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1495(.a(s_135), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1496(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1497(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1498(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1765(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1766(.a(gate259inter0), .b(s_174), .O(gate259inter1));
  and2  gate1767(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1768(.a(s_174), .O(gate259inter3));
  inv1  gate1769(.a(s_175), .O(gate259inter4));
  nand2 gate1770(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1771(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1772(.a(G758), .O(gate259inter7));
  inv1  gate1773(.a(G759), .O(gate259inter8));
  nand2 gate1774(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1775(.a(s_175), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1776(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1777(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1778(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1639(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1640(.a(gate262inter0), .b(s_156), .O(gate262inter1));
  and2  gate1641(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1642(.a(s_156), .O(gate262inter3));
  inv1  gate1643(.a(s_157), .O(gate262inter4));
  nand2 gate1644(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1645(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1646(.a(G764), .O(gate262inter7));
  inv1  gate1647(.a(G765), .O(gate262inter8));
  nand2 gate1648(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1649(.a(s_157), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1650(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1651(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1652(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate981(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate982(.a(gate264inter0), .b(s_62), .O(gate264inter1));
  and2  gate983(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate984(.a(s_62), .O(gate264inter3));
  inv1  gate985(.a(s_63), .O(gate264inter4));
  nand2 gate986(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate987(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate988(.a(G768), .O(gate264inter7));
  inv1  gate989(.a(G769), .O(gate264inter8));
  nand2 gate990(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate991(.a(s_63), .b(gate264inter3), .O(gate264inter10));
  nor2  gate992(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate993(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate994(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2017(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2018(.a(gate269inter0), .b(s_210), .O(gate269inter1));
  and2  gate2019(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2020(.a(s_210), .O(gate269inter3));
  inv1  gate2021(.a(s_211), .O(gate269inter4));
  nand2 gate2022(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2023(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2024(.a(G654), .O(gate269inter7));
  inv1  gate2025(.a(G782), .O(gate269inter8));
  nand2 gate2026(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2027(.a(s_211), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2028(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2029(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2030(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2045(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2046(.a(gate271inter0), .b(s_214), .O(gate271inter1));
  and2  gate2047(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2048(.a(s_214), .O(gate271inter3));
  inv1  gate2049(.a(s_215), .O(gate271inter4));
  nand2 gate2050(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2051(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2052(.a(G660), .O(gate271inter7));
  inv1  gate2053(.a(G788), .O(gate271inter8));
  nand2 gate2054(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2055(.a(s_215), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2056(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2057(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2058(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1065(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1066(.a(gate272inter0), .b(s_74), .O(gate272inter1));
  and2  gate1067(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1068(.a(s_74), .O(gate272inter3));
  inv1  gate1069(.a(s_75), .O(gate272inter4));
  nand2 gate1070(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1071(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1072(.a(G663), .O(gate272inter7));
  inv1  gate1073(.a(G791), .O(gate272inter8));
  nand2 gate1074(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1075(.a(s_75), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1076(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1077(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1078(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1863(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1864(.a(gate273inter0), .b(s_188), .O(gate273inter1));
  and2  gate1865(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1866(.a(s_188), .O(gate273inter3));
  inv1  gate1867(.a(s_189), .O(gate273inter4));
  nand2 gate1868(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1869(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1870(.a(G642), .O(gate273inter7));
  inv1  gate1871(.a(G794), .O(gate273inter8));
  nand2 gate1872(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1873(.a(s_189), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1874(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1875(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1876(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate603(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate604(.a(gate274inter0), .b(s_8), .O(gate274inter1));
  and2  gate605(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate606(.a(s_8), .O(gate274inter3));
  inv1  gate607(.a(s_9), .O(gate274inter4));
  nand2 gate608(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate609(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate610(.a(G770), .O(gate274inter7));
  inv1  gate611(.a(G794), .O(gate274inter8));
  nand2 gate612(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate613(.a(s_9), .b(gate274inter3), .O(gate274inter10));
  nor2  gate614(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate615(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate616(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate757(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate758(.a(gate278inter0), .b(s_30), .O(gate278inter1));
  and2  gate759(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate760(.a(s_30), .O(gate278inter3));
  inv1  gate761(.a(s_31), .O(gate278inter4));
  nand2 gate762(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate763(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate764(.a(G776), .O(gate278inter7));
  inv1  gate765(.a(G800), .O(gate278inter8));
  nand2 gate766(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate767(.a(s_31), .b(gate278inter3), .O(gate278inter10));
  nor2  gate768(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate769(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate770(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1149(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1150(.a(gate279inter0), .b(s_86), .O(gate279inter1));
  and2  gate1151(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1152(.a(s_86), .O(gate279inter3));
  inv1  gate1153(.a(s_87), .O(gate279inter4));
  nand2 gate1154(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1155(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1156(.a(G651), .O(gate279inter7));
  inv1  gate1157(.a(G803), .O(gate279inter8));
  nand2 gate1158(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1159(.a(s_87), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1160(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1161(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1162(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1079(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1080(.a(gate281inter0), .b(s_76), .O(gate281inter1));
  and2  gate1081(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1082(.a(s_76), .O(gate281inter3));
  inv1  gate1083(.a(s_77), .O(gate281inter4));
  nand2 gate1084(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1085(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1086(.a(G654), .O(gate281inter7));
  inv1  gate1087(.a(G806), .O(gate281inter8));
  nand2 gate1088(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1089(.a(s_77), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1090(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1091(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1092(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2353(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2354(.a(gate282inter0), .b(s_258), .O(gate282inter1));
  and2  gate2355(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2356(.a(s_258), .O(gate282inter3));
  inv1  gate2357(.a(s_259), .O(gate282inter4));
  nand2 gate2358(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2359(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2360(.a(G782), .O(gate282inter7));
  inv1  gate2361(.a(G806), .O(gate282inter8));
  nand2 gate2362(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2363(.a(s_259), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2364(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2365(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2366(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate771(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate772(.a(gate291inter0), .b(s_32), .O(gate291inter1));
  and2  gate773(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate774(.a(s_32), .O(gate291inter3));
  inv1  gate775(.a(s_33), .O(gate291inter4));
  nand2 gate776(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate777(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate778(.a(G822), .O(gate291inter7));
  inv1  gate779(.a(G823), .O(gate291inter8));
  nand2 gate780(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate781(.a(s_33), .b(gate291inter3), .O(gate291inter10));
  nor2  gate782(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate783(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate784(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate547(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate548(.a(gate292inter0), .b(s_0), .O(gate292inter1));
  and2  gate549(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate550(.a(s_0), .O(gate292inter3));
  inv1  gate551(.a(s_1), .O(gate292inter4));
  nand2 gate552(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate553(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate554(.a(G824), .O(gate292inter7));
  inv1  gate555(.a(G825), .O(gate292inter8));
  nand2 gate556(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate557(.a(s_1), .b(gate292inter3), .O(gate292inter10));
  nor2  gate558(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate559(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate560(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate2101(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2102(.a(gate293inter0), .b(s_222), .O(gate293inter1));
  and2  gate2103(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2104(.a(s_222), .O(gate293inter3));
  inv1  gate2105(.a(s_223), .O(gate293inter4));
  nand2 gate2106(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2107(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2108(.a(G828), .O(gate293inter7));
  inv1  gate2109(.a(G829), .O(gate293inter8));
  nand2 gate2110(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2111(.a(s_223), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2112(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2113(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2114(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1933(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1934(.a(gate389inter0), .b(s_198), .O(gate389inter1));
  and2  gate1935(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1936(.a(s_198), .O(gate389inter3));
  inv1  gate1937(.a(s_199), .O(gate389inter4));
  nand2 gate1938(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1939(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1940(.a(G3), .O(gate389inter7));
  inv1  gate1941(.a(G1042), .O(gate389inter8));
  nand2 gate1942(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1943(.a(s_199), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1944(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1945(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1946(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1569(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1570(.a(gate395inter0), .b(s_146), .O(gate395inter1));
  and2  gate1571(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1572(.a(s_146), .O(gate395inter3));
  inv1  gate1573(.a(s_147), .O(gate395inter4));
  nand2 gate1574(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1575(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1576(.a(G9), .O(gate395inter7));
  inv1  gate1577(.a(G1060), .O(gate395inter8));
  nand2 gate1578(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1579(.a(s_147), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1580(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1581(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1582(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1947(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1948(.a(gate399inter0), .b(s_200), .O(gate399inter1));
  and2  gate1949(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1950(.a(s_200), .O(gate399inter3));
  inv1  gate1951(.a(s_201), .O(gate399inter4));
  nand2 gate1952(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1953(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1954(.a(G13), .O(gate399inter7));
  inv1  gate1955(.a(G1072), .O(gate399inter8));
  nand2 gate1956(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1957(.a(s_201), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1958(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1959(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1960(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate589(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate590(.a(gate400inter0), .b(s_6), .O(gate400inter1));
  and2  gate591(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate592(.a(s_6), .O(gate400inter3));
  inv1  gate593(.a(s_7), .O(gate400inter4));
  nand2 gate594(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate595(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate596(.a(G14), .O(gate400inter7));
  inv1  gate597(.a(G1075), .O(gate400inter8));
  nand2 gate598(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate599(.a(s_7), .b(gate400inter3), .O(gate400inter10));
  nor2  gate600(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate601(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate602(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1499(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1500(.a(gate404inter0), .b(s_136), .O(gate404inter1));
  and2  gate1501(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1502(.a(s_136), .O(gate404inter3));
  inv1  gate1503(.a(s_137), .O(gate404inter4));
  nand2 gate1504(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1505(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1506(.a(G18), .O(gate404inter7));
  inv1  gate1507(.a(G1087), .O(gate404inter8));
  nand2 gate1508(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1509(.a(s_137), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1510(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1511(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1512(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1247(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1248(.a(gate405inter0), .b(s_100), .O(gate405inter1));
  and2  gate1249(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1250(.a(s_100), .O(gate405inter3));
  inv1  gate1251(.a(s_101), .O(gate405inter4));
  nand2 gate1252(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1253(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1254(.a(G19), .O(gate405inter7));
  inv1  gate1255(.a(G1090), .O(gate405inter8));
  nand2 gate1256(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1257(.a(s_101), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1258(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1259(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1260(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1093(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1094(.a(gate406inter0), .b(s_78), .O(gate406inter1));
  and2  gate1095(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1096(.a(s_78), .O(gate406inter3));
  inv1  gate1097(.a(s_79), .O(gate406inter4));
  nand2 gate1098(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1099(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1100(.a(G20), .O(gate406inter7));
  inv1  gate1101(.a(G1093), .O(gate406inter8));
  nand2 gate1102(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1103(.a(s_79), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1104(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1105(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1106(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate953(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate954(.a(gate410inter0), .b(s_58), .O(gate410inter1));
  and2  gate955(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate956(.a(s_58), .O(gate410inter3));
  inv1  gate957(.a(s_59), .O(gate410inter4));
  nand2 gate958(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate959(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate960(.a(G24), .O(gate410inter7));
  inv1  gate961(.a(G1105), .O(gate410inter8));
  nand2 gate962(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate963(.a(s_59), .b(gate410inter3), .O(gate410inter10));
  nor2  gate964(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate965(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate966(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1793(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1794(.a(gate411inter0), .b(s_178), .O(gate411inter1));
  and2  gate1795(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1796(.a(s_178), .O(gate411inter3));
  inv1  gate1797(.a(s_179), .O(gate411inter4));
  nand2 gate1798(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1799(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1800(.a(G25), .O(gate411inter7));
  inv1  gate1801(.a(G1108), .O(gate411inter8));
  nand2 gate1802(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1803(.a(s_179), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1804(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1805(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1806(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate897(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate898(.a(gate412inter0), .b(s_50), .O(gate412inter1));
  and2  gate899(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate900(.a(s_50), .O(gate412inter3));
  inv1  gate901(.a(s_51), .O(gate412inter4));
  nand2 gate902(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate903(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate904(.a(G26), .O(gate412inter7));
  inv1  gate905(.a(G1111), .O(gate412inter8));
  nand2 gate906(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate907(.a(s_51), .b(gate412inter3), .O(gate412inter10));
  nor2  gate908(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate909(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate910(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1415(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1416(.a(gate413inter0), .b(s_124), .O(gate413inter1));
  and2  gate1417(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1418(.a(s_124), .O(gate413inter3));
  inv1  gate1419(.a(s_125), .O(gate413inter4));
  nand2 gate1420(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1421(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1422(.a(G27), .O(gate413inter7));
  inv1  gate1423(.a(G1114), .O(gate413inter8));
  nand2 gate1424(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1425(.a(s_125), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1426(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1427(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1428(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1891(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1892(.a(gate416inter0), .b(s_192), .O(gate416inter1));
  and2  gate1893(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1894(.a(s_192), .O(gate416inter3));
  inv1  gate1895(.a(s_193), .O(gate416inter4));
  nand2 gate1896(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1897(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1898(.a(G30), .O(gate416inter7));
  inv1  gate1899(.a(G1123), .O(gate416inter8));
  nand2 gate1900(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1901(.a(s_193), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1902(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1903(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1904(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2143(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2144(.a(gate426inter0), .b(s_228), .O(gate426inter1));
  and2  gate2145(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2146(.a(s_228), .O(gate426inter3));
  inv1  gate2147(.a(s_229), .O(gate426inter4));
  nand2 gate2148(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2149(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2150(.a(G1045), .O(gate426inter7));
  inv1  gate2151(.a(G1141), .O(gate426inter8));
  nand2 gate2152(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2153(.a(s_229), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2154(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2155(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2156(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate869(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate870(.a(gate430inter0), .b(s_46), .O(gate430inter1));
  and2  gate871(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate872(.a(s_46), .O(gate430inter3));
  inv1  gate873(.a(s_47), .O(gate430inter4));
  nand2 gate874(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate875(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate876(.a(G1051), .O(gate430inter7));
  inv1  gate877(.a(G1147), .O(gate430inter8));
  nand2 gate878(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate879(.a(s_47), .b(gate430inter3), .O(gate430inter10));
  nor2  gate880(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate881(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate882(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1373(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1374(.a(gate432inter0), .b(s_118), .O(gate432inter1));
  and2  gate1375(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1376(.a(s_118), .O(gate432inter3));
  inv1  gate1377(.a(s_119), .O(gate432inter4));
  nand2 gate1378(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1379(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1380(.a(G1054), .O(gate432inter7));
  inv1  gate1381(.a(G1150), .O(gate432inter8));
  nand2 gate1382(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1383(.a(s_119), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1384(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1385(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1386(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate1989(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate1990(.a(gate436inter0), .b(s_206), .O(gate436inter1));
  and2  gate1991(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate1992(.a(s_206), .O(gate436inter3));
  inv1  gate1993(.a(s_207), .O(gate436inter4));
  nand2 gate1994(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate1995(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate1996(.a(G1060), .O(gate436inter7));
  inv1  gate1997(.a(G1156), .O(gate436inter8));
  nand2 gate1998(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate1999(.a(s_207), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2000(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2001(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2002(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate645(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate646(.a(gate439inter0), .b(s_14), .O(gate439inter1));
  and2  gate647(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate648(.a(s_14), .O(gate439inter3));
  inv1  gate649(.a(s_15), .O(gate439inter4));
  nand2 gate650(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate651(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate652(.a(G11), .O(gate439inter7));
  inv1  gate653(.a(G1162), .O(gate439inter8));
  nand2 gate654(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate655(.a(s_15), .b(gate439inter3), .O(gate439inter10));
  nor2  gate656(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate657(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate658(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate813(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate814(.a(gate440inter0), .b(s_38), .O(gate440inter1));
  and2  gate815(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate816(.a(s_38), .O(gate440inter3));
  inv1  gate817(.a(s_39), .O(gate440inter4));
  nand2 gate818(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate819(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate820(.a(G1066), .O(gate440inter7));
  inv1  gate821(.a(G1162), .O(gate440inter8));
  nand2 gate822(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate823(.a(s_39), .b(gate440inter3), .O(gate440inter10));
  nor2  gate824(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate825(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate826(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1709(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1710(.a(gate441inter0), .b(s_166), .O(gate441inter1));
  and2  gate1711(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1712(.a(s_166), .O(gate441inter3));
  inv1  gate1713(.a(s_167), .O(gate441inter4));
  nand2 gate1714(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1715(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1716(.a(G12), .O(gate441inter7));
  inv1  gate1717(.a(G1165), .O(gate441inter8));
  nand2 gate1718(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1719(.a(s_167), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1720(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1721(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1722(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1975(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1976(.a(gate442inter0), .b(s_204), .O(gate442inter1));
  and2  gate1977(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1978(.a(s_204), .O(gate442inter3));
  inv1  gate1979(.a(s_205), .O(gate442inter4));
  nand2 gate1980(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1981(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1982(.a(G1069), .O(gate442inter7));
  inv1  gate1983(.a(G1165), .O(gate442inter8));
  nand2 gate1984(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1985(.a(s_205), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1986(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1987(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1988(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate2185(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2186(.a(gate443inter0), .b(s_234), .O(gate443inter1));
  and2  gate2187(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2188(.a(s_234), .O(gate443inter3));
  inv1  gate2189(.a(s_235), .O(gate443inter4));
  nand2 gate2190(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2191(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2192(.a(G13), .O(gate443inter7));
  inv1  gate2193(.a(G1168), .O(gate443inter8));
  nand2 gate2194(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2195(.a(s_235), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2196(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2197(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2198(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2073(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2074(.a(gate445inter0), .b(s_218), .O(gate445inter1));
  and2  gate2075(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2076(.a(s_218), .O(gate445inter3));
  inv1  gate2077(.a(s_219), .O(gate445inter4));
  nand2 gate2078(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2079(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2080(.a(G14), .O(gate445inter7));
  inv1  gate2081(.a(G1171), .O(gate445inter8));
  nand2 gate2082(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2083(.a(s_219), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2084(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2085(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2086(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1443(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1444(.a(gate448inter0), .b(s_128), .O(gate448inter1));
  and2  gate1445(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1446(.a(s_128), .O(gate448inter3));
  inv1  gate1447(.a(s_129), .O(gate448inter4));
  nand2 gate1448(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1449(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1450(.a(G1078), .O(gate448inter7));
  inv1  gate1451(.a(G1174), .O(gate448inter8));
  nand2 gate1452(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1453(.a(s_129), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1454(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1455(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1456(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2227(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2228(.a(gate451inter0), .b(s_240), .O(gate451inter1));
  and2  gate2229(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2230(.a(s_240), .O(gate451inter3));
  inv1  gate2231(.a(s_241), .O(gate451inter4));
  nand2 gate2232(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2233(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2234(.a(G17), .O(gate451inter7));
  inv1  gate2235(.a(G1180), .O(gate451inter8));
  nand2 gate2236(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2237(.a(s_241), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2238(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2239(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2240(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate855(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate856(.a(gate453inter0), .b(s_44), .O(gate453inter1));
  and2  gate857(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate858(.a(s_44), .O(gate453inter3));
  inv1  gate859(.a(s_45), .O(gate453inter4));
  nand2 gate860(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate861(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate862(.a(G18), .O(gate453inter7));
  inv1  gate863(.a(G1183), .O(gate453inter8));
  nand2 gate864(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate865(.a(s_45), .b(gate453inter3), .O(gate453inter10));
  nor2  gate866(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate867(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate868(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate673(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate674(.a(gate455inter0), .b(s_18), .O(gate455inter1));
  and2  gate675(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate676(.a(s_18), .O(gate455inter3));
  inv1  gate677(.a(s_19), .O(gate455inter4));
  nand2 gate678(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate679(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate680(.a(G19), .O(gate455inter7));
  inv1  gate681(.a(G1186), .O(gate455inter8));
  nand2 gate682(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate683(.a(s_19), .b(gate455inter3), .O(gate455inter10));
  nor2  gate684(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate685(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate686(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1177(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1178(.a(gate457inter0), .b(s_90), .O(gate457inter1));
  and2  gate1179(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1180(.a(s_90), .O(gate457inter3));
  inv1  gate1181(.a(s_91), .O(gate457inter4));
  nand2 gate1182(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1183(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1184(.a(G20), .O(gate457inter7));
  inv1  gate1185(.a(G1189), .O(gate457inter8));
  nand2 gate1186(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1187(.a(s_91), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1188(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1189(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1190(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate2157(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate2158(.a(gate459inter0), .b(s_230), .O(gate459inter1));
  and2  gate2159(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate2160(.a(s_230), .O(gate459inter3));
  inv1  gate2161(.a(s_231), .O(gate459inter4));
  nand2 gate2162(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate2163(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate2164(.a(G21), .O(gate459inter7));
  inv1  gate2165(.a(G1192), .O(gate459inter8));
  nand2 gate2166(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate2167(.a(s_231), .b(gate459inter3), .O(gate459inter10));
  nor2  gate2168(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate2169(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate2170(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1583(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1584(.a(gate460inter0), .b(s_148), .O(gate460inter1));
  and2  gate1585(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1586(.a(s_148), .O(gate460inter3));
  inv1  gate1587(.a(s_149), .O(gate460inter4));
  nand2 gate1588(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1589(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1590(.a(G1096), .O(gate460inter7));
  inv1  gate1591(.a(G1192), .O(gate460inter8));
  nand2 gate1592(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1593(.a(s_149), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1594(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1595(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1596(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate925(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate926(.a(gate463inter0), .b(s_54), .O(gate463inter1));
  and2  gate927(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate928(.a(s_54), .O(gate463inter3));
  inv1  gate929(.a(s_55), .O(gate463inter4));
  nand2 gate930(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate931(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate932(.a(G23), .O(gate463inter7));
  inv1  gate933(.a(G1198), .O(gate463inter8));
  nand2 gate934(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate935(.a(s_55), .b(gate463inter3), .O(gate463inter10));
  nor2  gate936(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate937(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate938(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1695(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1696(.a(gate468inter0), .b(s_164), .O(gate468inter1));
  and2  gate1697(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1698(.a(s_164), .O(gate468inter3));
  inv1  gate1699(.a(s_165), .O(gate468inter4));
  nand2 gate1700(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1701(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1702(.a(G1108), .O(gate468inter7));
  inv1  gate1703(.a(G1204), .O(gate468inter8));
  nand2 gate1704(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1705(.a(s_165), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1706(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1707(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1708(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1541(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1542(.a(gate475inter0), .b(s_142), .O(gate475inter1));
  and2  gate1543(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1544(.a(s_142), .O(gate475inter3));
  inv1  gate1545(.a(s_143), .O(gate475inter4));
  nand2 gate1546(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1547(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1548(.a(G29), .O(gate475inter7));
  inv1  gate1549(.a(G1216), .O(gate475inter8));
  nand2 gate1550(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1551(.a(s_143), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1552(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1553(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1554(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate2171(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2172(.a(gate476inter0), .b(s_232), .O(gate476inter1));
  and2  gate2173(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2174(.a(s_232), .O(gate476inter3));
  inv1  gate2175(.a(s_233), .O(gate476inter4));
  nand2 gate2176(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2177(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2178(.a(G1120), .O(gate476inter7));
  inv1  gate2179(.a(G1216), .O(gate476inter8));
  nand2 gate2180(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2181(.a(s_233), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2182(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2183(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2184(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2087(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2088(.a(gate482inter0), .b(s_220), .O(gate482inter1));
  and2  gate2089(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2090(.a(s_220), .O(gate482inter3));
  inv1  gate2091(.a(s_221), .O(gate482inter4));
  nand2 gate2092(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2093(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2094(.a(G1129), .O(gate482inter7));
  inv1  gate2095(.a(G1225), .O(gate482inter8));
  nand2 gate2096(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2097(.a(s_221), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2098(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2099(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2100(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1457(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1458(.a(gate485inter0), .b(s_130), .O(gate485inter1));
  and2  gate1459(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1460(.a(s_130), .O(gate485inter3));
  inv1  gate1461(.a(s_131), .O(gate485inter4));
  nand2 gate1462(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1463(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1464(.a(G1232), .O(gate485inter7));
  inv1  gate1465(.a(G1233), .O(gate485inter8));
  nand2 gate1466(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1467(.a(s_131), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1468(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1469(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1470(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1051(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1052(.a(gate487inter0), .b(s_72), .O(gate487inter1));
  and2  gate1053(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1054(.a(s_72), .O(gate487inter3));
  inv1  gate1055(.a(s_73), .O(gate487inter4));
  nand2 gate1056(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1057(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1058(.a(G1236), .O(gate487inter7));
  inv1  gate1059(.a(G1237), .O(gate487inter8));
  nand2 gate1060(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1061(.a(s_73), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1062(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1063(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1064(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2325(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2326(.a(gate490inter0), .b(s_254), .O(gate490inter1));
  and2  gate2327(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2328(.a(s_254), .O(gate490inter3));
  inv1  gate2329(.a(s_255), .O(gate490inter4));
  nand2 gate2330(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2331(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2332(.a(G1242), .O(gate490inter7));
  inv1  gate2333(.a(G1243), .O(gate490inter8));
  nand2 gate2334(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2335(.a(s_255), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2336(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2337(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2338(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate827(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate828(.a(gate491inter0), .b(s_40), .O(gate491inter1));
  and2  gate829(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate830(.a(s_40), .O(gate491inter3));
  inv1  gate831(.a(s_41), .O(gate491inter4));
  nand2 gate832(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate833(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate834(.a(G1244), .O(gate491inter7));
  inv1  gate835(.a(G1245), .O(gate491inter8));
  nand2 gate836(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate837(.a(s_41), .b(gate491inter3), .O(gate491inter10));
  nor2  gate838(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate839(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate840(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate785(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate786(.a(gate492inter0), .b(s_34), .O(gate492inter1));
  and2  gate787(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate788(.a(s_34), .O(gate492inter3));
  inv1  gate789(.a(s_35), .O(gate492inter4));
  nand2 gate790(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate791(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate792(.a(G1246), .O(gate492inter7));
  inv1  gate793(.a(G1247), .O(gate492inter8));
  nand2 gate794(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate795(.a(s_35), .b(gate492inter3), .O(gate492inter10));
  nor2  gate796(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate797(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate798(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2129(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2130(.a(gate497inter0), .b(s_226), .O(gate497inter1));
  and2  gate2131(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2132(.a(s_226), .O(gate497inter3));
  inv1  gate2133(.a(s_227), .O(gate497inter4));
  nand2 gate2134(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2135(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2136(.a(G1256), .O(gate497inter7));
  inv1  gate2137(.a(G1257), .O(gate497inter8));
  nand2 gate2138(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2139(.a(s_227), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2140(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2141(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2142(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1527(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1528(.a(gate510inter0), .b(s_140), .O(gate510inter1));
  and2  gate1529(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1530(.a(s_140), .O(gate510inter3));
  inv1  gate1531(.a(s_141), .O(gate510inter4));
  nand2 gate1532(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1533(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1534(.a(G1282), .O(gate510inter7));
  inv1  gate1535(.a(G1283), .O(gate510inter8));
  nand2 gate1536(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1537(.a(s_141), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1538(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1539(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1540(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate729(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate730(.a(gate511inter0), .b(s_26), .O(gate511inter1));
  and2  gate731(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate732(.a(s_26), .O(gate511inter3));
  inv1  gate733(.a(s_27), .O(gate511inter4));
  nand2 gate734(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate735(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate736(.a(G1284), .O(gate511inter7));
  inv1  gate737(.a(G1285), .O(gate511inter8));
  nand2 gate738(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate739(.a(s_27), .b(gate511inter3), .O(gate511inter10));
  nor2  gate740(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate741(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate742(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule