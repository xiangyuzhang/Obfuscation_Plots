module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1723(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1724(.a(gate9inter0), .b(s_168), .O(gate9inter1));
  and2  gate1725(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1726(.a(s_168), .O(gate9inter3));
  inv1  gate1727(.a(s_169), .O(gate9inter4));
  nand2 gate1728(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1729(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1730(.a(G1), .O(gate9inter7));
  inv1  gate1731(.a(G2), .O(gate9inter8));
  nand2 gate1732(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1733(.a(s_169), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1734(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1735(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1736(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1947(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1948(.a(gate10inter0), .b(s_200), .O(gate10inter1));
  and2  gate1949(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1950(.a(s_200), .O(gate10inter3));
  inv1  gate1951(.a(s_201), .O(gate10inter4));
  nand2 gate1952(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1953(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1954(.a(G3), .O(gate10inter7));
  inv1  gate1955(.a(G4), .O(gate10inter8));
  nand2 gate1956(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1957(.a(s_201), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1958(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1959(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1960(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1247(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1248(.a(gate23inter0), .b(s_100), .O(gate23inter1));
  and2  gate1249(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1250(.a(s_100), .O(gate23inter3));
  inv1  gate1251(.a(s_101), .O(gate23inter4));
  nand2 gate1252(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1253(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1254(.a(G29), .O(gate23inter7));
  inv1  gate1255(.a(G30), .O(gate23inter8));
  nand2 gate1256(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1257(.a(s_101), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1258(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1259(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1260(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1191(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1192(.a(gate26inter0), .b(s_92), .O(gate26inter1));
  and2  gate1193(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1194(.a(s_92), .O(gate26inter3));
  inv1  gate1195(.a(s_93), .O(gate26inter4));
  nand2 gate1196(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1197(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1198(.a(G9), .O(gate26inter7));
  inv1  gate1199(.a(G13), .O(gate26inter8));
  nand2 gate1200(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1201(.a(s_93), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1202(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1203(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1204(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate1961(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1962(.a(gate27inter0), .b(s_202), .O(gate27inter1));
  and2  gate1963(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1964(.a(s_202), .O(gate27inter3));
  inv1  gate1965(.a(s_203), .O(gate27inter4));
  nand2 gate1966(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1967(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1968(.a(G2), .O(gate27inter7));
  inv1  gate1969(.a(G6), .O(gate27inter8));
  nand2 gate1970(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1971(.a(s_203), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1972(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1973(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1974(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1275(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1276(.a(gate33inter0), .b(s_104), .O(gate33inter1));
  and2  gate1277(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1278(.a(s_104), .O(gate33inter3));
  inv1  gate1279(.a(s_105), .O(gate33inter4));
  nand2 gate1280(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1281(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1282(.a(G17), .O(gate33inter7));
  inv1  gate1283(.a(G21), .O(gate33inter8));
  nand2 gate1284(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1285(.a(s_105), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1286(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1287(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1288(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate771(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate772(.a(gate34inter0), .b(s_32), .O(gate34inter1));
  and2  gate773(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate774(.a(s_32), .O(gate34inter3));
  inv1  gate775(.a(s_33), .O(gate34inter4));
  nand2 gate776(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate777(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate778(.a(G25), .O(gate34inter7));
  inv1  gate779(.a(G29), .O(gate34inter8));
  nand2 gate780(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate781(.a(s_33), .b(gate34inter3), .O(gate34inter10));
  nor2  gate782(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate783(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate784(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate631(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate632(.a(gate37inter0), .b(s_12), .O(gate37inter1));
  and2  gate633(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate634(.a(s_12), .O(gate37inter3));
  inv1  gate635(.a(s_13), .O(gate37inter4));
  nand2 gate636(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate637(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate638(.a(G19), .O(gate37inter7));
  inv1  gate639(.a(G23), .O(gate37inter8));
  nand2 gate640(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate641(.a(s_13), .b(gate37inter3), .O(gate37inter10));
  nor2  gate642(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate643(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate644(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1065(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1066(.a(gate40inter0), .b(s_74), .O(gate40inter1));
  and2  gate1067(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1068(.a(s_74), .O(gate40inter3));
  inv1  gate1069(.a(s_75), .O(gate40inter4));
  nand2 gate1070(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1071(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1072(.a(G28), .O(gate40inter7));
  inv1  gate1073(.a(G32), .O(gate40inter8));
  nand2 gate1074(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1075(.a(s_75), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1076(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1077(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1078(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1079(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1080(.a(gate41inter0), .b(s_76), .O(gate41inter1));
  and2  gate1081(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1082(.a(s_76), .O(gate41inter3));
  inv1  gate1083(.a(s_77), .O(gate41inter4));
  nand2 gate1084(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1085(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1086(.a(G1), .O(gate41inter7));
  inv1  gate1087(.a(G266), .O(gate41inter8));
  nand2 gate1088(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1089(.a(s_77), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1090(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1091(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1092(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate743(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate744(.a(gate43inter0), .b(s_28), .O(gate43inter1));
  and2  gate745(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate746(.a(s_28), .O(gate43inter3));
  inv1  gate747(.a(s_29), .O(gate43inter4));
  nand2 gate748(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate749(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate750(.a(G3), .O(gate43inter7));
  inv1  gate751(.a(G269), .O(gate43inter8));
  nand2 gate752(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate753(.a(s_29), .b(gate43inter3), .O(gate43inter10));
  nor2  gate754(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate755(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate756(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1387(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1388(.a(gate44inter0), .b(s_120), .O(gate44inter1));
  and2  gate1389(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1390(.a(s_120), .O(gate44inter3));
  inv1  gate1391(.a(s_121), .O(gate44inter4));
  nand2 gate1392(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1393(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1394(.a(G4), .O(gate44inter7));
  inv1  gate1395(.a(G269), .O(gate44inter8));
  nand2 gate1396(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1397(.a(s_121), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1398(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1399(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1400(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate547(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate548(.a(gate45inter0), .b(s_0), .O(gate45inter1));
  and2  gate549(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate550(.a(s_0), .O(gate45inter3));
  inv1  gate551(.a(s_1), .O(gate45inter4));
  nand2 gate552(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate553(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate554(.a(G5), .O(gate45inter7));
  inv1  gate555(.a(G272), .O(gate45inter8));
  nand2 gate556(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate557(.a(s_1), .b(gate45inter3), .O(gate45inter10));
  nor2  gate558(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate559(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate560(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1317(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1318(.a(gate53inter0), .b(s_110), .O(gate53inter1));
  and2  gate1319(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1320(.a(s_110), .O(gate53inter3));
  inv1  gate1321(.a(s_111), .O(gate53inter4));
  nand2 gate1322(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1323(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1324(.a(G13), .O(gate53inter7));
  inv1  gate1325(.a(G284), .O(gate53inter8));
  nand2 gate1326(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1327(.a(s_111), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1328(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1329(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1330(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1093(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1094(.a(gate58inter0), .b(s_78), .O(gate58inter1));
  and2  gate1095(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1096(.a(s_78), .O(gate58inter3));
  inv1  gate1097(.a(s_79), .O(gate58inter4));
  nand2 gate1098(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1099(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1100(.a(G18), .O(gate58inter7));
  inv1  gate1101(.a(G290), .O(gate58inter8));
  nand2 gate1102(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1103(.a(s_79), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1104(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1105(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1106(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate687(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate688(.a(gate62inter0), .b(s_20), .O(gate62inter1));
  and2  gate689(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate690(.a(s_20), .O(gate62inter3));
  inv1  gate691(.a(s_21), .O(gate62inter4));
  nand2 gate692(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate693(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate694(.a(G22), .O(gate62inter7));
  inv1  gate695(.a(G296), .O(gate62inter8));
  nand2 gate696(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate697(.a(s_21), .b(gate62inter3), .O(gate62inter10));
  nor2  gate698(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate699(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate700(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1289(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1290(.a(gate64inter0), .b(s_106), .O(gate64inter1));
  and2  gate1291(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1292(.a(s_106), .O(gate64inter3));
  inv1  gate1293(.a(s_107), .O(gate64inter4));
  nand2 gate1294(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1295(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1296(.a(G24), .O(gate64inter7));
  inv1  gate1297(.a(G299), .O(gate64inter8));
  nand2 gate1298(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1299(.a(s_107), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1300(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1301(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1302(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate953(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate954(.a(gate66inter0), .b(s_58), .O(gate66inter1));
  and2  gate955(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate956(.a(s_58), .O(gate66inter3));
  inv1  gate957(.a(s_59), .O(gate66inter4));
  nand2 gate958(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate959(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate960(.a(G26), .O(gate66inter7));
  inv1  gate961(.a(G302), .O(gate66inter8));
  nand2 gate962(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate963(.a(s_59), .b(gate66inter3), .O(gate66inter10));
  nor2  gate964(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate965(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate966(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1401(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1402(.a(gate68inter0), .b(s_122), .O(gate68inter1));
  and2  gate1403(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1404(.a(s_122), .O(gate68inter3));
  inv1  gate1405(.a(s_123), .O(gate68inter4));
  nand2 gate1406(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1407(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1408(.a(G28), .O(gate68inter7));
  inv1  gate1409(.a(G305), .O(gate68inter8));
  nand2 gate1410(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1411(.a(s_123), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1412(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1413(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1414(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1541(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1542(.a(gate71inter0), .b(s_142), .O(gate71inter1));
  and2  gate1543(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1544(.a(s_142), .O(gate71inter3));
  inv1  gate1545(.a(s_143), .O(gate71inter4));
  nand2 gate1546(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1547(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1548(.a(G31), .O(gate71inter7));
  inv1  gate1549(.a(G311), .O(gate71inter8));
  nand2 gate1550(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1551(.a(s_143), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1552(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1553(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1554(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1457(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1458(.a(gate74inter0), .b(s_130), .O(gate74inter1));
  and2  gate1459(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1460(.a(s_130), .O(gate74inter3));
  inv1  gate1461(.a(s_131), .O(gate74inter4));
  nand2 gate1462(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1463(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1464(.a(G5), .O(gate74inter7));
  inv1  gate1465(.a(G314), .O(gate74inter8));
  nand2 gate1466(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1467(.a(s_131), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1468(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1469(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1470(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate981(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate982(.a(gate79inter0), .b(s_62), .O(gate79inter1));
  and2  gate983(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate984(.a(s_62), .O(gate79inter3));
  inv1  gate985(.a(s_63), .O(gate79inter4));
  nand2 gate986(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate987(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate988(.a(G10), .O(gate79inter7));
  inv1  gate989(.a(G323), .O(gate79inter8));
  nand2 gate990(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate991(.a(s_63), .b(gate79inter3), .O(gate79inter10));
  nor2  gate992(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate993(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate994(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate673(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate674(.a(gate81inter0), .b(s_18), .O(gate81inter1));
  and2  gate675(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate676(.a(s_18), .O(gate81inter3));
  inv1  gate677(.a(s_19), .O(gate81inter4));
  nand2 gate678(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate679(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate680(.a(G3), .O(gate81inter7));
  inv1  gate681(.a(G326), .O(gate81inter8));
  nand2 gate682(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate683(.a(s_19), .b(gate81inter3), .O(gate81inter10));
  nor2  gate684(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate685(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate686(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1779(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1780(.a(gate93inter0), .b(s_176), .O(gate93inter1));
  and2  gate1781(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1782(.a(s_176), .O(gate93inter3));
  inv1  gate1783(.a(s_177), .O(gate93inter4));
  nand2 gate1784(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1785(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1786(.a(G18), .O(gate93inter7));
  inv1  gate1787(.a(G344), .O(gate93inter8));
  nand2 gate1788(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1789(.a(s_177), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1790(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1791(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1792(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1163(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1164(.a(gate106inter0), .b(s_88), .O(gate106inter1));
  and2  gate1165(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1166(.a(s_88), .O(gate106inter3));
  inv1  gate1167(.a(s_89), .O(gate106inter4));
  nand2 gate1168(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1169(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1170(.a(G364), .O(gate106inter7));
  inv1  gate1171(.a(G365), .O(gate106inter8));
  nand2 gate1172(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1173(.a(s_89), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1174(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1175(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1176(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1611(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1612(.a(gate107inter0), .b(s_152), .O(gate107inter1));
  and2  gate1613(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1614(.a(s_152), .O(gate107inter3));
  inv1  gate1615(.a(s_153), .O(gate107inter4));
  nand2 gate1616(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1617(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1618(.a(G366), .O(gate107inter7));
  inv1  gate1619(.a(G367), .O(gate107inter8));
  nand2 gate1620(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1621(.a(s_153), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1622(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1623(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1624(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1989(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1990(.a(gate110inter0), .b(s_206), .O(gate110inter1));
  and2  gate1991(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1992(.a(s_206), .O(gate110inter3));
  inv1  gate1993(.a(s_207), .O(gate110inter4));
  nand2 gate1994(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1995(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1996(.a(G372), .O(gate110inter7));
  inv1  gate1997(.a(G373), .O(gate110inter8));
  nand2 gate1998(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1999(.a(s_207), .b(gate110inter3), .O(gate110inter10));
  nor2  gate2000(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate2001(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate2002(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate855(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate856(.a(gate112inter0), .b(s_44), .O(gate112inter1));
  and2  gate857(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate858(.a(s_44), .O(gate112inter3));
  inv1  gate859(.a(s_45), .O(gate112inter4));
  nand2 gate860(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate861(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate862(.a(G376), .O(gate112inter7));
  inv1  gate863(.a(G377), .O(gate112inter8));
  nand2 gate864(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate865(.a(s_45), .b(gate112inter3), .O(gate112inter10));
  nor2  gate866(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate867(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate868(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1681(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1682(.a(gate116inter0), .b(s_162), .O(gate116inter1));
  and2  gate1683(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1684(.a(s_162), .O(gate116inter3));
  inv1  gate1685(.a(s_163), .O(gate116inter4));
  nand2 gate1686(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1687(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1688(.a(G384), .O(gate116inter7));
  inv1  gate1689(.a(G385), .O(gate116inter8));
  nand2 gate1690(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1691(.a(s_163), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1692(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1693(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1694(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate1821(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1822(.a(gate117inter0), .b(s_182), .O(gate117inter1));
  and2  gate1823(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1824(.a(s_182), .O(gate117inter3));
  inv1  gate1825(.a(s_183), .O(gate117inter4));
  nand2 gate1826(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1827(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1828(.a(G386), .O(gate117inter7));
  inv1  gate1829(.a(G387), .O(gate117inter8));
  nand2 gate1830(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1831(.a(s_183), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1832(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1833(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1834(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate603(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate604(.a(gate124inter0), .b(s_8), .O(gate124inter1));
  and2  gate605(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate606(.a(s_8), .O(gate124inter3));
  inv1  gate607(.a(s_9), .O(gate124inter4));
  nand2 gate608(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate609(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate610(.a(G400), .O(gate124inter7));
  inv1  gate611(.a(G401), .O(gate124inter8));
  nand2 gate612(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate613(.a(s_9), .b(gate124inter3), .O(gate124inter10));
  nor2  gate614(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate615(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate616(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1331(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1332(.a(gate127inter0), .b(s_112), .O(gate127inter1));
  and2  gate1333(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1334(.a(s_112), .O(gate127inter3));
  inv1  gate1335(.a(s_113), .O(gate127inter4));
  nand2 gate1336(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1337(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1338(.a(G406), .O(gate127inter7));
  inv1  gate1339(.a(G407), .O(gate127inter8));
  nand2 gate1340(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1341(.a(s_113), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1342(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1343(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1344(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1219(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1220(.a(gate137inter0), .b(s_96), .O(gate137inter1));
  and2  gate1221(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1222(.a(s_96), .O(gate137inter3));
  inv1  gate1223(.a(s_97), .O(gate137inter4));
  nand2 gate1224(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1225(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1226(.a(G426), .O(gate137inter7));
  inv1  gate1227(.a(G429), .O(gate137inter8));
  nand2 gate1228(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1229(.a(s_97), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1230(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1231(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1232(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate2073(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2074(.a(gate138inter0), .b(s_218), .O(gate138inter1));
  and2  gate2075(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2076(.a(s_218), .O(gate138inter3));
  inv1  gate2077(.a(s_219), .O(gate138inter4));
  nand2 gate2078(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2079(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2080(.a(G432), .O(gate138inter7));
  inv1  gate2081(.a(G435), .O(gate138inter8));
  nand2 gate2082(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2083(.a(s_219), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2084(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2085(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2086(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate659(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate660(.a(gate147inter0), .b(s_16), .O(gate147inter1));
  and2  gate661(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate662(.a(s_16), .O(gate147inter3));
  inv1  gate663(.a(s_17), .O(gate147inter4));
  nand2 gate664(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate665(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate666(.a(G486), .O(gate147inter7));
  inv1  gate667(.a(G489), .O(gate147inter8));
  nand2 gate668(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate669(.a(s_17), .b(gate147inter3), .O(gate147inter10));
  nor2  gate670(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate671(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate672(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1037(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1038(.a(gate150inter0), .b(s_70), .O(gate150inter1));
  and2  gate1039(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1040(.a(s_70), .O(gate150inter3));
  inv1  gate1041(.a(s_71), .O(gate150inter4));
  nand2 gate1042(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1043(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1044(.a(G504), .O(gate150inter7));
  inv1  gate1045(.a(G507), .O(gate150inter8));
  nand2 gate1046(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1047(.a(s_71), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1048(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1049(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1050(.a(gate150inter12), .b(gate150inter1), .O(G561));

  xor2  gate897(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate898(.a(gate151inter0), .b(s_50), .O(gate151inter1));
  and2  gate899(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate900(.a(s_50), .O(gate151inter3));
  inv1  gate901(.a(s_51), .O(gate151inter4));
  nand2 gate902(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate903(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate904(.a(G510), .O(gate151inter7));
  inv1  gate905(.a(G513), .O(gate151inter8));
  nand2 gate906(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate907(.a(s_51), .b(gate151inter3), .O(gate151inter10));
  nor2  gate908(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate909(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate910(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate575(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate576(.a(gate155inter0), .b(s_4), .O(gate155inter1));
  and2  gate577(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate578(.a(s_4), .O(gate155inter3));
  inv1  gate579(.a(s_5), .O(gate155inter4));
  nand2 gate580(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate581(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate582(.a(G432), .O(gate155inter7));
  inv1  gate583(.a(G525), .O(gate155inter8));
  nand2 gate584(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate585(.a(s_5), .b(gate155inter3), .O(gate155inter10));
  nor2  gate586(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate587(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate588(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate2087(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate2088(.a(gate156inter0), .b(s_220), .O(gate156inter1));
  and2  gate2089(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate2090(.a(s_220), .O(gate156inter3));
  inv1  gate2091(.a(s_221), .O(gate156inter4));
  nand2 gate2092(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate2093(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate2094(.a(G435), .O(gate156inter7));
  inv1  gate2095(.a(G525), .O(gate156inter8));
  nand2 gate2096(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate2097(.a(s_221), .b(gate156inter3), .O(gate156inter10));
  nor2  gate2098(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate2099(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate2100(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate939(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate940(.a(gate159inter0), .b(s_56), .O(gate159inter1));
  and2  gate941(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate942(.a(s_56), .O(gate159inter3));
  inv1  gate943(.a(s_57), .O(gate159inter4));
  nand2 gate944(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate945(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate946(.a(G444), .O(gate159inter7));
  inv1  gate947(.a(G531), .O(gate159inter8));
  nand2 gate948(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate949(.a(s_57), .b(gate159inter3), .O(gate159inter10));
  nor2  gate950(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate951(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate952(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2045(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2046(.a(gate160inter0), .b(s_214), .O(gate160inter1));
  and2  gate2047(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2048(.a(s_214), .O(gate160inter3));
  inv1  gate2049(.a(s_215), .O(gate160inter4));
  nand2 gate2050(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2051(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2052(.a(G447), .O(gate160inter7));
  inv1  gate2053(.a(G531), .O(gate160inter8));
  nand2 gate2054(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2055(.a(s_215), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2056(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2057(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2058(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1877(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1878(.a(gate165inter0), .b(s_190), .O(gate165inter1));
  and2  gate1879(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1880(.a(s_190), .O(gate165inter3));
  inv1  gate1881(.a(s_191), .O(gate165inter4));
  nand2 gate1882(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1883(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1884(.a(G462), .O(gate165inter7));
  inv1  gate1885(.a(G540), .O(gate165inter8));
  nand2 gate1886(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1887(.a(s_191), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1888(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1889(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1890(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1485(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1486(.a(gate170inter0), .b(s_134), .O(gate170inter1));
  and2  gate1487(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1488(.a(s_134), .O(gate170inter3));
  inv1  gate1489(.a(s_135), .O(gate170inter4));
  nand2 gate1490(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1491(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1492(.a(G477), .O(gate170inter7));
  inv1  gate1493(.a(G546), .O(gate170inter8));
  nand2 gate1494(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1495(.a(s_135), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1496(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1497(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1498(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1107(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1108(.a(gate176inter0), .b(s_80), .O(gate176inter1));
  and2  gate1109(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1110(.a(s_80), .O(gate176inter3));
  inv1  gate1111(.a(s_81), .O(gate176inter4));
  nand2 gate1112(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1113(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1114(.a(G495), .O(gate176inter7));
  inv1  gate1115(.a(G555), .O(gate176inter8));
  nand2 gate1116(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1117(.a(s_81), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1118(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1119(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1120(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1807(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1808(.a(gate183inter0), .b(s_180), .O(gate183inter1));
  and2  gate1809(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1810(.a(s_180), .O(gate183inter3));
  inv1  gate1811(.a(s_181), .O(gate183inter4));
  nand2 gate1812(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1813(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1814(.a(G516), .O(gate183inter7));
  inv1  gate1815(.a(G567), .O(gate183inter8));
  nand2 gate1816(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1817(.a(s_181), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1818(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1819(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1820(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1051(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1052(.a(gate187inter0), .b(s_72), .O(gate187inter1));
  and2  gate1053(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1054(.a(s_72), .O(gate187inter3));
  inv1  gate1055(.a(s_73), .O(gate187inter4));
  nand2 gate1056(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1057(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1058(.a(G574), .O(gate187inter7));
  inv1  gate1059(.a(G575), .O(gate187inter8));
  nand2 gate1060(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1061(.a(s_73), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1062(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1063(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1064(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1177(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1178(.a(gate189inter0), .b(s_90), .O(gate189inter1));
  and2  gate1179(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1180(.a(s_90), .O(gate189inter3));
  inv1  gate1181(.a(s_91), .O(gate189inter4));
  nand2 gate1182(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1183(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1184(.a(G578), .O(gate189inter7));
  inv1  gate1185(.a(G579), .O(gate189inter8));
  nand2 gate1186(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1187(.a(s_91), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1188(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1189(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1190(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1919(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1920(.a(gate190inter0), .b(s_196), .O(gate190inter1));
  and2  gate1921(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1922(.a(s_196), .O(gate190inter3));
  inv1  gate1923(.a(s_197), .O(gate190inter4));
  nand2 gate1924(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1925(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1926(.a(G580), .O(gate190inter7));
  inv1  gate1927(.a(G581), .O(gate190inter8));
  nand2 gate1928(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1929(.a(s_197), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1930(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1931(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1932(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate813(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate814(.a(gate192inter0), .b(s_38), .O(gate192inter1));
  and2  gate815(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate816(.a(s_38), .O(gate192inter3));
  inv1  gate817(.a(s_39), .O(gate192inter4));
  nand2 gate818(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate819(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate820(.a(G584), .O(gate192inter7));
  inv1  gate821(.a(G585), .O(gate192inter8));
  nand2 gate822(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate823(.a(s_39), .b(gate192inter3), .O(gate192inter10));
  nor2  gate824(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate825(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate826(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate925(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate926(.a(gate196inter0), .b(s_54), .O(gate196inter1));
  and2  gate927(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate928(.a(s_54), .O(gate196inter3));
  inv1  gate929(.a(s_55), .O(gate196inter4));
  nand2 gate930(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate931(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate932(.a(G592), .O(gate196inter7));
  inv1  gate933(.a(G593), .O(gate196inter8));
  nand2 gate934(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate935(.a(s_55), .b(gate196inter3), .O(gate196inter10));
  nor2  gate936(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate937(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate938(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1639(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1640(.a(gate201inter0), .b(s_156), .O(gate201inter1));
  and2  gate1641(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1642(.a(s_156), .O(gate201inter3));
  inv1  gate1643(.a(s_157), .O(gate201inter4));
  nand2 gate1644(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1645(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1646(.a(G602), .O(gate201inter7));
  inv1  gate1647(.a(G607), .O(gate201inter8));
  nand2 gate1648(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1649(.a(s_157), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1650(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1651(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1652(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate617(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate618(.a(gate202inter0), .b(s_10), .O(gate202inter1));
  and2  gate619(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate620(.a(s_10), .O(gate202inter3));
  inv1  gate621(.a(s_11), .O(gate202inter4));
  nand2 gate622(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate623(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate624(.a(G612), .O(gate202inter7));
  inv1  gate625(.a(G617), .O(gate202inter8));
  nand2 gate626(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate627(.a(s_11), .b(gate202inter3), .O(gate202inter10));
  nor2  gate628(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate629(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate630(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1751(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1752(.a(gate209inter0), .b(s_172), .O(gate209inter1));
  and2  gate1753(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1754(.a(s_172), .O(gate209inter3));
  inv1  gate1755(.a(s_173), .O(gate209inter4));
  nand2 gate1756(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1757(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1758(.a(G602), .O(gate209inter7));
  inv1  gate1759(.a(G666), .O(gate209inter8));
  nand2 gate1760(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1761(.a(s_173), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1762(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1763(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1764(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1597(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1598(.a(gate212inter0), .b(s_150), .O(gate212inter1));
  and2  gate1599(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1600(.a(s_150), .O(gate212inter3));
  inv1  gate1601(.a(s_151), .O(gate212inter4));
  nand2 gate1602(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1603(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1604(.a(G617), .O(gate212inter7));
  inv1  gate1605(.a(G669), .O(gate212inter8));
  nand2 gate1606(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1607(.a(s_151), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1608(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1609(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1610(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate827(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate828(.a(gate223inter0), .b(s_40), .O(gate223inter1));
  and2  gate829(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate830(.a(s_40), .O(gate223inter3));
  inv1  gate831(.a(s_41), .O(gate223inter4));
  nand2 gate832(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate833(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate834(.a(G627), .O(gate223inter7));
  inv1  gate835(.a(G687), .O(gate223inter8));
  nand2 gate836(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate837(.a(s_41), .b(gate223inter3), .O(gate223inter10));
  nor2  gate838(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate839(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate840(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate561(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate562(.a(gate227inter0), .b(s_2), .O(gate227inter1));
  and2  gate563(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate564(.a(s_2), .O(gate227inter3));
  inv1  gate565(.a(s_3), .O(gate227inter4));
  nand2 gate566(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate567(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate568(.a(G694), .O(gate227inter7));
  inv1  gate569(.a(G695), .O(gate227inter8));
  nand2 gate570(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate571(.a(s_3), .b(gate227inter3), .O(gate227inter10));
  nor2  gate572(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate573(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate574(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate799(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate800(.a(gate228inter0), .b(s_36), .O(gate228inter1));
  and2  gate801(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate802(.a(s_36), .O(gate228inter3));
  inv1  gate803(.a(s_37), .O(gate228inter4));
  nand2 gate804(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate805(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate806(.a(G696), .O(gate228inter7));
  inv1  gate807(.a(G697), .O(gate228inter8));
  nand2 gate808(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate809(.a(s_37), .b(gate228inter3), .O(gate228inter10));
  nor2  gate810(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate811(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate812(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1443(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1444(.a(gate232inter0), .b(s_128), .O(gate232inter1));
  and2  gate1445(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1446(.a(s_128), .O(gate232inter3));
  inv1  gate1447(.a(s_129), .O(gate232inter4));
  nand2 gate1448(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1449(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1450(.a(G704), .O(gate232inter7));
  inv1  gate1451(.a(G705), .O(gate232inter8));
  nand2 gate1452(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1453(.a(s_129), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1454(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1455(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1456(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate1737(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1738(.a(gate233inter0), .b(s_170), .O(gate233inter1));
  and2  gate1739(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1740(.a(s_170), .O(gate233inter3));
  inv1  gate1741(.a(s_171), .O(gate233inter4));
  nand2 gate1742(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1743(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1744(.a(G242), .O(gate233inter7));
  inv1  gate1745(.a(G718), .O(gate233inter8));
  nand2 gate1746(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1747(.a(s_171), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1748(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1749(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1750(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1667(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1668(.a(gate238inter0), .b(s_160), .O(gate238inter1));
  and2  gate1669(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1670(.a(s_160), .O(gate238inter3));
  inv1  gate1671(.a(s_161), .O(gate238inter4));
  nand2 gate1672(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1673(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1674(.a(G257), .O(gate238inter7));
  inv1  gate1675(.a(G709), .O(gate238inter8));
  nand2 gate1676(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1677(.a(s_161), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1678(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1679(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1680(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1023(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1024(.a(gate239inter0), .b(s_68), .O(gate239inter1));
  and2  gate1025(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1026(.a(s_68), .O(gate239inter3));
  inv1  gate1027(.a(s_69), .O(gate239inter4));
  nand2 gate1028(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1029(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1030(.a(G260), .O(gate239inter7));
  inv1  gate1031(.a(G712), .O(gate239inter8));
  nand2 gate1032(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1033(.a(s_69), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1034(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1035(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1036(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate1905(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1906(.a(gate240inter0), .b(s_194), .O(gate240inter1));
  and2  gate1907(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1908(.a(s_194), .O(gate240inter3));
  inv1  gate1909(.a(s_195), .O(gate240inter4));
  nand2 gate1910(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1911(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1912(.a(G263), .O(gate240inter7));
  inv1  gate1913(.a(G715), .O(gate240inter8));
  nand2 gate1914(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1915(.a(s_195), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1916(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1917(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1918(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1975(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1976(.a(gate242inter0), .b(s_204), .O(gate242inter1));
  and2  gate1977(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1978(.a(s_204), .O(gate242inter3));
  inv1  gate1979(.a(s_205), .O(gate242inter4));
  nand2 gate1980(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1981(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1982(.a(G718), .O(gate242inter7));
  inv1  gate1983(.a(G730), .O(gate242inter8));
  nand2 gate1984(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1985(.a(s_205), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1986(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1987(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1988(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1415(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1416(.a(gate243inter0), .b(s_124), .O(gate243inter1));
  and2  gate1417(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1418(.a(s_124), .O(gate243inter3));
  inv1  gate1419(.a(s_125), .O(gate243inter4));
  nand2 gate1420(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1421(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1422(.a(G245), .O(gate243inter7));
  inv1  gate1423(.a(G733), .O(gate243inter8));
  nand2 gate1424(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1425(.a(s_125), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1426(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1427(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1428(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1933(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1934(.a(gate244inter0), .b(s_198), .O(gate244inter1));
  and2  gate1935(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1936(.a(s_198), .O(gate244inter3));
  inv1  gate1937(.a(s_199), .O(gate244inter4));
  nand2 gate1938(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1939(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1940(.a(G721), .O(gate244inter7));
  inv1  gate1941(.a(G733), .O(gate244inter8));
  nand2 gate1942(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1943(.a(s_199), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1944(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1945(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1946(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1149(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1150(.a(gate250inter0), .b(s_86), .O(gate250inter1));
  and2  gate1151(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1152(.a(s_86), .O(gate250inter3));
  inv1  gate1153(.a(s_87), .O(gate250inter4));
  nand2 gate1154(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1155(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1156(.a(G706), .O(gate250inter7));
  inv1  gate1157(.a(G742), .O(gate250inter8));
  nand2 gate1158(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1159(.a(s_87), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1160(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1161(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1162(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2031(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2032(.a(gate253inter0), .b(s_212), .O(gate253inter1));
  and2  gate2033(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2034(.a(s_212), .O(gate253inter3));
  inv1  gate2035(.a(s_213), .O(gate253inter4));
  nand2 gate2036(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2037(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2038(.a(G260), .O(gate253inter7));
  inv1  gate2039(.a(G748), .O(gate253inter8));
  nand2 gate2040(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2041(.a(s_213), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2042(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2043(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2044(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2059(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2060(.a(gate256inter0), .b(s_216), .O(gate256inter1));
  and2  gate2061(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2062(.a(s_216), .O(gate256inter3));
  inv1  gate2063(.a(s_217), .O(gate256inter4));
  nand2 gate2064(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2065(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2066(.a(G715), .O(gate256inter7));
  inv1  gate2067(.a(G751), .O(gate256inter8));
  nand2 gate2068(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2069(.a(s_217), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2070(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2071(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2072(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1303(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1304(.a(gate260inter0), .b(s_108), .O(gate260inter1));
  and2  gate1305(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1306(.a(s_108), .O(gate260inter3));
  inv1  gate1307(.a(s_109), .O(gate260inter4));
  nand2 gate1308(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1309(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1310(.a(G760), .O(gate260inter7));
  inv1  gate1311(.a(G761), .O(gate260inter8));
  nand2 gate1312(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1313(.a(s_109), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1314(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1315(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1316(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1527(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1528(.a(gate267inter0), .b(s_140), .O(gate267inter1));
  and2  gate1529(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1530(.a(s_140), .O(gate267inter3));
  inv1  gate1531(.a(s_141), .O(gate267inter4));
  nand2 gate1532(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1533(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1534(.a(G648), .O(gate267inter7));
  inv1  gate1535(.a(G776), .O(gate267inter8));
  nand2 gate1536(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1537(.a(s_141), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1538(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1539(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1540(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate701(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate702(.a(gate268inter0), .b(s_22), .O(gate268inter1));
  and2  gate703(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate704(.a(s_22), .O(gate268inter3));
  inv1  gate705(.a(s_23), .O(gate268inter4));
  nand2 gate706(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate707(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate708(.a(G651), .O(gate268inter7));
  inv1  gate709(.a(G779), .O(gate268inter8));
  nand2 gate710(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate711(.a(s_23), .b(gate268inter3), .O(gate268inter10));
  nor2  gate712(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate713(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate714(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1555(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1556(.a(gate271inter0), .b(s_144), .O(gate271inter1));
  and2  gate1557(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1558(.a(s_144), .O(gate271inter3));
  inv1  gate1559(.a(s_145), .O(gate271inter4));
  nand2 gate1560(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1561(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1562(.a(G660), .O(gate271inter7));
  inv1  gate1563(.a(G788), .O(gate271inter8));
  nand2 gate1564(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1565(.a(s_145), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1566(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1567(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1568(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1233(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1234(.a(gate273inter0), .b(s_98), .O(gate273inter1));
  and2  gate1235(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1236(.a(s_98), .O(gate273inter3));
  inv1  gate1237(.a(s_99), .O(gate273inter4));
  nand2 gate1238(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1239(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1240(.a(G642), .O(gate273inter7));
  inv1  gate1241(.a(G794), .O(gate273inter8));
  nand2 gate1242(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1243(.a(s_99), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1244(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1245(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1246(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate883(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate884(.a(gate274inter0), .b(s_48), .O(gate274inter1));
  and2  gate885(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate886(.a(s_48), .O(gate274inter3));
  inv1  gate887(.a(s_49), .O(gate274inter4));
  nand2 gate888(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate889(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate890(.a(G770), .O(gate274inter7));
  inv1  gate891(.a(G794), .O(gate274inter8));
  nand2 gate892(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate893(.a(s_49), .b(gate274inter3), .O(gate274inter10));
  nor2  gate894(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate895(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate896(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate967(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate968(.a(gate276inter0), .b(s_60), .O(gate276inter1));
  and2  gate969(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate970(.a(s_60), .O(gate276inter3));
  inv1  gate971(.a(s_61), .O(gate276inter4));
  nand2 gate972(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate973(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate974(.a(G773), .O(gate276inter7));
  inv1  gate975(.a(G797), .O(gate276inter8));
  nand2 gate976(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate977(.a(s_61), .b(gate276inter3), .O(gate276inter10));
  nor2  gate978(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate979(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate980(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1625(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1626(.a(gate282inter0), .b(s_154), .O(gate282inter1));
  and2  gate1627(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1628(.a(s_154), .O(gate282inter3));
  inv1  gate1629(.a(s_155), .O(gate282inter4));
  nand2 gate1630(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1631(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1632(.a(G782), .O(gate282inter7));
  inv1  gate1633(.a(G806), .O(gate282inter8));
  nand2 gate1634(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1635(.a(s_155), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1636(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1637(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1638(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1513(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1514(.a(gate289inter0), .b(s_138), .O(gate289inter1));
  and2  gate1515(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1516(.a(s_138), .O(gate289inter3));
  inv1  gate1517(.a(s_139), .O(gate289inter4));
  nand2 gate1518(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1519(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1520(.a(G818), .O(gate289inter7));
  inv1  gate1521(.a(G819), .O(gate289inter8));
  nand2 gate1522(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1523(.a(s_139), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1524(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1525(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1526(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate715(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate716(.a(gate388inter0), .b(s_24), .O(gate388inter1));
  and2  gate717(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate718(.a(s_24), .O(gate388inter3));
  inv1  gate719(.a(s_25), .O(gate388inter4));
  nand2 gate720(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate721(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate722(.a(G2), .O(gate388inter7));
  inv1  gate723(.a(G1039), .O(gate388inter8));
  nand2 gate724(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate725(.a(s_25), .b(gate388inter3), .O(gate388inter10));
  nor2  gate726(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate727(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate728(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1695(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1696(.a(gate395inter0), .b(s_164), .O(gate395inter1));
  and2  gate1697(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1698(.a(s_164), .O(gate395inter3));
  inv1  gate1699(.a(s_165), .O(gate395inter4));
  nand2 gate1700(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1701(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1702(.a(G9), .O(gate395inter7));
  inv1  gate1703(.a(G1060), .O(gate395inter8));
  nand2 gate1704(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1705(.a(s_165), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1706(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1707(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1708(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate757(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate758(.a(gate398inter0), .b(s_30), .O(gate398inter1));
  and2  gate759(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate760(.a(s_30), .O(gate398inter3));
  inv1  gate761(.a(s_31), .O(gate398inter4));
  nand2 gate762(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate763(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate764(.a(G12), .O(gate398inter7));
  inv1  gate765(.a(G1069), .O(gate398inter8));
  nand2 gate766(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate767(.a(s_31), .b(gate398inter3), .O(gate398inter10));
  nor2  gate768(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate769(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate770(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate869(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate870(.a(gate403inter0), .b(s_46), .O(gate403inter1));
  and2  gate871(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate872(.a(s_46), .O(gate403inter3));
  inv1  gate873(.a(s_47), .O(gate403inter4));
  nand2 gate874(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate875(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate876(.a(G17), .O(gate403inter7));
  inv1  gate877(.a(G1084), .O(gate403inter8));
  nand2 gate878(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate879(.a(s_47), .b(gate403inter3), .O(gate403inter10));
  nor2  gate880(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate881(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate882(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate645(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate646(.a(gate411inter0), .b(s_14), .O(gate411inter1));
  and2  gate647(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate648(.a(s_14), .O(gate411inter3));
  inv1  gate649(.a(s_15), .O(gate411inter4));
  nand2 gate650(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate651(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate652(.a(G25), .O(gate411inter7));
  inv1  gate653(.a(G1108), .O(gate411inter8));
  nand2 gate654(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate655(.a(s_15), .b(gate411inter3), .O(gate411inter10));
  nor2  gate656(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate657(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate658(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1135(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1136(.a(gate412inter0), .b(s_84), .O(gate412inter1));
  and2  gate1137(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1138(.a(s_84), .O(gate412inter3));
  inv1  gate1139(.a(s_85), .O(gate412inter4));
  nand2 gate1140(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1141(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1142(.a(G26), .O(gate412inter7));
  inv1  gate1143(.a(G1111), .O(gate412inter8));
  nand2 gate1144(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1145(.a(s_85), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1146(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1147(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1148(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate729(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate730(.a(gate417inter0), .b(s_26), .O(gate417inter1));
  and2  gate731(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate732(.a(s_26), .O(gate417inter3));
  inv1  gate733(.a(s_27), .O(gate417inter4));
  nand2 gate734(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate735(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate736(.a(G31), .O(gate417inter7));
  inv1  gate737(.a(G1126), .O(gate417inter8));
  nand2 gate738(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate739(.a(s_27), .b(gate417inter3), .O(gate417inter10));
  nor2  gate740(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate741(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate742(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1429(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1430(.a(gate418inter0), .b(s_126), .O(gate418inter1));
  and2  gate1431(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1432(.a(s_126), .O(gate418inter3));
  inv1  gate1433(.a(s_127), .O(gate418inter4));
  nand2 gate1434(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1435(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1436(.a(G32), .O(gate418inter7));
  inv1  gate1437(.a(G1129), .O(gate418inter8));
  nand2 gate1438(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1439(.a(s_127), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1440(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1441(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1442(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1863(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1864(.a(gate419inter0), .b(s_188), .O(gate419inter1));
  and2  gate1865(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1866(.a(s_188), .O(gate419inter3));
  inv1  gate1867(.a(s_189), .O(gate419inter4));
  nand2 gate1868(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1869(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1870(.a(G1), .O(gate419inter7));
  inv1  gate1871(.a(G1132), .O(gate419inter8));
  nand2 gate1872(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1873(.a(s_189), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1874(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1875(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1876(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1359(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1360(.a(gate420inter0), .b(s_116), .O(gate420inter1));
  and2  gate1361(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1362(.a(s_116), .O(gate420inter3));
  inv1  gate1363(.a(s_117), .O(gate420inter4));
  nand2 gate1364(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1365(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1366(.a(G1036), .O(gate420inter7));
  inv1  gate1367(.a(G1132), .O(gate420inter8));
  nand2 gate1368(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1369(.a(s_117), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1370(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1371(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1372(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2017(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2018(.a(gate424inter0), .b(s_210), .O(gate424inter1));
  and2  gate2019(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2020(.a(s_210), .O(gate424inter3));
  inv1  gate2021(.a(s_211), .O(gate424inter4));
  nand2 gate2022(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2023(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2024(.a(G1042), .O(gate424inter7));
  inv1  gate2025(.a(G1138), .O(gate424inter8));
  nand2 gate2026(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2027(.a(s_211), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2028(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2029(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2030(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1009(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1010(.a(gate428inter0), .b(s_66), .O(gate428inter1));
  and2  gate1011(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1012(.a(s_66), .O(gate428inter3));
  inv1  gate1013(.a(s_67), .O(gate428inter4));
  nand2 gate1014(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1015(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1016(.a(G1048), .O(gate428inter7));
  inv1  gate1017(.a(G1144), .O(gate428inter8));
  nand2 gate1018(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1019(.a(s_67), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1020(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1021(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1022(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate995(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate996(.a(gate434inter0), .b(s_64), .O(gate434inter1));
  and2  gate997(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate998(.a(s_64), .O(gate434inter3));
  inv1  gate999(.a(s_65), .O(gate434inter4));
  nand2 gate1000(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1001(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1002(.a(G1057), .O(gate434inter7));
  inv1  gate1003(.a(G1153), .O(gate434inter8));
  nand2 gate1004(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1005(.a(s_65), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1006(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1007(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1008(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1653(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1654(.a(gate435inter0), .b(s_158), .O(gate435inter1));
  and2  gate1655(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1656(.a(s_158), .O(gate435inter3));
  inv1  gate1657(.a(s_159), .O(gate435inter4));
  nand2 gate1658(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1659(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1660(.a(G9), .O(gate435inter7));
  inv1  gate1661(.a(G1156), .O(gate435inter8));
  nand2 gate1662(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1663(.a(s_159), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1664(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1665(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1666(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1205(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1206(.a(gate437inter0), .b(s_94), .O(gate437inter1));
  and2  gate1207(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1208(.a(s_94), .O(gate437inter3));
  inv1  gate1209(.a(s_95), .O(gate437inter4));
  nand2 gate1210(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1211(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1212(.a(G10), .O(gate437inter7));
  inv1  gate1213(.a(G1159), .O(gate437inter8));
  nand2 gate1214(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1215(.a(s_95), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1216(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1217(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1218(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate589(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate590(.a(gate446inter0), .b(s_6), .O(gate446inter1));
  and2  gate591(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate592(.a(s_6), .O(gate446inter3));
  inv1  gate593(.a(s_7), .O(gate446inter4));
  nand2 gate594(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate595(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate596(.a(G1075), .O(gate446inter7));
  inv1  gate597(.a(G1171), .O(gate446inter8));
  nand2 gate598(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate599(.a(s_7), .b(gate446inter3), .O(gate446inter10));
  nor2  gate600(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate601(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate602(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1345(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1346(.a(gate447inter0), .b(s_114), .O(gate447inter1));
  and2  gate1347(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1348(.a(s_114), .O(gate447inter3));
  inv1  gate1349(.a(s_115), .O(gate447inter4));
  nand2 gate1350(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1351(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1352(.a(G15), .O(gate447inter7));
  inv1  gate1353(.a(G1174), .O(gate447inter8));
  nand2 gate1354(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1355(.a(s_115), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1356(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1357(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1358(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1793(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1794(.a(gate448inter0), .b(s_178), .O(gate448inter1));
  and2  gate1795(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1796(.a(s_178), .O(gate448inter3));
  inv1  gate1797(.a(s_179), .O(gate448inter4));
  nand2 gate1798(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1799(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1800(.a(G1078), .O(gate448inter7));
  inv1  gate1801(.a(G1174), .O(gate448inter8));
  nand2 gate1802(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1803(.a(s_179), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1804(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1805(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1806(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1849(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1850(.a(gate451inter0), .b(s_186), .O(gate451inter1));
  and2  gate1851(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1852(.a(s_186), .O(gate451inter3));
  inv1  gate1853(.a(s_187), .O(gate451inter4));
  nand2 gate1854(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1855(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1856(.a(G17), .O(gate451inter7));
  inv1  gate1857(.a(G1180), .O(gate451inter8));
  nand2 gate1858(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1859(.a(s_187), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1860(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1861(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1862(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1261(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1262(.a(gate457inter0), .b(s_102), .O(gate457inter1));
  and2  gate1263(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1264(.a(s_102), .O(gate457inter3));
  inv1  gate1265(.a(s_103), .O(gate457inter4));
  nand2 gate1266(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1267(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1268(.a(G20), .O(gate457inter7));
  inv1  gate1269(.a(G1189), .O(gate457inter8));
  nand2 gate1270(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1271(.a(s_103), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1272(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1273(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1274(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1373(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1374(.a(gate458inter0), .b(s_118), .O(gate458inter1));
  and2  gate1375(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1376(.a(s_118), .O(gate458inter3));
  inv1  gate1377(.a(s_119), .O(gate458inter4));
  nand2 gate1378(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1379(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1380(.a(G1093), .O(gate458inter7));
  inv1  gate1381(.a(G1189), .O(gate458inter8));
  nand2 gate1382(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1383(.a(s_119), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1384(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1385(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1386(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1583(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1584(.a(gate460inter0), .b(s_148), .O(gate460inter1));
  and2  gate1585(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1586(.a(s_148), .O(gate460inter3));
  inv1  gate1587(.a(s_149), .O(gate460inter4));
  nand2 gate1588(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1589(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1590(.a(G1096), .O(gate460inter7));
  inv1  gate1591(.a(G1192), .O(gate460inter8));
  nand2 gate1592(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1593(.a(s_149), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1594(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1595(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1596(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate785(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate786(.a(gate465inter0), .b(s_34), .O(gate465inter1));
  and2  gate787(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate788(.a(s_34), .O(gate465inter3));
  inv1  gate789(.a(s_35), .O(gate465inter4));
  nand2 gate790(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate791(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate792(.a(G24), .O(gate465inter7));
  inv1  gate793(.a(G1201), .O(gate465inter8));
  nand2 gate794(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate795(.a(s_35), .b(gate465inter3), .O(gate465inter10));
  nor2  gate796(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate797(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate798(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1121(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1122(.a(gate477inter0), .b(s_82), .O(gate477inter1));
  and2  gate1123(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1124(.a(s_82), .O(gate477inter3));
  inv1  gate1125(.a(s_83), .O(gate477inter4));
  nand2 gate1126(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1127(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1128(.a(G30), .O(gate477inter7));
  inv1  gate1129(.a(G1219), .O(gate477inter8));
  nand2 gate1130(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1131(.a(s_83), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1132(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1133(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1134(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1499(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1500(.a(gate483inter0), .b(s_136), .O(gate483inter1));
  and2  gate1501(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1502(.a(s_136), .O(gate483inter3));
  inv1  gate1503(.a(s_137), .O(gate483inter4));
  nand2 gate1504(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1505(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1506(.a(G1228), .O(gate483inter7));
  inv1  gate1507(.a(G1229), .O(gate483inter8));
  nand2 gate1508(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1509(.a(s_137), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1510(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1511(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1512(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1709(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1710(.a(gate490inter0), .b(s_166), .O(gate490inter1));
  and2  gate1711(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1712(.a(s_166), .O(gate490inter3));
  inv1  gate1713(.a(s_167), .O(gate490inter4));
  nand2 gate1714(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1715(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1716(.a(G1242), .O(gate490inter7));
  inv1  gate1717(.a(G1243), .O(gate490inter8));
  nand2 gate1718(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1719(.a(s_167), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1720(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1721(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1722(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate841(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate842(.a(gate492inter0), .b(s_42), .O(gate492inter1));
  and2  gate843(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate844(.a(s_42), .O(gate492inter3));
  inv1  gate845(.a(s_43), .O(gate492inter4));
  nand2 gate846(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate847(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate848(.a(G1246), .O(gate492inter7));
  inv1  gate849(.a(G1247), .O(gate492inter8));
  nand2 gate850(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate851(.a(s_43), .b(gate492inter3), .O(gate492inter10));
  nor2  gate852(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate853(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate854(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate911(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate912(.a(gate493inter0), .b(s_52), .O(gate493inter1));
  and2  gate913(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate914(.a(s_52), .O(gate493inter3));
  inv1  gate915(.a(s_53), .O(gate493inter4));
  nand2 gate916(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate917(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate918(.a(G1248), .O(gate493inter7));
  inv1  gate919(.a(G1249), .O(gate493inter8));
  nand2 gate920(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate921(.a(s_53), .b(gate493inter3), .O(gate493inter10));
  nor2  gate922(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate923(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate924(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1569(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1570(.a(gate494inter0), .b(s_146), .O(gate494inter1));
  and2  gate1571(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1572(.a(s_146), .O(gate494inter3));
  inv1  gate1573(.a(s_147), .O(gate494inter4));
  nand2 gate1574(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1575(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1576(.a(G1250), .O(gate494inter7));
  inv1  gate1577(.a(G1251), .O(gate494inter8));
  nand2 gate1578(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1579(.a(s_147), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1580(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1581(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1582(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1835(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1836(.a(gate497inter0), .b(s_184), .O(gate497inter1));
  and2  gate1837(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1838(.a(s_184), .O(gate497inter3));
  inv1  gate1839(.a(s_185), .O(gate497inter4));
  nand2 gate1840(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1841(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1842(.a(G1256), .O(gate497inter7));
  inv1  gate1843(.a(G1257), .O(gate497inter8));
  nand2 gate1844(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1845(.a(s_185), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1846(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1847(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1848(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1891(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1892(.a(gate501inter0), .b(s_192), .O(gate501inter1));
  and2  gate1893(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1894(.a(s_192), .O(gate501inter3));
  inv1  gate1895(.a(s_193), .O(gate501inter4));
  nand2 gate1896(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1897(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1898(.a(G1264), .O(gate501inter7));
  inv1  gate1899(.a(G1265), .O(gate501inter8));
  nand2 gate1900(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1901(.a(s_193), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1902(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1903(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1904(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1765(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1766(.a(gate502inter0), .b(s_174), .O(gate502inter1));
  and2  gate1767(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1768(.a(s_174), .O(gate502inter3));
  inv1  gate1769(.a(s_175), .O(gate502inter4));
  nand2 gate1770(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1771(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1772(.a(G1266), .O(gate502inter7));
  inv1  gate1773(.a(G1267), .O(gate502inter8));
  nand2 gate1774(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1775(.a(s_175), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1776(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1777(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1778(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2003(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2004(.a(gate503inter0), .b(s_208), .O(gate503inter1));
  and2  gate2005(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2006(.a(s_208), .O(gate503inter3));
  inv1  gate2007(.a(s_209), .O(gate503inter4));
  nand2 gate2008(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2009(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2010(.a(G1268), .O(gate503inter7));
  inv1  gate2011(.a(G1269), .O(gate503inter8));
  nand2 gate2012(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2013(.a(s_209), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2014(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2015(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2016(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1471(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1472(.a(gate505inter0), .b(s_132), .O(gate505inter1));
  and2  gate1473(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1474(.a(s_132), .O(gate505inter3));
  inv1  gate1475(.a(s_133), .O(gate505inter4));
  nand2 gate1476(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1477(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1478(.a(G1272), .O(gate505inter7));
  inv1  gate1479(.a(G1273), .O(gate505inter8));
  nand2 gate1480(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1481(.a(s_133), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1482(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1483(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1484(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule