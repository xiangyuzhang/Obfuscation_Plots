module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate1inter0, gate1inter1, gate1inter2, gate1inter3, gate1inter4, gate1inter5, gate1inter6, gate1inter7, gate1inter8, gate1inter9, gate1inter10, gate1inter11, gate1inter12, gate6inter0, gate6inter1, gate6inter2, gate6inter3, gate6inter4, gate6inter5, gate6inter6, gate6inter7, gate6inter8, gate6inter9, gate6inter10, gate6inter11, gate6inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate4inter0, gate4inter1, gate4inter2, gate4inter3, gate4inter4, gate4inter5, gate4inter6, gate4inter7, gate4inter8, gate4inter9, gate4inter10, gate4inter11, gate4inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12;

  xor2  gate329(.a(N5), .b(N1), .O(gate1inter0));
  nand2 gate330(.a(gate1inter0), .b(s_18), .O(gate1inter1));
  and2  gate331(.a(N5), .b(N1), .O(gate1inter2));
  inv1  gate332(.a(s_18), .O(gate1inter3));
  inv1  gate333(.a(s_19), .O(gate1inter4));
  nand2 gate334(.a(gate1inter4), .b(gate1inter3), .O(gate1inter5));
  nor2  gate335(.a(gate1inter5), .b(gate1inter2), .O(gate1inter6));
  inv1  gate336(.a(N1), .O(gate1inter7));
  inv1  gate337(.a(N5), .O(gate1inter8));
  nand2 gate338(.a(gate1inter8), .b(gate1inter7), .O(gate1inter9));
  nand2 gate339(.a(s_19), .b(gate1inter3), .O(gate1inter10));
  nor2  gate340(.a(gate1inter10), .b(gate1inter9), .O(gate1inter11));
  nor2  gate341(.a(gate1inter11), .b(gate1inter6), .O(gate1inter12));
  nand2 gate342(.a(gate1inter12), .b(gate1inter1), .O(N250));
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );

  xor2  gate511(.a(N29), .b(N25), .O(gate4inter0));
  nand2 gate512(.a(gate4inter0), .b(s_44), .O(gate4inter1));
  and2  gate513(.a(N29), .b(N25), .O(gate4inter2));
  inv1  gate514(.a(s_44), .O(gate4inter3));
  inv1  gate515(.a(s_45), .O(gate4inter4));
  nand2 gate516(.a(gate4inter4), .b(gate4inter3), .O(gate4inter5));
  nor2  gate517(.a(gate4inter5), .b(gate4inter2), .O(gate4inter6));
  inv1  gate518(.a(N25), .O(gate4inter7));
  inv1  gate519(.a(N29), .O(gate4inter8));
  nand2 gate520(.a(gate4inter8), .b(gate4inter7), .O(gate4inter9));
  nand2 gate521(.a(s_45), .b(gate4inter3), .O(gate4inter10));
  nor2  gate522(.a(gate4inter10), .b(gate4inter9), .O(gate4inter11));
  nor2  gate523(.a(gate4inter11), .b(gate4inter6), .O(gate4inter12));
  nand2 gate524(.a(gate4inter12), .b(gate4inter1), .O(N253));
xor2 gate5( .a(N33), .b(N37), .O(N254) );

  xor2  gate343(.a(N45), .b(N41), .O(gate6inter0));
  nand2 gate344(.a(gate6inter0), .b(s_20), .O(gate6inter1));
  and2  gate345(.a(N45), .b(N41), .O(gate6inter2));
  inv1  gate346(.a(s_20), .O(gate6inter3));
  inv1  gate347(.a(s_21), .O(gate6inter4));
  nand2 gate348(.a(gate6inter4), .b(gate6inter3), .O(gate6inter5));
  nor2  gate349(.a(gate6inter5), .b(gate6inter2), .O(gate6inter6));
  inv1  gate350(.a(N41), .O(gate6inter7));
  inv1  gate351(.a(N45), .O(gate6inter8));
  nand2 gate352(.a(gate6inter8), .b(gate6inter7), .O(gate6inter9));
  nand2 gate353(.a(s_21), .b(gate6inter3), .O(gate6inter10));
  nor2  gate354(.a(gate6inter10), .b(gate6inter9), .O(gate6inter11));
  nor2  gate355(.a(gate6inter11), .b(gate6inter6), .O(gate6inter12));
  nand2 gate356(.a(gate6inter12), .b(gate6inter1), .O(N255));
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );

  xor2  gate231(.a(N125), .b(N121), .O(gate16inter0));
  nand2 gate232(.a(gate16inter0), .b(s_4), .O(gate16inter1));
  and2  gate233(.a(N125), .b(N121), .O(gate16inter2));
  inv1  gate234(.a(s_4), .O(gate16inter3));
  inv1  gate235(.a(s_5), .O(gate16inter4));
  nand2 gate236(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate237(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate238(.a(N121), .O(gate16inter7));
  inv1  gate239(.a(N125), .O(gate16inter8));
  nand2 gate240(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate241(.a(s_5), .b(gate16inter3), .O(gate16inter10));
  nor2  gate242(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate243(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate244(.a(gate16inter12), .b(gate16inter1), .O(N265));
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate273(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate274(.a(gate25inter0), .b(s_10), .O(gate25inter1));
  and2  gate275(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate276(.a(s_10), .O(gate25inter3));
  inv1  gate277(.a(s_11), .O(gate25inter4));
  nand2 gate278(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate279(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate280(.a(N1), .O(gate25inter7));
  inv1  gate281(.a(N17), .O(gate25inter8));
  nand2 gate282(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate283(.a(s_11), .b(gate25inter3), .O(gate25inter10));
  nor2  gate284(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate285(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate286(.a(gate25inter12), .b(gate25inter1), .O(N274));
xor2 gate26( .a(N33), .b(N49), .O(N275) );

  xor2  gate315(.a(N21), .b(N5), .O(gate27inter0));
  nand2 gate316(.a(gate27inter0), .b(s_16), .O(gate27inter1));
  and2  gate317(.a(N21), .b(N5), .O(gate27inter2));
  inv1  gate318(.a(s_16), .O(gate27inter3));
  inv1  gate319(.a(s_17), .O(gate27inter4));
  nand2 gate320(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate321(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate322(.a(N5), .O(gate27inter7));
  inv1  gate323(.a(N21), .O(gate27inter8));
  nand2 gate324(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate325(.a(s_17), .b(gate27inter3), .O(gate27inter10));
  nor2  gate326(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate327(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate328(.a(gate27inter12), .b(gate27inter1), .O(N276));

  xor2  gate259(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate260(.a(gate28inter0), .b(s_8), .O(gate28inter1));
  and2  gate261(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate262(.a(s_8), .O(gate28inter3));
  inv1  gate263(.a(s_9), .O(gate28inter4));
  nand2 gate264(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate265(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate266(.a(N37), .O(gate28inter7));
  inv1  gate267(.a(N53), .O(gate28inter8));
  nand2 gate268(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate269(.a(s_9), .b(gate28inter3), .O(gate28inter10));
  nor2  gate270(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate271(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate272(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );

  xor2  gate217(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate218(.a(gate40inter0), .b(s_2), .O(gate40inter1));
  and2  gate219(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate220(.a(s_2), .O(gate40inter3));
  inv1  gate221(.a(s_3), .O(gate40inter4));
  nand2 gate222(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate223(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate224(.a(N109), .O(gate40inter7));
  inv1  gate225(.a(N125), .O(gate40inter8));
  nand2 gate226(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate227(.a(s_3), .b(gate40inter3), .O(gate40inter10));
  nor2  gate228(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate229(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate230(.a(gate40inter12), .b(gate40inter1), .O(N289));
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate469(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate470(.a(gate42inter0), .b(s_38), .O(gate42inter1));
  and2  gate471(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate472(.a(s_38), .O(gate42inter3));
  inv1  gate473(.a(s_39), .O(gate42inter4));
  nand2 gate474(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate475(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate476(.a(N252), .O(gate42inter7));
  inv1  gate477(.a(N253), .O(gate42inter8));
  nand2 gate478(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate479(.a(s_39), .b(gate42inter3), .O(gate42inter10));
  nor2  gate480(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate481(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate482(.a(gate42inter12), .b(gate42inter1), .O(N293));
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );

  xor2  gate385(.a(N265), .b(N264), .O(gate48inter0));
  nand2 gate386(.a(gate48inter0), .b(s_26), .O(gate48inter1));
  and2  gate387(.a(N265), .b(N264), .O(gate48inter2));
  inv1  gate388(.a(s_26), .O(gate48inter3));
  inv1  gate389(.a(s_27), .O(gate48inter4));
  nand2 gate390(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate391(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate392(.a(N264), .O(gate48inter7));
  inv1  gate393(.a(N265), .O(gate48inter8));
  nand2 gate394(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate395(.a(s_27), .b(gate48inter3), .O(gate48inter10));
  nor2  gate396(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate397(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate398(.a(gate48inter12), .b(gate48inter1), .O(N311));
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate553(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate554(.a(gate50inter0), .b(s_50), .O(gate50inter1));
  and2  gate555(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate556(.a(s_50), .O(gate50inter3));
  inv1  gate557(.a(s_51), .O(gate50inter4));
  nand2 gate558(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate559(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate560(.a(N276), .O(gate50inter7));
  inv1  gate561(.a(N277), .O(gate50inter8));
  nand2 gate562(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate563(.a(s_51), .b(gate50inter3), .O(gate50inter10));
  nor2  gate564(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate565(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate566(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );

  xor2  gate371(.a(N283), .b(N282), .O(gate53inter0));
  nand2 gate372(.a(gate53inter0), .b(s_24), .O(gate53inter1));
  and2  gate373(.a(N283), .b(N282), .O(gate53inter2));
  inv1  gate374(.a(s_24), .O(gate53inter3));
  inv1  gate375(.a(s_25), .O(gate53inter4));
  nand2 gate376(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate377(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate378(.a(N282), .O(gate53inter7));
  inv1  gate379(.a(N283), .O(gate53inter8));
  nand2 gate380(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate381(.a(s_25), .b(gate53inter3), .O(gate53inter10));
  nor2  gate382(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate383(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate384(.a(gate53inter12), .b(gate53inter1), .O(N318));
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate399(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate400(.a(gate55inter0), .b(s_28), .O(gate55inter1));
  and2  gate401(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate402(.a(s_28), .O(gate55inter3));
  inv1  gate403(.a(s_29), .O(gate55inter4));
  nand2 gate404(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate405(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate406(.a(N286), .O(gate55inter7));
  inv1  gate407(.a(N287), .O(gate55inter8));
  nand2 gate408(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate409(.a(s_29), .b(gate55inter3), .O(gate55inter10));
  nor2  gate410(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate411(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate412(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );

  xor2  gate441(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate442(.a(gate57inter0), .b(s_34), .O(gate57inter1));
  and2  gate443(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate444(.a(s_34), .O(gate57inter3));
  inv1  gate445(.a(s_35), .O(gate57inter4));
  nand2 gate446(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate447(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate448(.a(N290), .O(gate57inter7));
  inv1  gate449(.a(N293), .O(gate57inter8));
  nand2 gate450(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate451(.a(s_35), .b(gate57inter3), .O(gate57inter10));
  nor2  gate452(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate453(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate454(.a(gate57inter12), .b(gate57inter1), .O(N338));
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );

  xor2  gate357(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate358(.a(gate67inter0), .b(s_22), .O(gate67inter1));
  and2  gate359(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate360(.a(s_22), .O(gate67inter3));
  inv1  gate361(.a(s_23), .O(gate67inter4));
  nand2 gate362(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate363(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate364(.a(N268), .O(gate67inter7));
  inv1  gate365(.a(N344), .O(gate67inter8));
  nand2 gate366(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate367(.a(s_23), .b(gate67inter3), .O(gate67inter10));
  nor2  gate368(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate369(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate370(.a(gate67inter12), .b(gate67inter1), .O(N348));

  xor2  gate497(.a(N345), .b(N269), .O(gate68inter0));
  nand2 gate498(.a(gate68inter0), .b(s_42), .O(gate68inter1));
  and2  gate499(.a(N345), .b(N269), .O(gate68inter2));
  inv1  gate500(.a(s_42), .O(gate68inter3));
  inv1  gate501(.a(s_43), .O(gate68inter4));
  nand2 gate502(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate503(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate504(.a(N269), .O(gate68inter7));
  inv1  gate505(.a(N345), .O(gate68inter8));
  nand2 gate506(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate507(.a(s_43), .b(gate68inter3), .O(gate68inter10));
  nor2  gate508(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate509(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate510(.a(gate68inter12), .b(gate68inter1), .O(N349));
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate525(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate526(.a(gate75inter0), .b(s_46), .O(gate75inter1));
  and2  gate527(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate528(.a(s_46), .O(gate75inter3));
  inv1  gate529(.a(s_47), .O(gate75inter4));
  nand2 gate530(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate531(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate532(.a(N316), .O(gate75inter7));
  inv1  gate533(.a(N348), .O(gate75inter8));
  nand2 gate534(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate535(.a(s_47), .b(gate75inter3), .O(gate75inter10));
  nor2  gate536(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate537(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate538(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );

  xor2  gate483(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate484(.a(gate79inter0), .b(s_40), .O(gate79inter1));
  and2  gate485(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate486(.a(s_40), .O(gate79inter3));
  inv1  gate487(.a(s_41), .O(gate79inter4));
  nand2 gate488(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate489(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate490(.a(N320), .O(gate79inter7));
  inv1  gate491(.a(N352), .O(gate79inter8));
  nand2 gate492(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate493(.a(s_41), .b(gate79inter3), .O(gate79inter10));
  nor2  gate494(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate495(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate496(.a(gate79inter12), .b(gate79inter1), .O(N432));
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );

  xor2  gate301(.a(N696), .b(N17), .O(gate175inter0));
  nand2 gate302(.a(gate175inter0), .b(s_14), .O(gate175inter1));
  and2  gate303(.a(N696), .b(N17), .O(gate175inter2));
  inv1  gate304(.a(s_14), .O(gate175inter3));
  inv1  gate305(.a(s_15), .O(gate175inter4));
  nand2 gate306(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate307(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate308(.a(N17), .O(gate175inter7));
  inv1  gate309(.a(N696), .O(gate175inter8));
  nand2 gate310(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate311(.a(s_15), .b(gate175inter3), .O(gate175inter10));
  nor2  gate312(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate313(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate314(.a(gate175inter12), .b(gate175inter1), .O(N728));
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate203(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate204(.a(gate177inter0), .b(s_0), .O(gate177inter1));
  and2  gate205(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate206(.a(s_0), .O(gate177inter3));
  inv1  gate207(.a(s_1), .O(gate177inter4));
  nand2 gate208(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate209(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate210(.a(N25), .O(gate177inter7));
  inv1  gate211(.a(N698), .O(gate177inter8));
  nand2 gate212(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate213(.a(s_1), .b(gate177inter3), .O(gate177inter10));
  nor2  gate214(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate215(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate216(.a(gate177inter12), .b(gate177inter1), .O(N730));
xor2 gate178( .a(N29), .b(N699), .O(N731) );
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );

  xor2  gate455(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate456(.a(gate181inter0), .b(s_36), .O(gate181inter1));
  and2  gate457(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate458(.a(s_36), .O(gate181inter3));
  inv1  gate459(.a(s_37), .O(gate181inter4));
  nand2 gate460(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate461(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate462(.a(N41), .O(gate181inter7));
  inv1  gate463(.a(N702), .O(gate181inter8));
  nand2 gate464(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate465(.a(s_37), .b(gate181inter3), .O(gate181inter10));
  nor2  gate466(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate467(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate468(.a(gate181inter12), .b(gate181inter1), .O(N734));
xor2 gate182( .a(N45), .b(N703), .O(N735) );

  xor2  gate427(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate428(.a(gate183inter0), .b(s_32), .O(gate183inter1));
  and2  gate429(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate430(.a(s_32), .O(gate183inter3));
  inv1  gate431(.a(s_33), .O(gate183inter4));
  nand2 gate432(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate433(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate434(.a(N49), .O(gate183inter7));
  inv1  gate435(.a(N704), .O(gate183inter8));
  nand2 gate436(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate437(.a(s_33), .b(gate183inter3), .O(gate183inter10));
  nor2  gate438(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate439(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate440(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );
xor2 gate190( .a(N77), .b(N711), .O(N743) );
xor2 gate191( .a(N81), .b(N712), .O(N744) );

  xor2  gate539(.a(N713), .b(N85), .O(gate192inter0));
  nand2 gate540(.a(gate192inter0), .b(s_48), .O(gate192inter1));
  and2  gate541(.a(N713), .b(N85), .O(gate192inter2));
  inv1  gate542(.a(s_48), .O(gate192inter3));
  inv1  gate543(.a(s_49), .O(gate192inter4));
  nand2 gate544(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate545(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate546(.a(N85), .O(gate192inter7));
  inv1  gate547(.a(N713), .O(gate192inter8));
  nand2 gate548(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate549(.a(s_49), .b(gate192inter3), .O(gate192inter10));
  nor2  gate550(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate551(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate552(.a(gate192inter12), .b(gate192inter1), .O(N745));

  xor2  gate287(.a(N714), .b(N89), .O(gate193inter0));
  nand2 gate288(.a(gate193inter0), .b(s_12), .O(gate193inter1));
  and2  gate289(.a(N714), .b(N89), .O(gate193inter2));
  inv1  gate290(.a(s_12), .O(gate193inter3));
  inv1  gate291(.a(s_13), .O(gate193inter4));
  nand2 gate292(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate293(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate294(.a(N89), .O(gate193inter7));
  inv1  gate295(.a(N714), .O(gate193inter8));
  nand2 gate296(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate297(.a(s_13), .b(gate193inter3), .O(gate193inter10));
  nor2  gate298(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate299(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate300(.a(gate193inter12), .b(gate193inter1), .O(N746));
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );

  xor2  gate245(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate246(.a(gate198inter0), .b(s_6), .O(gate198inter1));
  and2  gate247(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate248(.a(s_6), .O(gate198inter3));
  inv1  gate249(.a(s_7), .O(gate198inter4));
  nand2 gate250(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate251(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate252(.a(N109), .O(gate198inter7));
  inv1  gate253(.a(N719), .O(gate198inter8));
  nand2 gate254(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate255(.a(s_7), .b(gate198inter3), .O(gate198inter10));
  nor2  gate256(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate257(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate258(.a(gate198inter12), .b(gate198inter1), .O(N751));
xor2 gate199( .a(N113), .b(N720), .O(N752) );

  xor2  gate413(.a(N721), .b(N117), .O(gate200inter0));
  nand2 gate414(.a(gate200inter0), .b(s_30), .O(gate200inter1));
  and2  gate415(.a(N721), .b(N117), .O(gate200inter2));
  inv1  gate416(.a(s_30), .O(gate200inter3));
  inv1  gate417(.a(s_31), .O(gate200inter4));
  nand2 gate418(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate419(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate420(.a(N117), .O(gate200inter7));
  inv1  gate421(.a(N721), .O(gate200inter8));
  nand2 gate422(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate423(.a(s_31), .b(gate200inter3), .O(gate200inter10));
  nor2  gate424(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate425(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate426(.a(gate200inter12), .b(gate200inter1), .O(N753));
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule